magic
tech sky130B
magscale 1 2
timestamp 1680008478
<< viali >>
rect 2973 42245 3007 42279
rect 6929 42245 6963 42279
rect 13369 42245 13403 42279
rect 28549 42245 28583 42279
rect 32413 42245 32447 42279
rect 35541 42245 35575 42279
rect 41889 42245 41923 42279
rect 2421 42177 2455 42211
rect 5917 42177 5951 42211
rect 9781 42177 9815 42211
rect 12449 42177 12483 42211
rect 13461 42177 13495 42211
rect 14657 42177 14691 42211
rect 14749 42177 14783 42211
rect 17233 42177 17267 42211
rect 18153 42177 18187 42211
rect 20821 42177 20855 42211
rect 24593 42177 24627 42211
rect 27261 42177 27295 42211
rect 28181 42177 28215 42211
rect 30573 42177 30607 42211
rect 31585 42177 31619 42211
rect 41613 42177 41647 42211
rect 42717 42177 42751 42211
rect 5641 42109 5675 42143
rect 7021 42109 7055 42143
rect 7205 42109 7239 42143
rect 10333 42109 10367 42143
rect 12173 42109 12207 42143
rect 13645 42109 13679 42143
rect 14933 42109 14967 42143
rect 17325 42109 17359 42143
rect 17509 42109 17543 42143
rect 18705 42109 18739 42143
rect 21373 42109 21407 42143
rect 24961 42109 24995 42143
rect 30389 42109 30423 42143
rect 42993 42109 43027 42143
rect 32597 42041 32631 42075
rect 6561 41973 6595 42007
rect 13001 41973 13035 42007
rect 14289 41973 14323 42007
rect 16865 41973 16899 42007
rect 27537 41973 27571 42007
rect 31677 41973 31711 42007
rect 35633 41973 35667 42007
rect 6929 41769 6963 41803
rect 26341 41769 26375 41803
rect 24593 41633 24627 41667
rect 27629 41633 27663 41667
rect 32137 41633 32171 41667
rect 32413 41633 32447 41667
rect 34897 41633 34931 41667
rect 5549 41565 5583 41599
rect 5816 41565 5850 41599
rect 9137 41565 9171 41599
rect 12357 41565 12391 41599
rect 12624 41565 12658 41599
rect 16425 41565 16459 41599
rect 16681 41565 16715 41599
rect 17141 41565 17175 41599
rect 19625 41565 19659 41599
rect 21281 41565 21315 41599
rect 23857 41565 23891 41599
rect 28733 41565 28767 41599
rect 32873 41565 32907 41599
rect 34007 41565 34041 41599
rect 34161 41565 34195 41599
rect 37933 41565 37967 41599
rect 40049 41565 40083 41599
rect 42257 41565 42291 41599
rect 42349 41565 42383 41599
rect 42901 41565 42935 41599
rect 9404 41497 9438 41531
rect 17417 41497 17451 41531
rect 19533 41497 19567 41531
rect 21557 41497 21591 41531
rect 24869 41497 24903 41531
rect 27077 41497 27111 41531
rect 29009 41497 29043 41531
rect 33149 41497 33183 41531
rect 35164 41497 35198 41531
rect 38178 41497 38212 41531
rect 40294 41497 40328 41531
rect 43177 41497 43211 41531
rect 10517 41429 10551 41463
rect 13737 41429 13771 41463
rect 15301 41429 15335 41463
rect 18889 41429 18923 41463
rect 23029 41429 23063 41463
rect 23949 41429 23983 41463
rect 30665 41429 30699 41463
rect 33793 41429 33827 41463
rect 36277 41429 36311 41463
rect 39313 41429 39347 41463
rect 41429 41429 41463 41463
rect 9597 41225 9631 41259
rect 12173 41225 12207 41259
rect 17417 41225 17451 41259
rect 22385 41225 22419 41259
rect 38025 41225 38059 41259
rect 39957 41225 39991 41259
rect 14188 41157 14222 41191
rect 17233 41157 17267 41191
rect 19717 41157 19751 41191
rect 32321 41157 32355 41191
rect 35786 41157 35820 41191
rect 38761 41157 38795 41191
rect 7665 41089 7699 41123
rect 7932 41089 7966 41123
rect 9965 41089 9999 41123
rect 12081 41089 12115 41123
rect 15853 41089 15887 41123
rect 17509 41089 17543 41123
rect 18061 41089 18095 41123
rect 22293 41089 22327 41123
rect 23213 41089 23247 41123
rect 24133 41089 24167 41123
rect 25237 41089 25271 41123
rect 25513 41089 25547 41123
rect 26433 41089 26467 41123
rect 27261 41089 27295 41123
rect 28365 41089 28399 41123
rect 28549 41089 28583 41123
rect 28641 41089 28675 41123
rect 28733 41089 28767 41123
rect 30297 41089 30331 41123
rect 30389 41089 30423 41123
rect 31125 41089 31159 41123
rect 31677 41089 31711 41123
rect 32468 41089 32502 41123
rect 33701 41089 33735 41123
rect 33885 41089 33919 41123
rect 34559 41089 34593 41123
rect 34713 41089 34747 41123
rect 35541 41089 35575 41123
rect 37657 41089 37691 41123
rect 38945 41089 38979 41123
rect 39129 41089 39163 41123
rect 39773 41089 39807 41123
rect 40857 41089 40891 41123
rect 42901 41089 42935 41123
rect 10057 41021 10091 41055
rect 10149 41021 10183 41055
rect 12265 41021 12299 41055
rect 13921 41021 13955 41055
rect 16129 41021 16163 41055
rect 18337 41021 18371 41055
rect 19441 41021 19475 41055
rect 21189 41021 21223 41055
rect 24685 41021 24719 41055
rect 26249 41021 26283 41055
rect 27813 41021 27847 41055
rect 29469 41021 29503 41055
rect 29837 41021 29871 41055
rect 32689 41021 32723 41055
rect 37565 41021 37599 41055
rect 39589 41021 39623 41055
rect 40601 41021 40635 41055
rect 43177 41021 43211 41055
rect 29929 40953 29963 40987
rect 32597 40953 32631 40987
rect 34345 40953 34379 40987
rect 9045 40885 9079 40919
rect 11713 40885 11747 40919
rect 15301 40885 15335 40919
rect 16957 40885 16991 40919
rect 23489 40885 23523 40919
rect 26617 40885 26651 40919
rect 29009 40885 29043 40919
rect 31585 40885 31619 40919
rect 32781 40885 32815 40919
rect 33517 40885 33551 40919
rect 36921 40885 36955 40919
rect 41981 40885 42015 40919
rect 12265 40681 12299 40715
rect 16221 40681 16255 40715
rect 20361 40681 20395 40715
rect 22983 40681 23017 40715
rect 30297 40681 30331 40715
rect 32413 40681 32447 40715
rect 35081 40681 35115 40715
rect 36093 40681 36127 40715
rect 38485 40681 38519 40715
rect 40601 40681 40635 40715
rect 15117 40613 15151 40647
rect 18245 40613 18279 40647
rect 26341 40613 26375 40647
rect 30205 40613 30239 40647
rect 35633 40613 35667 40647
rect 5917 40545 5951 40579
rect 7113 40545 7147 40579
rect 16865 40545 16899 40579
rect 21189 40545 21223 40579
rect 27445 40545 27479 40579
rect 30113 40545 30147 40579
rect 32505 40545 32539 40579
rect 35173 40545 35207 40579
rect 40141 40545 40175 40579
rect 5641 40477 5675 40511
rect 9597 40477 9631 40511
rect 9781 40477 9815 40511
rect 9873 40477 9907 40511
rect 10885 40477 10919 40511
rect 16405 40477 16439 40511
rect 17141 40477 17175 40511
rect 20269 40477 20303 40511
rect 21557 40477 21591 40511
rect 23857 40477 23891 40511
rect 24041 40477 24075 40511
rect 24593 40477 24627 40511
rect 24869 40477 24903 40511
rect 25697 40477 25731 40511
rect 25973 40477 26007 40511
rect 26985 40477 27019 40511
rect 27077 40477 27111 40511
rect 27905 40477 27939 40511
rect 28089 40477 28123 40511
rect 28733 40477 28767 40511
rect 28825 40477 28859 40511
rect 30665 40477 30699 40511
rect 31309 40477 31343 40511
rect 31953 40477 31987 40511
rect 32045 40477 32079 40511
rect 33333 40477 33367 40511
rect 33517 40477 33551 40511
rect 34161 40477 34195 40511
rect 34253 40477 34287 40511
rect 34897 40477 34931 40511
rect 34989 40477 35023 40511
rect 35909 40477 35943 40511
rect 36185 40477 36219 40511
rect 38393 40477 38427 40511
rect 38577 40477 38611 40511
rect 40233 40477 40267 40511
rect 41889 40477 41923 40511
rect 6929 40409 6963 40443
rect 9137 40409 9171 40443
rect 11152 40409 11186 40443
rect 14565 40409 14599 40443
rect 14657 40409 14691 40443
rect 14841 40409 14875 40443
rect 26065 40409 26099 40443
rect 26182 40409 26216 40443
rect 27169 40409 27203 40443
rect 27307 40409 27341 40443
rect 27997 40409 28031 40443
rect 29101 40409 29135 40443
rect 29193 40409 29227 40443
rect 31217 40409 31251 40443
rect 33701 40409 33735 40443
rect 42156 40409 42190 40443
rect 5273 40341 5307 40375
rect 5733 40341 5767 40375
rect 6469 40341 6503 40375
rect 6837 40341 6871 40375
rect 23949 40341 23983 40375
rect 26801 40341 26835 40375
rect 28549 40341 28583 40375
rect 29837 40341 29871 40375
rect 32781 40341 32815 40375
rect 43269 40341 43303 40375
rect 6009 40137 6043 40171
rect 7021 40137 7055 40171
rect 8401 40137 8435 40171
rect 8861 40137 8895 40171
rect 12081 40137 12115 40171
rect 12173 40137 12207 40171
rect 14289 40137 14323 40171
rect 26417 40137 26451 40171
rect 35633 40137 35667 40171
rect 42625 40137 42659 40171
rect 4896 40069 4930 40103
rect 6929 40069 6963 40103
rect 8769 40069 8803 40103
rect 17049 40069 17083 40103
rect 18337 40069 18371 40103
rect 26617 40069 26651 40103
rect 29929 40069 29963 40103
rect 38729 40069 38763 40103
rect 38945 40069 38979 40103
rect 42993 40069 43027 40103
rect 10425 40001 10459 40035
rect 10609 40001 10643 40035
rect 17233 40001 17267 40035
rect 17325 40001 17359 40035
rect 17785 40001 17819 40035
rect 18153 40001 18187 40035
rect 22293 40001 22327 40035
rect 22385 40001 22419 40035
rect 23397 40001 23431 40035
rect 23857 40001 23891 40035
rect 24409 40001 24443 40035
rect 24961 40001 24995 40035
rect 27629 40001 27663 40035
rect 27997 40001 28031 40035
rect 30205 40001 30239 40035
rect 31033 40001 31067 40035
rect 31493 40001 31527 40035
rect 33425 40001 33459 40035
rect 34253 40001 34287 40035
rect 34520 40001 34554 40035
rect 4629 39933 4663 39967
rect 7113 39933 7147 39967
rect 8953 39933 8987 39967
rect 9965 39933 9999 39967
rect 10701 39933 10735 39967
rect 12265 39933 12299 39967
rect 13277 39933 13311 39967
rect 23949 39933 23983 39967
rect 27537 39933 27571 39967
rect 27905 39933 27939 39967
rect 32873 39933 32907 39967
rect 43085 39933 43119 39967
rect 43177 39933 43211 39967
rect 17049 39865 17083 39899
rect 6561 39797 6595 39831
rect 11713 39797 11747 39831
rect 26249 39797 26283 39831
rect 26433 39797 26467 39831
rect 27353 39797 27387 39831
rect 31677 39797 31711 39831
rect 38577 39797 38611 39831
rect 38761 39797 38795 39831
rect 18337 39593 18371 39627
rect 21005 39593 21039 39627
rect 21189 39593 21223 39627
rect 23857 39593 23891 39627
rect 24041 39593 24075 39627
rect 27629 39593 27663 39627
rect 31769 39593 31803 39627
rect 33057 39593 33091 39627
rect 34345 39593 34379 39627
rect 37749 39593 37783 39627
rect 38669 39593 38703 39627
rect 32229 39525 32263 39559
rect 6561 39457 6595 39491
rect 27261 39457 27295 39491
rect 31953 39457 31987 39491
rect 6653 39389 6687 39423
rect 9137 39389 9171 39423
rect 9413 39389 9447 39423
rect 10425 39389 10459 39423
rect 10609 39389 10643 39423
rect 11621 39389 11655 39423
rect 16221 39389 16255 39423
rect 16405 39389 16439 39423
rect 17509 39389 17543 39423
rect 18245 39389 18279 39423
rect 18429 39389 18463 39423
rect 20177 39389 20211 39423
rect 20361 39389 20395 39423
rect 20821 39389 20855 39423
rect 20913 39389 20947 39423
rect 22937 39389 22971 39423
rect 23121 39389 23155 39423
rect 23765 39389 23799 39423
rect 23857 39389 23891 39423
rect 27445 39389 27479 39423
rect 30113 39389 30147 39423
rect 30389 39389 30423 39423
rect 30481 39389 30515 39423
rect 32045 39389 32079 39423
rect 33885 39389 33919 39423
rect 34161 39389 34195 39423
rect 34989 39389 35023 39423
rect 36553 39389 36587 39423
rect 37105 39389 37139 39423
rect 37198 39389 37232 39423
rect 37381 39389 37415 39423
rect 37611 39389 37645 39423
rect 38945 39389 38979 39423
rect 40049 39389 40083 39423
rect 42901 39389 42935 39423
rect 7113 39321 7147 39355
rect 9505 39321 9539 39355
rect 11897 39321 11931 39355
rect 23581 39321 23615 39355
rect 31769 39321 31803 39355
rect 32781 39321 32815 39355
rect 35357 39321 35391 39355
rect 36277 39321 36311 39355
rect 37473 39321 37507 39355
rect 38669 39321 38703 39355
rect 38853 39321 38887 39355
rect 40294 39321 40328 39355
rect 43177 39321 43211 39355
rect 10793 39253 10827 39287
rect 16313 39253 16347 39287
rect 17693 39253 17727 39287
rect 20269 39253 20303 39287
rect 23029 39253 23063 39287
rect 30573 39253 30607 39287
rect 33977 39253 34011 39287
rect 41429 39253 41463 39287
rect 15761 39049 15795 39083
rect 16957 39049 16991 39083
rect 18521 39049 18555 39083
rect 20085 39049 20119 39083
rect 21465 39049 21499 39083
rect 25145 39049 25179 39083
rect 26525 39049 26559 39083
rect 27169 39049 27203 39083
rect 36921 39049 36955 39083
rect 38117 39049 38151 39083
rect 39129 39049 39163 39083
rect 8769 38981 8803 39015
rect 8953 38981 8987 39015
rect 13277 38981 13311 39015
rect 15301 38981 15335 39015
rect 28917 38981 28951 39015
rect 34161 38981 34195 39015
rect 36553 38981 36587 39015
rect 36645 38981 36679 39015
rect 37749 38981 37783 39015
rect 5825 38913 5859 38947
rect 6009 38913 6043 38947
rect 7389 38913 7423 38947
rect 7481 38913 7515 38947
rect 9965 38913 9999 38947
rect 10701 38913 10735 38947
rect 11897 38913 11931 38947
rect 13185 38913 13219 38947
rect 13461 38913 13495 38947
rect 14105 38913 14139 38947
rect 14841 38913 14875 38947
rect 15577 38913 15611 38947
rect 16865 38913 16899 38947
rect 17049 38913 17083 38947
rect 18705 38913 18739 38947
rect 18797 38913 18831 38947
rect 18889 38913 18923 38947
rect 19441 38913 19475 38947
rect 19901 38913 19935 38947
rect 20821 38913 20855 38947
rect 21281 38913 21315 38947
rect 23305 38913 23339 38947
rect 24501 38913 24535 38947
rect 24961 38913 24995 38947
rect 26341 38913 26375 38947
rect 26617 38913 26651 38947
rect 27353 38913 27387 38947
rect 27445 38913 27479 38947
rect 27629 38913 27663 38947
rect 27721 38913 27755 38947
rect 28181 38913 28215 38947
rect 28365 38913 28399 38947
rect 29193 38913 29227 38947
rect 30113 38913 30147 38947
rect 30389 38913 30423 38947
rect 31401 38913 31435 38947
rect 33149 38913 33183 38947
rect 33885 38913 33919 38947
rect 34805 38913 34839 38947
rect 36277 38913 36311 38947
rect 36425 38913 36459 38947
rect 36783 38913 36817 38947
rect 37473 38913 37507 38947
rect 37621 38913 37655 38947
rect 37841 38913 37875 38947
rect 37938 38913 37972 38947
rect 39037 38913 39071 38947
rect 39221 38913 39255 38947
rect 42993 38913 43027 38947
rect 6929 38845 6963 38879
rect 10977 38845 11011 38879
rect 12081 38845 12115 38879
rect 14473 38845 14507 38879
rect 15393 38845 15427 38879
rect 19809 38845 19843 38879
rect 21097 38845 21131 38879
rect 22845 38845 22879 38879
rect 23397 38845 23431 38879
rect 24869 38845 24903 38879
rect 29653 38845 29687 38879
rect 31493 38845 31527 38879
rect 32873 38845 32907 38879
rect 35081 38845 35115 38879
rect 43085 38845 43119 38879
rect 43177 38845 43211 38879
rect 22753 38777 22787 38811
rect 29101 38777 29135 38811
rect 30297 38777 30331 38811
rect 34897 38777 34931 38811
rect 5917 38709 5951 38743
rect 8585 38709 8619 38743
rect 8769 38709 8803 38743
rect 13645 38709 13679 38743
rect 15301 38709 15335 38743
rect 19533 38709 19567 38743
rect 20913 38709 20947 38743
rect 22937 38709 22971 38743
rect 24593 38709 24627 38743
rect 26157 38709 26191 38743
rect 28181 38709 28215 38743
rect 29009 38709 29043 38743
rect 31401 38709 31435 38743
rect 31769 38709 31803 38743
rect 35265 38709 35299 38743
rect 42625 38709 42659 38743
rect 14473 38505 14507 38539
rect 17693 38505 17727 38539
rect 19441 38505 19475 38539
rect 19809 38505 19843 38539
rect 20269 38505 20303 38539
rect 20729 38505 20763 38539
rect 21189 38505 21223 38539
rect 21373 38505 21407 38539
rect 23949 38505 23983 38539
rect 24869 38505 24903 38539
rect 36921 38505 36955 38539
rect 38117 38505 38151 38539
rect 40693 38505 40727 38539
rect 14933 38437 14967 38471
rect 23213 38437 23247 38471
rect 28365 38437 28399 38471
rect 30389 38437 30423 38471
rect 39497 38437 39531 38471
rect 10149 38369 10183 38403
rect 13001 38369 13035 38403
rect 13093 38369 13127 38403
rect 14657 38369 14691 38403
rect 18797 38369 18831 38403
rect 20453 38369 20487 38403
rect 21557 38369 21591 38403
rect 23765 38369 23799 38403
rect 24869 38369 24903 38403
rect 27261 38369 27295 38403
rect 29745 38369 29779 38403
rect 41797 38369 41831 38403
rect 5825 38301 5859 38335
rect 5917 38301 5951 38335
rect 7021 38301 7055 38335
rect 7113 38301 7147 38335
rect 7573 38301 7607 38335
rect 7941 38301 7975 38335
rect 8125 38301 8159 38335
rect 9229 38301 9263 38335
rect 10333 38301 10367 38335
rect 11529 38301 11563 38335
rect 11897 38301 11931 38335
rect 13461 38301 13495 38335
rect 14749 38301 14783 38335
rect 16129 38301 16163 38335
rect 16221 38301 16255 38335
rect 16405 38301 16439 38335
rect 16497 38301 16531 38335
rect 17509 38301 17543 38335
rect 17693 38301 17727 38335
rect 18705 38301 18739 38335
rect 18889 38301 18923 38335
rect 19717 38301 19751 38335
rect 19809 38301 19843 38335
rect 20269 38301 20303 38335
rect 20545 38301 20579 38335
rect 21373 38301 21407 38335
rect 23121 38301 23155 38335
rect 23305 38301 23339 38335
rect 24041 38301 24075 38335
rect 25053 38301 25087 38335
rect 27077 38301 27111 38335
rect 27169 38301 27203 38335
rect 27353 38301 27387 38335
rect 30205 38301 30239 38335
rect 30481 38301 30515 38335
rect 31493 38301 31527 38335
rect 31769 38301 31803 38335
rect 32689 38301 32723 38335
rect 32781 38301 32815 38335
rect 32873 38301 32907 38335
rect 33057 38301 33091 38335
rect 34253 38301 34287 38335
rect 34897 38301 34931 38335
rect 35081 38301 35115 38335
rect 36277 38301 36311 38335
rect 36370 38301 36404 38335
rect 36645 38301 36679 38335
rect 36742 38301 36776 38335
rect 37473 38301 37507 38335
rect 37621 38301 37655 38335
rect 37938 38301 37972 38335
rect 38945 38301 38979 38335
rect 39221 38301 39255 38335
rect 39313 38301 39347 38335
rect 40049 38301 40083 38335
rect 40142 38301 40176 38335
rect 40417 38301 40451 38335
rect 40555 38301 40589 38335
rect 42064 38301 42098 38335
rect 6561 38233 6595 38267
rect 12081 38233 12115 38267
rect 14473 38233 14507 38267
rect 21649 38233 21683 38267
rect 24593 38233 24627 38267
rect 27997 38233 28031 38267
rect 31677 38233 31711 38267
rect 33793 38233 33827 38267
rect 36553 38233 36587 38267
rect 37749 38233 37783 38267
rect 37841 38233 37875 38267
rect 39129 38233 39163 38267
rect 40325 38233 40359 38267
rect 6101 38165 6135 38199
rect 13277 38165 13311 38199
rect 13369 38165 13403 38199
rect 13737 38165 13771 38199
rect 16681 38165 16715 38199
rect 17877 38165 17911 38199
rect 23765 38165 23799 38199
rect 25237 38165 25271 38199
rect 26893 38165 26927 38199
rect 28457 38165 28491 38199
rect 32413 38165 32447 38199
rect 34989 38165 35023 38199
rect 43177 38165 43211 38199
rect 18245 37961 18279 37995
rect 23581 37961 23615 37995
rect 25053 37961 25087 37995
rect 29745 37961 29779 37995
rect 34621 37961 34655 37995
rect 36461 37961 36495 37995
rect 41245 37961 41279 37995
rect 7113 37893 7147 37927
rect 14565 37893 14599 37927
rect 16129 37893 16163 37927
rect 19717 37893 19751 37927
rect 34069 37893 34103 37927
rect 34989 37893 35023 37927
rect 40969 37893 41003 37927
rect 4261 37825 4295 37859
rect 4528 37825 4562 37859
rect 7297 37825 7331 37859
rect 7941 37825 7975 37859
rect 8125 37825 8159 37859
rect 8217 37825 8251 37859
rect 9045 37825 9079 37859
rect 10057 37825 10091 37859
rect 10977 37825 11011 37859
rect 11897 37825 11931 37859
rect 11989 37825 12023 37859
rect 12173 37825 12207 37859
rect 12265 37825 12299 37859
rect 12725 37825 12759 37859
rect 12909 37825 12943 37859
rect 13829 37825 13863 37859
rect 14013 37825 14047 37859
rect 14105 37825 14139 37859
rect 14381 37825 14415 37859
rect 15945 37825 15979 37859
rect 16037 37825 16071 37859
rect 16865 37825 16899 37859
rect 17049 37825 17083 37859
rect 17785 37825 17819 37859
rect 17969 37825 18003 37859
rect 18061 37825 18095 37859
rect 19901 37825 19935 37859
rect 20000 37825 20034 37859
rect 22201 37825 22235 37859
rect 22569 37825 22603 37859
rect 22753 37825 22787 37859
rect 23397 37825 23431 37859
rect 24409 37825 24443 37859
rect 24869 37825 24903 37859
rect 25881 37825 25915 37859
rect 26157 37825 26191 37859
rect 27169 37825 27203 37859
rect 27353 37825 27387 37859
rect 28733 37825 28767 37859
rect 28917 37825 28951 37859
rect 29377 37825 29411 37859
rect 30205 37825 30239 37859
rect 30389 37825 30423 37859
rect 31585 37825 31619 37859
rect 32321 37825 32355 37859
rect 32505 37825 32539 37859
rect 33793 37825 33827 37859
rect 33885 37825 33919 37859
rect 34805 37825 34839 37859
rect 35817 37825 35851 37859
rect 35910 37825 35944 37859
rect 36093 37825 36127 37859
rect 36185 37825 36219 37859
rect 36323 37825 36357 37859
rect 37565 37825 37599 37859
rect 38853 37825 38887 37859
rect 39037 37825 39071 37859
rect 39129 37825 39163 37859
rect 39221 37825 39255 37859
rect 40601 37825 40635 37859
rect 40694 37825 40728 37859
rect 40877 37825 40911 37859
rect 41107 37825 41141 37859
rect 42901 37825 42935 37859
rect 7481 37757 7515 37791
rect 10701 37757 10735 37791
rect 10793 37757 10827 37791
rect 14197 37757 14231 37791
rect 20085 37757 20119 37791
rect 22385 37757 22419 37791
rect 22477 37757 22511 37791
rect 23213 37757 23247 37791
rect 24777 37757 24811 37791
rect 25973 37757 26007 37791
rect 29469 37757 29503 37791
rect 31309 37757 31343 37791
rect 38117 37757 38151 37791
rect 43177 37757 43211 37791
rect 8401 37689 8435 37723
rect 13093 37689 13127 37723
rect 15761 37689 15795 37723
rect 17877 37689 17911 37723
rect 31769 37689 31803 37723
rect 39405 37689 39439 37723
rect 5641 37621 5675 37655
rect 8217 37621 8251 37655
rect 9965 37621 9999 37655
rect 11161 37621 11195 37655
rect 11713 37621 11747 37655
rect 16313 37621 16347 37655
rect 17233 37621 17267 37655
rect 22017 37621 22051 37655
rect 24777 37621 24811 37655
rect 25697 37621 25731 37655
rect 26157 37621 26191 37655
rect 27169 37621 27203 37655
rect 28733 37621 28767 37655
rect 29561 37621 29595 37655
rect 30205 37621 30239 37655
rect 31401 37621 31435 37655
rect 32597 37621 32631 37655
rect 4905 37417 4939 37451
rect 12449 37417 12483 37451
rect 12541 37417 12575 37451
rect 14565 37417 14599 37451
rect 20453 37417 20487 37451
rect 22569 37417 22603 37451
rect 25145 37417 25179 37451
rect 26893 37417 26927 37451
rect 37289 37417 37323 37451
rect 39497 37417 39531 37451
rect 9873 37349 9907 37383
rect 11529 37349 11563 37383
rect 11621 37349 11655 37383
rect 25605 37349 25639 37383
rect 35817 37349 35851 37383
rect 5457 37281 5491 37315
rect 6837 37281 6871 37315
rect 9961 37281 9995 37315
rect 12633 37281 12667 37315
rect 16589 37281 16623 37315
rect 17141 37281 17175 37315
rect 20545 37281 20579 37315
rect 26709 37281 26743 37315
rect 32781 37281 32815 37315
rect 35081 37281 35115 37315
rect 6561 37213 6595 37247
rect 6745 37213 6779 37247
rect 7389 37213 7423 37247
rect 7665 37213 7699 37247
rect 8217 37213 8251 37247
rect 9781 37213 9815 37247
rect 10057 37213 10091 37247
rect 10333 37213 10367 37247
rect 11437 37213 11471 37247
rect 11713 37213 11747 37247
rect 12357 37213 12391 37247
rect 14473 37213 14507 37247
rect 16773 37213 16807 37247
rect 20453 37213 20487 37247
rect 20729 37213 20763 37247
rect 22661 37213 22695 37247
rect 24869 37213 24903 37247
rect 24961 37213 24995 37247
rect 25789 37213 25823 37247
rect 26985 37213 27019 37247
rect 27813 37213 27847 37247
rect 28825 37213 28859 37247
rect 29101 37213 29135 37247
rect 29193 37213 29227 37247
rect 30021 37213 30055 37247
rect 30297 37213 30331 37247
rect 32137 37213 32171 37247
rect 32321 37213 32355 37247
rect 32689 37213 32723 37247
rect 33793 37213 33827 37247
rect 33885 37213 33919 37247
rect 33977 37213 34011 37247
rect 35265 37213 35299 37247
rect 35725 37213 35759 37247
rect 36645 37213 36679 37247
rect 36738 37213 36772 37247
rect 37151 37213 37185 37247
rect 38945 37213 38979 37247
rect 39221 37213 39255 37247
rect 39313 37213 39347 37247
rect 40141 37213 40175 37247
rect 40234 37213 40268 37247
rect 40509 37213 40543 37247
rect 40647 37213 40681 37247
rect 41705 37213 41739 37247
rect 5273 37145 5307 37179
rect 8401 37145 8435 37179
rect 8585 37145 8619 37179
rect 14289 37145 14323 37179
rect 17049 37145 17083 37179
rect 25145 37145 25179 37179
rect 25973 37145 26007 37179
rect 27445 37145 27479 37179
rect 27629 37145 27663 37179
rect 31309 37145 31343 37179
rect 31493 37145 31527 37179
rect 31677 37145 31711 37179
rect 33333 37145 33367 37179
rect 36921 37145 36955 37179
rect 37013 37145 37047 37179
rect 39129 37145 39163 37179
rect 40417 37145 40451 37179
rect 41972 37145 42006 37179
rect 5365 37077 5399 37111
rect 6377 37077 6411 37111
rect 7389 37077 7423 37111
rect 11897 37077 11931 37111
rect 20913 37077 20947 37111
rect 24685 37077 24719 37111
rect 26709 37077 26743 37111
rect 29837 37077 29871 37111
rect 40785 37077 40819 37111
rect 43085 37077 43119 37111
rect 13737 36873 13771 36907
rect 15853 36873 15887 36907
rect 17141 36873 17175 36907
rect 20269 36873 20303 36907
rect 24685 36873 24719 36907
rect 42625 36873 42659 36907
rect 43085 36873 43119 36907
rect 6653 36805 6687 36839
rect 17601 36805 17635 36839
rect 6837 36737 6871 36771
rect 6929 36737 6963 36771
rect 7849 36737 7883 36771
rect 8033 36737 8067 36771
rect 8953 36737 8987 36771
rect 9137 36737 9171 36771
rect 9229 36737 9263 36771
rect 10333 36737 10367 36771
rect 10977 36737 11011 36771
rect 11069 36737 11103 36771
rect 12725 36737 12759 36771
rect 13553 36737 13587 36771
rect 14662 36737 14696 36771
rect 15485 36737 15519 36771
rect 15577 36737 15611 36771
rect 16865 36737 16899 36771
rect 17233 36737 17267 36771
rect 17325 36737 17359 36771
rect 19165 36737 19199 36771
rect 20637 36737 20671 36771
rect 22109 36737 22143 36771
rect 22293 36737 22327 36771
rect 24041 36737 24075 36771
rect 24225 36737 24259 36771
rect 24869 36737 24903 36771
rect 25053 36737 25087 36771
rect 27353 36737 27387 36771
rect 27721 36737 27755 36771
rect 29745 36737 29779 36771
rect 30021 36737 30055 36771
rect 31033 36737 31067 36771
rect 31217 36737 31251 36771
rect 32321 36737 32355 36771
rect 32597 36737 32631 36771
rect 33517 36737 33551 36771
rect 33701 36737 33735 36771
rect 34345 36737 34379 36771
rect 34529 36737 34563 36771
rect 34897 36737 34931 36771
rect 36185 36737 36219 36771
rect 36369 36737 36403 36771
rect 36553 36737 36587 36771
rect 42993 36737 43027 36771
rect 9045 36669 9079 36703
rect 10057 36669 10091 36703
rect 10793 36669 10827 36703
rect 11989 36669 12023 36703
rect 13277 36669 13311 36703
rect 14749 36669 14783 36703
rect 19441 36669 19475 36703
rect 20545 36669 20579 36703
rect 22017 36669 22051 36703
rect 27261 36669 27295 36703
rect 29929 36669 29963 36703
rect 30757 36669 30791 36703
rect 33057 36669 33091 36703
rect 34805 36669 34839 36703
rect 43177 36669 43211 36703
rect 32413 36601 32447 36635
rect 33793 36601 33827 36635
rect 6745 36533 6779 36567
rect 7113 36533 7147 36567
rect 7665 36533 7699 36567
rect 9413 36533 9447 36567
rect 13369 36533 13403 36567
rect 14841 36533 14875 36567
rect 15025 36533 15059 36567
rect 15485 36533 15519 36567
rect 16957 36533 16991 36567
rect 20637 36533 20671 36567
rect 22477 36533 22511 36567
rect 24225 36533 24259 36567
rect 25053 36533 25087 36567
rect 27721 36533 27755 36567
rect 27905 36533 27939 36567
rect 35449 36533 35483 36567
rect 12449 36329 12483 36363
rect 13645 36329 13679 36363
rect 14565 36329 14599 36363
rect 14749 36329 14783 36363
rect 16037 36329 16071 36363
rect 17141 36329 17175 36363
rect 17233 36329 17267 36363
rect 17785 36329 17819 36363
rect 18521 36329 18555 36363
rect 19993 36329 20027 36363
rect 21189 36329 21223 36363
rect 23489 36329 23523 36363
rect 23949 36329 23983 36363
rect 27537 36329 27571 36363
rect 28641 36329 28675 36363
rect 30021 36329 30055 36363
rect 30316 36329 30350 36363
rect 37381 36329 37415 36363
rect 15669 36261 15703 36295
rect 16221 36261 16255 36295
rect 20959 36261 20993 36295
rect 30205 36261 30239 36295
rect 33241 36261 33275 36295
rect 34897 36261 34931 36295
rect 38117 36261 38151 36295
rect 6101 36193 6135 36227
rect 10425 36193 10459 36227
rect 14473 36193 14507 36227
rect 17325 36193 17359 36227
rect 21833 36193 21867 36227
rect 24593 36193 24627 36227
rect 27905 36193 27939 36227
rect 30113 36193 30147 36227
rect 31861 36193 31895 36227
rect 4077 36125 4111 36159
rect 6193 36125 6227 36159
rect 6837 36125 6871 36159
rect 6929 36125 6963 36159
rect 7021 36125 7055 36159
rect 7205 36125 7239 36159
rect 8309 36125 8343 36159
rect 8585 36125 8619 36159
rect 9873 36125 9907 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 11069 36125 11103 36159
rect 11345 36125 11379 36159
rect 11529 36125 11563 36159
rect 11713 36125 11747 36159
rect 12541 36125 12575 36159
rect 12633 36125 12667 36159
rect 13553 36125 13587 36159
rect 14565 36125 14599 36159
rect 17049 36125 17083 36159
rect 17785 36125 17819 36159
rect 17969 36125 18003 36159
rect 18521 36125 18555 36159
rect 18705 36125 18739 36159
rect 19441 36125 19475 36159
rect 19717 36125 19751 36159
rect 19809 36125 19843 36159
rect 20821 36125 20855 36159
rect 21097 36125 21131 36159
rect 21281 36125 21315 36159
rect 21741 36125 21775 36159
rect 21925 36125 21959 36159
rect 22569 36125 22603 36159
rect 23673 36125 23707 36159
rect 23765 36125 23799 36159
rect 24869 36125 24903 36159
rect 24961 36125 24995 36159
rect 25053 36125 25087 36159
rect 25237 36125 25271 36159
rect 27721 36125 27755 36159
rect 27813 36125 27847 36159
rect 27997 36125 28031 36159
rect 28549 36125 28583 36159
rect 28917 36125 28951 36159
rect 29009 36125 29043 36159
rect 30481 36125 30515 36159
rect 31769 36125 31803 36159
rect 32045 36125 32079 36159
rect 32965 36125 32999 36159
rect 34069 36125 34103 36159
rect 34253 36125 34287 36159
rect 35081 36125 35115 36159
rect 35633 36125 35667 36159
rect 35725 36125 35759 36159
rect 36737 36125 36771 36159
rect 36885 36125 36919 36159
rect 37105 36125 37139 36159
rect 37202 36125 37236 36159
rect 37841 36125 37875 36159
rect 38577 36125 38611 36159
rect 38761 36125 38795 36159
rect 40049 36125 40083 36159
rect 40417 36125 40451 36159
rect 41889 36125 41923 36159
rect 4344 36057 4378 36091
rect 9597 36057 9631 36091
rect 12357 36057 12391 36091
rect 13369 36057 13403 36091
rect 14289 36057 14323 36091
rect 16037 36057 16071 36091
rect 19625 36057 19659 36091
rect 22385 36057 22419 36091
rect 23489 36057 23523 36091
rect 32505 36057 32539 36091
rect 33241 36057 33275 36091
rect 37013 36057 37047 36091
rect 38117 36057 38151 36091
rect 40233 36057 40267 36091
rect 40325 36057 40359 36091
rect 42156 36057 42190 36091
rect 5457 35989 5491 36023
rect 6653 35989 6687 36023
rect 8493 35989 8527 36023
rect 11253 35989 11287 36023
rect 12817 35989 12851 36023
rect 18889 35989 18923 36023
rect 22661 35989 22695 36023
rect 29193 35989 29227 36023
rect 33057 35989 33091 36023
rect 34161 35989 34195 36023
rect 37933 35989 37967 36023
rect 38669 35989 38703 36023
rect 40601 35989 40635 36023
rect 43269 35989 43303 36023
rect 4997 35785 5031 35819
rect 8309 35785 8343 35819
rect 12081 35785 12115 35819
rect 12817 35785 12851 35819
rect 15577 35785 15611 35819
rect 20637 35785 20671 35819
rect 22017 35785 22051 35819
rect 23489 35785 23523 35819
rect 24961 35785 24995 35819
rect 31493 35785 31527 35819
rect 38301 35785 38335 35819
rect 42625 35785 42659 35819
rect 7389 35717 7423 35751
rect 7481 35717 7515 35751
rect 11897 35717 11931 35751
rect 14289 35717 14323 35751
rect 17969 35717 18003 35751
rect 18797 35717 18831 35751
rect 20177 35717 20211 35751
rect 37933 35717 37967 35751
rect 38117 35717 38151 35751
rect 7297 35649 7331 35683
rect 7665 35649 7699 35683
rect 8217 35649 8251 35683
rect 8401 35649 8435 35683
rect 8953 35649 8987 35683
rect 9229 35649 9263 35683
rect 9689 35649 9723 35683
rect 10149 35649 10183 35683
rect 11713 35649 11747 35683
rect 12909 35649 12943 35683
rect 13093 35649 13127 35683
rect 14565 35649 14599 35683
rect 15393 35649 15427 35683
rect 15577 35649 15611 35683
rect 16037 35649 16071 35683
rect 16221 35649 16255 35683
rect 16957 35649 16991 35683
rect 17141 35649 17175 35683
rect 17693 35649 17727 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 18705 35649 18739 35683
rect 18889 35649 18923 35683
rect 20453 35649 20487 35683
rect 22201 35649 22235 35683
rect 22293 35649 22327 35683
rect 22661 35649 22695 35683
rect 23489 35649 23523 35683
rect 23673 35649 23707 35683
rect 24225 35649 24259 35683
rect 25421 35649 25455 35683
rect 26065 35649 26099 35683
rect 26433 35649 26467 35683
rect 27675 35649 27709 35683
rect 29101 35649 29135 35683
rect 30113 35649 30147 35683
rect 31125 35649 31159 35683
rect 33241 35649 33275 35683
rect 33425 35649 33459 35683
rect 34161 35649 34195 35683
rect 34345 35649 34379 35683
rect 39293 35649 39327 35683
rect 40969 35649 41003 35683
rect 41062 35649 41096 35683
rect 41245 35649 41279 35683
rect 41337 35649 41371 35683
rect 41434 35649 41468 35683
rect 42993 35649 43027 35683
rect 5181 35581 5215 35615
rect 5273 35581 5307 35615
rect 5365 35581 5399 35615
rect 5457 35581 5491 35615
rect 14381 35581 14415 35615
rect 16129 35581 16163 35615
rect 17049 35581 17083 35615
rect 20361 35581 20395 35615
rect 22385 35581 22419 35615
rect 22477 35581 22511 35615
rect 25145 35581 25179 35615
rect 25973 35581 26007 35615
rect 27261 35581 27295 35615
rect 27537 35581 27571 35615
rect 30205 35581 30239 35615
rect 30389 35581 30423 35615
rect 30665 35581 30699 35615
rect 31217 35581 31251 35615
rect 33149 35581 33183 35615
rect 39037 35581 39071 35615
rect 43085 35581 43119 35615
rect 43269 35581 43303 35615
rect 9137 35513 9171 35547
rect 14749 35513 14783 35547
rect 25329 35513 25363 35547
rect 28089 35513 28123 35547
rect 41613 35513 41647 35547
rect 7113 35445 7147 35479
rect 10333 35445 10367 35479
rect 14289 35445 14323 35479
rect 18245 35445 18279 35479
rect 20453 35445 20487 35479
rect 24317 35445 24351 35479
rect 26341 35445 26375 35479
rect 26617 35445 26651 35479
rect 27721 35445 27755 35479
rect 29377 35445 29411 35479
rect 31309 35445 31343 35479
rect 34253 35445 34287 35479
rect 38117 35445 38151 35479
rect 40417 35445 40451 35479
rect 5365 35241 5399 35275
rect 14289 35241 14323 35275
rect 15669 35241 15703 35275
rect 19717 35241 19751 35275
rect 20177 35241 20211 35275
rect 22293 35241 22327 35275
rect 25145 35241 25179 35275
rect 27077 35241 27111 35275
rect 27905 35241 27939 35275
rect 29837 35241 29871 35275
rect 32321 35241 32355 35275
rect 33425 35241 33459 35275
rect 36461 35241 36495 35275
rect 14749 35173 14783 35207
rect 15853 35173 15887 35207
rect 30849 35173 30883 35207
rect 30941 35173 30975 35207
rect 33609 35173 33643 35207
rect 37565 35173 37599 35207
rect 7573 35105 7607 35139
rect 14381 35105 14415 35139
rect 26985 35105 27019 35139
rect 27169 35105 27203 35139
rect 28917 35105 28951 35139
rect 29193 35105 29227 35139
rect 30757 35105 30791 35139
rect 31861 35105 31895 35139
rect 32413 35105 32447 35139
rect 32781 35105 32815 35139
rect 38209 35105 38243 35139
rect 38669 35105 38703 35139
rect 40049 35105 40083 35139
rect 42257 35105 42291 35139
rect 5549 35037 5583 35071
rect 5641 35037 5675 35071
rect 7297 35037 7331 35071
rect 7481 35037 7515 35071
rect 7665 35037 7699 35071
rect 7849 35037 7883 35071
rect 9321 35037 9355 35071
rect 9505 35037 9539 35071
rect 10793 35037 10827 35071
rect 10977 35037 11011 35071
rect 12081 35037 12115 35071
rect 12541 35037 12575 35071
rect 14289 35037 14323 35071
rect 14565 35037 14599 35071
rect 19625 35037 19659 35071
rect 19993 35037 20027 35071
rect 22293 35037 22327 35071
rect 22477 35037 22511 35071
rect 22937 35037 22971 35071
rect 25513 35037 25547 35071
rect 26157 35037 26191 35071
rect 26249 35037 26283 35071
rect 27261 35037 27295 35071
rect 27721 35037 27755 35071
rect 27905 35037 27939 35071
rect 28733 35037 28767 35071
rect 28825 35037 28859 35071
rect 29009 35037 29043 35071
rect 29745 35037 29779 35071
rect 29929 35037 29963 35071
rect 31309 35037 31343 35071
rect 31953 35037 31987 35071
rect 34161 35037 34195 35071
rect 34345 35037 34379 35071
rect 35817 35037 35851 35071
rect 35910 35037 35944 35071
rect 36323 35037 36357 35071
rect 36921 35037 36955 35071
rect 37059 35037 37093 35071
rect 37427 35037 37461 35071
rect 38301 35037 38335 35071
rect 41981 35037 42015 35071
rect 42901 35037 42935 35071
rect 9137 34969 9171 35003
rect 15485 34969 15519 35003
rect 17233 34969 17267 35003
rect 17969 34969 18003 35003
rect 23121 34969 23155 35003
rect 23305 34969 23339 35003
rect 25329 34969 25363 35003
rect 33241 34969 33275 35003
rect 36093 34969 36127 35003
rect 36185 34969 36219 35003
rect 37197 34969 37231 35003
rect 37289 34969 37323 35003
rect 40294 34969 40328 35003
rect 43177 34969 43211 35003
rect 8033 34901 8067 34935
rect 11069 34901 11103 34935
rect 12173 34901 12207 34935
rect 15669 34901 15703 34935
rect 26065 34901 26099 34935
rect 30481 34901 30515 34935
rect 33425 34901 33459 34935
rect 34253 34901 34287 34935
rect 41429 34901 41463 34935
rect 19533 34697 19567 34731
rect 33057 34697 33091 34731
rect 36001 34697 36035 34731
rect 7573 34629 7607 34663
rect 9229 34629 9263 34663
rect 12909 34629 12943 34663
rect 13093 34629 13127 34663
rect 14473 34629 14507 34663
rect 18398 34629 18432 34663
rect 24869 34629 24903 34663
rect 25789 34629 25823 34663
rect 27813 34629 27847 34663
rect 34529 34629 34563 34663
rect 42809 34629 42843 34663
rect 4169 34561 4203 34595
rect 4436 34561 4470 34595
rect 7113 34561 7147 34595
rect 7297 34561 7331 34595
rect 8493 34561 8527 34595
rect 8677 34561 8711 34595
rect 9413 34561 9447 34595
rect 10057 34561 10091 34595
rect 10241 34561 10275 34595
rect 11713 34561 11747 34595
rect 11897 34561 11931 34595
rect 12725 34561 12759 34595
rect 13553 34561 13587 34595
rect 13829 34561 13863 34595
rect 14381 34561 14415 34595
rect 18153 34561 18187 34595
rect 23121 34561 23155 34595
rect 23213 34561 23247 34595
rect 23765 34561 23799 34595
rect 24133 34561 24167 34595
rect 25237 34561 25271 34595
rect 26157 34561 26191 34595
rect 27537 34561 27571 34595
rect 27629 34561 27663 34595
rect 28365 34561 28399 34595
rect 28733 34561 28767 34595
rect 31309 34561 31343 34595
rect 33241 34561 33275 34595
rect 33701 34561 33735 34595
rect 36139 34561 36173 34595
rect 36277 34561 36311 34595
rect 36369 34561 36403 34595
rect 36497 34561 36531 34595
rect 36645 34561 36679 34595
rect 8401 34493 8435 34527
rect 9597 34493 9631 34527
rect 11805 34493 11839 34527
rect 13921 34493 13955 34527
rect 25973 34493 26007 34527
rect 26065 34493 26099 34527
rect 28457 34493 28491 34527
rect 29009 34493 29043 34527
rect 33333 34493 33367 34527
rect 34897 34493 34931 34527
rect 35265 34493 35299 34527
rect 23029 34425 23063 34459
rect 34667 34425 34701 34459
rect 5549 34357 5583 34391
rect 6929 34357 6963 34391
rect 7481 34357 7515 34391
rect 10149 34357 10183 34391
rect 25973 34357 26007 34391
rect 28549 34357 28583 34391
rect 28641 34357 28675 34391
rect 30021 34357 30055 34391
rect 33609 34357 33643 34391
rect 34805 34357 34839 34391
rect 43085 34357 43119 34391
rect 5825 34153 5859 34187
rect 8033 34153 8067 34187
rect 26709 34153 26743 34187
rect 28181 34153 28215 34187
rect 31953 34153 31987 34187
rect 33793 34153 33827 34187
rect 35909 34153 35943 34187
rect 21649 34085 21683 34119
rect 30665 34085 30699 34119
rect 6193 34017 6227 34051
rect 10057 34017 10091 34051
rect 10241 34017 10275 34051
rect 10333 34017 10367 34051
rect 10885 34017 10919 34051
rect 13461 34017 13495 34051
rect 26617 34017 26651 34051
rect 27445 34017 27479 34051
rect 30113 34017 30147 34051
rect 35817 34017 35851 34051
rect 41889 34017 41923 34051
rect 6009 33949 6043 33983
rect 6101 33949 6135 33983
rect 6285 33949 6319 33983
rect 6469 33949 6503 33983
rect 6929 33949 6963 33983
rect 7113 33949 7147 33983
rect 8033 33949 8067 33983
rect 8309 33949 8343 33983
rect 10149 33949 10183 33983
rect 11253 33949 11287 33983
rect 11345 33949 11379 33983
rect 13369 33949 13403 33983
rect 13553 33949 13587 33983
rect 17049 33949 17083 33983
rect 19441 33949 19475 33983
rect 19533 33949 19567 33983
rect 19717 33949 19751 33983
rect 21465 33949 21499 33983
rect 21557 33949 21591 33983
rect 21741 33949 21775 33983
rect 22661 33949 22695 33983
rect 23029 33949 23063 33983
rect 23397 33949 23431 33983
rect 23765 33949 23799 33983
rect 24777 33949 24811 33983
rect 26525 33949 26559 33983
rect 27353 33949 27387 33983
rect 27537 33949 27571 33983
rect 27997 33949 28031 33983
rect 28181 33949 28215 33983
rect 29929 33949 29963 33983
rect 30573 33949 30607 33983
rect 30849 33949 30883 33983
rect 32597 33949 32631 33983
rect 32781 33949 32815 33983
rect 32873 33949 32907 33983
rect 32965 33949 32999 33983
rect 33977 33949 34011 33983
rect 34069 33949 34103 33983
rect 35081 33949 35115 33983
rect 35725 33949 35759 33983
rect 8217 33881 8251 33915
rect 11043 33881 11077 33915
rect 11161 33881 11195 33915
rect 12173 33881 12207 33915
rect 12909 33881 12943 33915
rect 16804 33881 16838 33915
rect 17509 33881 17543 33915
rect 18337 33881 18371 33915
rect 25789 33881 25823 33915
rect 32137 33881 32171 33915
rect 33793 33881 33827 33915
rect 34897 33881 34931 33915
rect 35265 33881 35299 33915
rect 42156 33881 42190 33915
rect 7021 33813 7055 33847
rect 9873 33813 9907 33847
rect 11529 33813 11563 33847
rect 15669 33813 15703 33847
rect 19901 33813 19935 33847
rect 21925 33813 21959 33847
rect 22477 33813 22511 33847
rect 26893 33813 26927 33847
rect 29745 33813 29779 33847
rect 31033 33813 31067 33847
rect 31769 33813 31803 33847
rect 31937 33813 31971 33847
rect 33241 33813 33275 33847
rect 34253 33813 34287 33847
rect 36093 33813 36127 33847
rect 43269 33813 43303 33847
rect 7113 33609 7147 33643
rect 8953 33609 8987 33643
rect 26065 33609 26099 33643
rect 27997 33609 28031 33643
rect 31769 33609 31803 33643
rect 42625 33609 42659 33643
rect 9965 33541 9999 33575
rect 12081 33541 12115 33575
rect 12909 33541 12943 33575
rect 19616 33541 19650 33575
rect 24961 33541 24995 33575
rect 26157 33541 26191 33575
rect 27537 33541 27571 33575
rect 33149 33541 33183 33575
rect 39313 33541 39347 33575
rect 39405 33541 39439 33575
rect 40785 33541 40819 33575
rect 42993 33541 43027 33575
rect 5089 33473 5123 33507
rect 6837 33473 6871 33507
rect 6929 33473 6963 33507
rect 9321 33473 9355 33507
rect 9781 33473 9815 33507
rect 10057 33473 10091 33507
rect 10609 33473 10643 33507
rect 10885 33473 10919 33507
rect 13553 33473 13587 33507
rect 13829 33473 13863 33507
rect 14289 33473 14323 33507
rect 14473 33473 14507 33507
rect 16865 33473 16899 33507
rect 17132 33473 17166 33507
rect 22109 33473 22143 33507
rect 22201 33473 22235 33507
rect 22569 33473 22603 33507
rect 24317 33473 24351 33507
rect 24777 33473 24811 33507
rect 25421 33473 25455 33507
rect 25973 33473 26007 33507
rect 27806 33473 27840 33507
rect 28641 33473 28675 33507
rect 28917 33473 28951 33507
rect 30297 33473 30331 33507
rect 30665 33473 30699 33507
rect 31125 33473 31159 33507
rect 31309 33473 31343 33507
rect 31401 33473 31435 33507
rect 31493 33473 31527 33507
rect 36481 33473 36515 33507
rect 39129 33473 39163 33507
rect 39497 33473 39531 33507
rect 40417 33473 40451 33507
rect 40510 33473 40544 33507
rect 40693 33473 40727 33507
rect 40923 33473 40957 33507
rect 5365 33405 5399 33439
rect 6653 33405 6687 33439
rect 6745 33405 6779 33439
rect 13645 33405 13679 33439
rect 19349 33405 19383 33439
rect 22477 33405 22511 33439
rect 25605 33405 25639 33439
rect 27629 33405 27663 33439
rect 28733 33405 28767 33439
rect 30205 33405 30239 33439
rect 36737 33405 36771 33439
rect 43085 33405 43119 33439
rect 43269 33405 43303 33439
rect 10793 33337 10827 33371
rect 20729 33337 20763 33371
rect 28457 33337 28491 33371
rect 39681 33337 39715 33371
rect 41061 33337 41095 33371
rect 4905 33269 4939 33303
rect 5273 33269 5307 33303
rect 8769 33269 8803 33303
rect 8953 33269 8987 33303
rect 9781 33269 9815 33303
rect 13369 33269 13403 33303
rect 13553 33269 13587 33303
rect 14289 33269 14323 33303
rect 18245 33269 18279 33303
rect 23121 33269 23155 33303
rect 27813 33269 27847 33303
rect 28641 33269 28675 33303
rect 30573 33269 30607 33303
rect 34437 33269 34471 33303
rect 35357 33269 35391 33303
rect 6285 33065 6319 33099
rect 7757 33065 7791 33099
rect 7849 33065 7883 33099
rect 7941 33065 7975 33099
rect 10793 33065 10827 33099
rect 10977 33065 11011 33099
rect 12265 33065 12299 33099
rect 17509 33065 17543 33099
rect 25789 33065 25823 33099
rect 27169 33065 27203 33099
rect 27353 33065 27387 33099
rect 28273 33065 28307 33099
rect 28733 33065 28767 33099
rect 38945 33065 38979 33099
rect 5457 32997 5491 33031
rect 25973 32997 26007 33031
rect 30481 32997 30515 33031
rect 6469 32929 6503 32963
rect 9137 32929 9171 32963
rect 9321 32929 9355 32963
rect 17969 32929 18003 32963
rect 18061 32929 18095 32963
rect 21005 32929 21039 32963
rect 22661 32929 22695 32963
rect 24593 32929 24627 32963
rect 25053 32929 25087 32963
rect 27077 32929 27111 32963
rect 34989 32929 35023 32963
rect 4077 32861 4111 32895
rect 4344 32861 4378 32895
rect 6561 32861 6595 32895
rect 6653 32861 6687 32895
rect 6745 32861 6779 32895
rect 8033 32861 8067 32895
rect 8217 32861 8251 32895
rect 9413 32861 9447 32895
rect 9505 32861 9539 32895
rect 9597 32861 9631 32895
rect 19625 32861 19659 32895
rect 19809 32861 19843 32895
rect 19993 32861 20027 32895
rect 21373 32861 21407 32895
rect 22042 32861 22076 32895
rect 22845 32861 22879 32895
rect 23029 32861 23063 32895
rect 23673 32861 23707 32895
rect 25145 32861 25179 32895
rect 26985 32861 27019 32895
rect 28457 32861 28491 32895
rect 28549 32861 28583 32895
rect 30297 32861 30331 32895
rect 30941 32861 30975 32895
rect 31217 32861 31251 32895
rect 33333 32861 33367 32895
rect 34069 32861 34103 32895
rect 35541 32861 35575 32895
rect 36093 32861 36127 32895
rect 36186 32861 36220 32895
rect 36558 32861 36592 32895
rect 37657 32861 37691 32895
rect 37805 32861 37839 32895
rect 38122 32861 38156 32895
rect 41429 32861 41463 32895
rect 42901 32861 42935 32895
rect 10609 32793 10643 32827
rect 12081 32793 12115 32827
rect 17877 32793 17911 32827
rect 19717 32793 19751 32827
rect 21281 32793 21315 32827
rect 26249 32793 26283 32827
rect 28273 32793 28307 32827
rect 36369 32793 36403 32827
rect 36461 32793 36495 32827
rect 37933 32793 37967 32827
rect 38025 32793 38059 32827
rect 38761 32793 38795 32827
rect 41162 32793 41196 32827
rect 43177 32793 43211 32827
rect 7481 32725 7515 32759
rect 10809 32725 10843 32759
rect 12281 32725 12315 32759
rect 12449 32725 12483 32759
rect 19441 32725 19475 32759
rect 21189 32725 21223 32759
rect 21557 32725 21591 32759
rect 24777 32725 24811 32759
rect 34069 32725 34103 32759
rect 36737 32725 36771 32759
rect 38301 32725 38335 32759
rect 38945 32725 38979 32759
rect 39129 32725 39163 32759
rect 40049 32725 40083 32759
rect 7113 32521 7147 32555
rect 7757 32521 7791 32555
rect 9229 32521 9263 32555
rect 11897 32521 11931 32555
rect 14381 32521 14415 32555
rect 20269 32521 20303 32555
rect 20637 32521 20671 32555
rect 26157 32521 26191 32555
rect 27261 32521 27295 32555
rect 29469 32521 29503 32555
rect 36921 32521 36955 32555
rect 39589 32521 39623 32555
rect 8677 32453 8711 32487
rect 9597 32453 9631 32487
rect 11713 32453 11747 32487
rect 13001 32453 13035 32487
rect 15086 32453 15120 32487
rect 28549 32453 28583 32487
rect 28733 32453 28767 32487
rect 32505 32453 32539 32487
rect 36553 32453 36587 32487
rect 36645 32453 36679 32487
rect 39037 32453 39071 32487
rect 4252 32385 4286 32419
rect 7297 32385 7331 32419
rect 7389 32385 7423 32419
rect 8585 32385 8619 32419
rect 8769 32385 8803 32419
rect 9413 32385 9447 32419
rect 12173 32385 12207 32419
rect 12817 32385 12851 32419
rect 13093 32385 13127 32419
rect 13185 32385 13219 32419
rect 13829 32385 13863 32419
rect 14013 32385 14047 32419
rect 14105 32385 14139 32419
rect 14197 32385 14231 32419
rect 18153 32385 18187 32419
rect 20453 32385 20487 32419
rect 20729 32385 20763 32419
rect 22845 32385 22879 32419
rect 23213 32385 23247 32419
rect 23397 32385 23431 32419
rect 23581 32385 23615 32419
rect 23857 32385 23891 32419
rect 25513 32385 25547 32419
rect 25697 32385 25731 32419
rect 26341 32385 26375 32419
rect 26525 32385 26559 32419
rect 26617 32385 26651 32419
rect 27445 32385 27479 32419
rect 27721 32385 27755 32419
rect 27905 32385 27939 32419
rect 28365 32385 28399 32419
rect 29285 32385 29319 32419
rect 29469 32385 29503 32419
rect 31125 32385 31159 32419
rect 31493 32385 31527 32419
rect 33517 32385 33551 32419
rect 34621 32385 34655 32419
rect 34989 32385 35023 32419
rect 35265 32385 35299 32419
rect 36277 32385 36311 32419
rect 36370 32385 36404 32419
rect 36742 32385 36776 32419
rect 38117 32385 38151 32419
rect 38761 32385 38795 32419
rect 38853 32385 38887 32419
rect 39497 32385 39531 32419
rect 39681 32385 39715 32419
rect 42993 32385 43027 32419
rect 3985 32317 4019 32351
rect 14841 32317 14875 32351
rect 18429 32317 18463 32351
rect 27629 32317 27663 32351
rect 30941 32317 30975 32351
rect 37749 32317 37783 32351
rect 38025 32317 38059 32351
rect 43085 32317 43119 32351
rect 43269 32317 43303 32351
rect 5365 32249 5399 32283
rect 25421 32249 25455 32283
rect 27537 32249 27571 32283
rect 39037 32249 39071 32283
rect 11897 32181 11931 32215
rect 13369 32181 13403 32215
rect 16221 32181 16255 32215
rect 19717 32181 19751 32215
rect 24225 32181 24259 32215
rect 42625 32181 42659 32215
rect 4629 31977 4663 32011
rect 10333 31977 10367 32011
rect 26893 31977 26927 32011
rect 32321 31977 32355 32011
rect 35909 31977 35943 32011
rect 37473 31977 37507 32011
rect 40969 31977 41003 32011
rect 13369 31909 13403 31943
rect 13461 31909 13495 31943
rect 15669 31909 15703 31943
rect 17785 31909 17819 31943
rect 23213 31909 23247 31943
rect 33517 31909 33551 31943
rect 42901 31909 42935 31943
rect 5273 31841 5307 31875
rect 10517 31841 10551 31875
rect 13185 31841 13219 31875
rect 14289 31841 14323 31875
rect 23397 31841 23431 31875
rect 28641 31841 28675 31875
rect 33379 31841 33413 31875
rect 37933 31841 37967 31875
rect 41521 31841 41555 31875
rect 5089 31773 5123 31807
rect 6101 31773 6135 31807
rect 6277 31751 6311 31785
rect 6377 31773 6411 31807
rect 6561 31773 6595 31807
rect 6653 31773 6687 31807
rect 7113 31773 7147 31807
rect 7297 31773 7331 31807
rect 9321 31773 9355 31807
rect 9505 31773 9539 31807
rect 9597 31773 9631 31807
rect 10333 31773 10367 31807
rect 10609 31773 10643 31807
rect 12357 31773 12391 31807
rect 13461 31773 13495 31807
rect 14556 31773 14590 31807
rect 16405 31773 16439 31807
rect 20269 31773 20303 31807
rect 20637 31773 20671 31807
rect 21097 31773 21131 31807
rect 21925 31773 21959 31807
rect 22017 31773 22051 31807
rect 23121 31773 23155 31807
rect 23305 31773 23339 31807
rect 23581 31773 23615 31807
rect 24961 31773 24995 31807
rect 25099 31773 25133 31807
rect 25329 31773 25363 31807
rect 26157 31773 26191 31807
rect 26801 31773 26835 31807
rect 26985 31773 27019 31807
rect 28273 31773 28307 31807
rect 28457 31773 28491 31807
rect 28549 31773 28583 31807
rect 28825 31773 28859 31807
rect 29745 31773 29779 31807
rect 29929 31773 29963 31807
rect 31309 31773 31343 31807
rect 32413 31773 32447 31807
rect 33241 31773 33275 31807
rect 33609 31773 33643 31807
rect 35265 31773 35299 31807
rect 35413 31773 35447 31807
rect 35541 31773 35575 31807
rect 35633 31773 35667 31807
rect 35730 31773 35764 31807
rect 36829 31773 36863 31807
rect 36922 31773 36956 31807
rect 37294 31773 37328 31807
rect 38301 31773 38335 31807
rect 38485 31773 38519 31807
rect 40325 31773 40359 31807
rect 40418 31773 40452 31807
rect 40831 31773 40865 31807
rect 41788 31773 41822 31807
rect 4997 31705 5031 31739
rect 7205 31705 7239 31739
rect 12449 31705 12483 31739
rect 16650 31705 16684 31739
rect 21741 31705 21775 31739
rect 25789 31705 25823 31739
rect 26341 31705 26375 31739
rect 37105 31705 37139 31739
rect 37197 31705 37231 31739
rect 40601 31705 40635 31739
rect 40693 31705 40727 31739
rect 9137 31637 9171 31671
rect 10793 31637 10827 31671
rect 22937 31637 22971 31671
rect 25237 31637 25271 31671
rect 29009 31637 29043 31671
rect 29837 31637 29871 31671
rect 6929 31433 6963 31467
rect 9413 31433 9447 31467
rect 9505 31433 9539 31467
rect 10793 31433 10827 31467
rect 34161 31433 34195 31467
rect 38485 31433 38519 31467
rect 41061 31433 41095 31467
rect 8677 31365 8711 31399
rect 11989 31365 12023 31399
rect 13737 31365 13771 31399
rect 13937 31365 13971 31399
rect 25697 31365 25731 31399
rect 32597 31365 32631 31399
rect 6837 31297 6871 31331
rect 7113 31297 7147 31331
rect 8217 31297 8251 31331
rect 8309 31297 8343 31331
rect 8493 31297 8527 31331
rect 9321 31297 9355 31331
rect 10149 31297 10183 31331
rect 10333 31297 10367 31331
rect 10425 31297 10459 31331
rect 10517 31297 10551 31331
rect 11713 31297 11747 31331
rect 12725 31297 12759 31331
rect 12909 31297 12943 31331
rect 19073 31297 19107 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 23949 31297 23983 31331
rect 25237 31297 25271 31331
rect 25329 31297 25363 31331
rect 26617 31297 26651 31331
rect 28089 31297 28123 31331
rect 28457 31297 28491 31331
rect 30849 31297 30883 31331
rect 31033 31297 31067 31331
rect 32413 31297 32447 31331
rect 33333 31297 33367 31331
rect 34253 31297 34287 31331
rect 35234 31297 35268 31331
rect 35357 31297 35391 31331
rect 36369 31297 36403 31331
rect 36461 31297 36495 31331
rect 36599 31297 36633 31331
rect 36737 31297 36771 31331
rect 37933 31297 37967 31331
rect 38117 31297 38151 31331
rect 38209 31297 38243 31331
rect 38301 31297 38335 31331
rect 40877 31297 40911 31331
rect 42901 31297 42935 31331
rect 23121 31229 23155 31263
rect 26433 31229 26467 31263
rect 27721 31229 27755 31263
rect 32781 31229 32815 31263
rect 35633 31229 35667 31263
rect 35725 31229 35759 31263
rect 43177 31229 43211 31263
rect 8401 31161 8435 31195
rect 9137 31161 9171 31195
rect 23213 31161 23247 31195
rect 23489 31161 23523 31195
rect 7297 31093 7331 31127
rect 9689 31093 9723 31127
rect 12725 31093 12759 31127
rect 13921 31093 13955 31127
rect 14105 31093 14139 31127
rect 19165 31093 19199 31127
rect 24041 31093 24075 31127
rect 25053 31093 25087 31127
rect 25237 31093 25271 31127
rect 31125 31093 31159 31127
rect 35081 31093 35115 31127
rect 36185 31093 36219 31127
rect 7021 30889 7055 30923
rect 7389 30889 7423 30923
rect 25053 30889 25087 30923
rect 43269 30889 43303 30923
rect 19717 30821 19751 30855
rect 24685 30821 24719 30855
rect 33057 30821 33091 30855
rect 33977 30821 34011 30855
rect 5457 30753 5491 30787
rect 7481 30753 7515 30787
rect 9689 30753 9723 30787
rect 9781 30753 9815 30787
rect 11621 30753 11655 30787
rect 17877 30753 17911 30787
rect 21373 30753 21407 30787
rect 23673 30753 23707 30787
rect 23857 30753 23891 30787
rect 25145 30753 25179 30787
rect 27629 30753 27663 30787
rect 27721 30753 27755 30787
rect 28457 30753 28491 30787
rect 35633 30753 35667 30787
rect 40049 30753 40083 30787
rect 40141 30753 40175 30787
rect 41889 30753 41923 30787
rect 5273 30685 5307 30719
rect 7205 30685 7239 30719
rect 8125 30685 8159 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 9873 30685 9907 30719
rect 9965 30685 9999 30719
rect 10609 30685 10643 30719
rect 10977 30685 11011 30719
rect 14565 30685 14599 30719
rect 17969 30685 18003 30719
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 20361 30685 20395 30719
rect 21005 30685 21039 30719
rect 24869 30685 24903 30719
rect 25881 30685 25915 30719
rect 26157 30685 26191 30719
rect 27353 30685 27387 30719
rect 28733 30685 28767 30719
rect 30665 30685 30699 30719
rect 31309 30685 31343 30719
rect 32965 30685 32999 30719
rect 33149 30685 33183 30719
rect 33241 30685 33275 30719
rect 34253 30685 34287 30719
rect 34897 30685 34931 30719
rect 34989 30685 35023 30719
rect 35173 30685 35207 30719
rect 36093 30685 36127 30719
rect 36185 30685 36219 30719
rect 36369 30685 36403 30719
rect 36461 30685 36495 30719
rect 37749 30685 37783 30719
rect 38761 30685 38795 30719
rect 38945 30685 38979 30719
rect 39129 30685 39163 30719
rect 40325 30685 40359 30719
rect 10793 30617 10827 30651
rect 10885 30617 10919 30651
rect 11866 30617 11900 30651
rect 14810 30617 14844 30651
rect 18245 30617 18279 30651
rect 18337 30617 18371 30651
rect 20821 30617 20855 30651
rect 27838 30617 27872 30651
rect 28825 30617 28859 30651
rect 29193 30617 29227 30651
rect 33977 30617 34011 30651
rect 37381 30617 37415 30651
rect 39037 30617 39071 30651
rect 42156 30617 42190 30651
rect 4813 30549 4847 30583
rect 5181 30549 5215 30583
rect 8585 30549 8619 30583
rect 9505 30549 9539 30583
rect 11161 30549 11195 30583
rect 13001 30549 13035 30583
rect 15945 30549 15979 30583
rect 17693 30549 17727 30583
rect 19533 30549 19567 30583
rect 20269 30549 20303 30583
rect 23213 30549 23247 30583
rect 23581 30549 23615 30583
rect 25697 30549 25731 30583
rect 27997 30549 28031 30583
rect 28641 30549 28675 30583
rect 31493 30549 31527 30583
rect 33425 30549 33459 30583
rect 34161 30549 34195 30583
rect 36645 30549 36679 30583
rect 39313 30549 39347 30583
rect 40509 30549 40543 30583
rect 5549 30345 5583 30379
rect 14565 30345 14599 30379
rect 20085 30345 20119 30379
rect 29469 30345 29503 30379
rect 30665 30345 30699 30379
rect 36001 30345 36035 30379
rect 42625 30345 42659 30379
rect 42993 30345 43027 30379
rect 43085 30345 43119 30379
rect 9505 30277 9539 30311
rect 14197 30277 14231 30311
rect 18889 30277 18923 30311
rect 39589 30277 39623 30311
rect 4169 30209 4203 30243
rect 4436 30209 4470 30243
rect 9597 30209 9631 30243
rect 10885 30209 10919 30243
rect 11069 30209 11103 30243
rect 11161 30209 11195 30243
rect 13001 30209 13035 30243
rect 13277 30209 13311 30243
rect 14013 30209 14047 30243
rect 14289 30209 14323 30243
rect 14381 30209 14415 30243
rect 17969 30209 18003 30243
rect 18797 30209 18831 30243
rect 19599 30209 19633 30243
rect 19717 30209 19751 30243
rect 19809 30209 19843 30243
rect 19901 30209 19935 30243
rect 21281 30209 21315 30243
rect 21465 30209 21499 30243
rect 22017 30209 22051 30243
rect 22273 30209 22307 30243
rect 24317 30209 24351 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 26341 30209 26375 30243
rect 26525 30209 26559 30243
rect 28089 30209 28123 30243
rect 28365 30209 28399 30243
rect 28733 30209 28767 30243
rect 29469 30209 29503 30243
rect 29653 30209 29687 30243
rect 30665 30209 30699 30243
rect 31309 30209 31343 30243
rect 32781 30209 32815 30243
rect 33609 30209 33643 30243
rect 34989 30209 35023 30243
rect 35449 30209 35483 30243
rect 35541 30209 35575 30243
rect 35725 30209 35759 30243
rect 35817 30209 35851 30243
rect 36461 30209 36495 30243
rect 37841 30209 37875 30243
rect 39037 30209 39071 30243
rect 39129 30209 39163 30243
rect 39313 30209 39347 30243
rect 39405 30209 39439 30243
rect 40325 30209 40359 30243
rect 40969 30209 41003 30243
rect 41153 30209 41187 30243
rect 17785 30141 17819 30175
rect 19441 30141 19475 30175
rect 21097 30141 21131 30175
rect 24409 30141 24443 30175
rect 24501 30141 24535 30175
rect 25697 30141 25731 30175
rect 31585 30141 31619 30175
rect 32321 30141 32355 30175
rect 33149 30141 33183 30175
rect 34253 30141 34287 30175
rect 36737 30141 36771 30175
rect 37933 30141 37967 30175
rect 38117 30141 38151 30175
rect 40141 30141 40175 30175
rect 40509 30141 40543 30175
rect 43177 30141 43211 30175
rect 23949 30073 23983 30107
rect 26341 30073 26375 30107
rect 10701 30005 10735 30039
rect 23397 30005 23431 30039
rect 27813 30005 27847 30039
rect 37473 30005 37507 30039
rect 41153 30005 41187 30039
rect 11621 29801 11655 29835
rect 18797 29801 18831 29835
rect 23581 29801 23615 29835
rect 32413 29801 32447 29835
rect 33609 29801 33643 29835
rect 36461 29801 36495 29835
rect 17877 29733 17911 29767
rect 16865 29665 16899 29699
rect 17417 29665 17451 29699
rect 19441 29665 19475 29699
rect 22937 29665 22971 29699
rect 23121 29665 23155 29699
rect 27537 29665 27571 29699
rect 30113 29665 30147 29699
rect 30389 29665 30423 29699
rect 30573 29665 30607 29699
rect 41981 29665 42015 29699
rect 6837 29597 6871 29631
rect 6929 29597 6963 29631
rect 7205 29597 7239 29631
rect 7941 29597 7975 29631
rect 8033 29597 8067 29631
rect 10241 29597 10275 29631
rect 12633 29597 12667 29631
rect 12817 29597 12851 29631
rect 17601 29597 17635 29631
rect 17693 29597 17727 29631
rect 17969 29597 18003 29631
rect 18705 29597 18739 29631
rect 18797 29597 18831 29631
rect 19717 29597 19751 29631
rect 19809 29597 19843 29631
rect 19901 29597 19935 29631
rect 20085 29597 20119 29631
rect 20545 29597 20579 29631
rect 20729 29597 20763 29631
rect 26617 29597 26651 29631
rect 26985 29597 27019 29631
rect 27997 29597 28031 29631
rect 28641 29597 28675 29631
rect 30665 29597 30699 29631
rect 31493 29597 31527 29631
rect 31677 29597 31711 29631
rect 31861 29597 31895 29631
rect 32321 29597 32355 29631
rect 32965 29597 32999 29631
rect 33113 29597 33147 29631
rect 33333 29597 33367 29631
rect 33449 29597 33483 29631
rect 34897 29597 34931 29631
rect 34989 29597 35023 29631
rect 35173 29597 35207 29631
rect 37841 29597 37875 29631
rect 41714 29597 41748 29631
rect 42901 29597 42935 29631
rect 7021 29529 7055 29563
rect 10508 29529 10542 29563
rect 19599 29529 19633 29563
rect 26433 29529 26467 29563
rect 27629 29529 27663 29563
rect 31585 29529 31619 29563
rect 33241 29529 33275 29563
rect 35633 29529 35667 29563
rect 37574 29529 37608 29563
rect 43177 29529 43211 29563
rect 6653 29461 6687 29495
rect 7757 29461 7791 29495
rect 12725 29461 12759 29495
rect 16221 29461 16255 29495
rect 16589 29461 16623 29495
rect 16681 29461 16715 29495
rect 18429 29461 18463 29495
rect 20637 29461 20671 29495
rect 23213 29461 23247 29495
rect 28733 29461 28767 29495
rect 31309 29461 31343 29495
rect 40601 29461 40635 29495
rect 9045 29257 9079 29291
rect 16865 29257 16899 29291
rect 18061 29257 18095 29291
rect 25697 29257 25731 29291
rect 27721 29257 27755 29291
rect 28457 29257 28491 29291
rect 32965 29257 32999 29291
rect 39589 29257 39623 29291
rect 41061 29257 41095 29291
rect 17233 29189 17267 29223
rect 28365 29189 28399 29223
rect 29929 29189 29963 29223
rect 30113 29189 30147 29223
rect 32873 29189 32907 29223
rect 34621 29189 34655 29223
rect 35633 29189 35667 29223
rect 38209 29189 38243 29223
rect 40417 29189 40451 29223
rect 40877 29189 40911 29223
rect 7665 29121 7699 29155
rect 7932 29121 7966 29155
rect 13369 29121 13403 29155
rect 13636 29121 13670 29155
rect 18245 29121 18279 29155
rect 18521 29121 18555 29155
rect 19441 29121 19475 29155
rect 19625 29121 19659 29155
rect 25329 29121 25363 29155
rect 27629 29121 27663 29155
rect 27813 29121 27847 29155
rect 28641 29121 28675 29155
rect 29745 29121 29779 29155
rect 31033 29121 31067 29155
rect 33149 29121 33183 29155
rect 34437 29121 34471 29155
rect 34713 29121 34747 29155
rect 34805 29121 34839 29155
rect 36369 29121 36403 29155
rect 37473 29121 37507 29155
rect 37703 29121 37737 29155
rect 38945 29121 38979 29155
rect 39093 29121 39127 29155
rect 39221 29121 39255 29155
rect 39313 29121 39347 29155
rect 39410 29121 39444 29155
rect 40141 29121 40175 29155
rect 40325 29121 40359 29155
rect 41153 29121 41187 29155
rect 17325 29053 17359 29087
rect 17417 29053 17451 29087
rect 18337 29053 18371 29087
rect 19257 29053 19291 29087
rect 25421 29053 25455 29087
rect 28733 29053 28767 29087
rect 30849 29053 30883 29087
rect 33333 29053 33367 29087
rect 37841 29053 37875 29087
rect 14749 28985 14783 29019
rect 34989 28985 35023 29019
rect 40877 28985 40911 29019
rect 18521 28917 18555 28951
rect 28549 28917 28583 28951
rect 37611 28917 37645 28951
rect 8033 28713 8067 28747
rect 13737 28713 13771 28747
rect 20913 28713 20947 28747
rect 22845 28713 22879 28747
rect 32781 28713 32815 28747
rect 43269 28713 43303 28747
rect 6929 28645 6963 28679
rect 16865 28645 16899 28679
rect 28089 28645 28123 28679
rect 30481 28645 30515 28679
rect 39497 28645 39531 28679
rect 18429 28577 18463 28611
rect 33149 28577 33183 28611
rect 40141 28577 40175 28611
rect 5549 28509 5583 28543
rect 8217 28509 8251 28543
rect 8309 28509 8343 28543
rect 8585 28509 8619 28543
rect 9137 28509 9171 28543
rect 9404 28509 9438 28543
rect 13185 28509 13219 28543
rect 13461 28509 13495 28543
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 14657 28509 14691 28543
rect 15485 28509 15519 28543
rect 19901 28509 19935 28543
rect 22845 28509 22879 28543
rect 22937 28509 22971 28543
rect 24869 28509 24903 28543
rect 26801 28509 26835 28543
rect 27997 28509 28031 28543
rect 28549 28509 28583 28543
rect 28733 28509 28767 28543
rect 30205 28509 30239 28543
rect 30481 28509 30515 28543
rect 31309 28509 31343 28543
rect 31493 28509 31527 28543
rect 31677 28509 31711 28543
rect 32965 28509 32999 28543
rect 33241 28509 33275 28543
rect 34897 28509 34931 28543
rect 34989 28509 35023 28543
rect 35173 28509 35207 28543
rect 35633 28509 35667 28543
rect 36921 28509 36955 28543
rect 37197 28509 37231 28543
rect 37381 28509 37415 28543
rect 37565 28509 37599 28543
rect 38853 28509 38887 28543
rect 38946 28509 38980 28543
rect 39221 28509 39255 28543
rect 39318 28509 39352 28543
rect 40049 28509 40083 28543
rect 40325 28509 40359 28543
rect 40417 28509 40451 28543
rect 41889 28509 41923 28543
rect 5816 28441 5850 28475
rect 8401 28441 8435 28475
rect 13369 28441 13403 28475
rect 14473 28441 14507 28475
rect 15752 28441 15786 28475
rect 19993 28441 20027 28475
rect 20361 28441 20395 28475
rect 23121 28441 23155 28475
rect 25114 28441 25148 28475
rect 27169 28441 27203 28475
rect 31401 28441 31435 28475
rect 39129 28441 39163 28475
rect 42156 28441 42190 28475
rect 10517 28373 10551 28407
rect 14841 28373 14875 28407
rect 17785 28373 17819 28407
rect 18153 28373 18187 28407
rect 18245 28373 18279 28407
rect 19625 28373 19659 28407
rect 20729 28373 20763 28407
rect 22661 28373 22695 28407
rect 26249 28373 26283 28407
rect 30297 28373 30331 28407
rect 31125 28373 31159 28407
rect 37473 28373 37507 28407
rect 40601 28373 40635 28407
rect 7021 28169 7055 28203
rect 17325 28169 17359 28203
rect 17693 28169 17727 28203
rect 21189 28169 21223 28203
rect 22845 28169 22879 28203
rect 23213 28169 23247 28203
rect 24225 28169 24259 28203
rect 38117 28169 38151 28203
rect 42625 28169 42659 28203
rect 42993 28169 43027 28203
rect 43085 28169 43119 28203
rect 12265 28101 12299 28135
rect 14942 28101 14976 28135
rect 26525 28101 26559 28135
rect 31033 28101 31067 28135
rect 32689 28101 32723 28135
rect 33517 28101 33551 28135
rect 36829 28101 36863 28135
rect 37473 28101 37507 28135
rect 39221 28101 39255 28135
rect 6929 28033 6963 28067
rect 8125 28033 8159 28067
rect 8309 28033 8343 28067
rect 11989 28033 12023 28067
rect 12173 28033 12207 28067
rect 12357 28033 12391 28067
rect 15209 28033 15243 28067
rect 21097 28033 21131 28067
rect 24593 28033 24627 28067
rect 26157 28033 26191 28067
rect 26341 28033 26375 28067
rect 28181 28033 28215 28067
rect 30849 28033 30883 28067
rect 30941 28033 30975 28067
rect 31217 28033 31251 28067
rect 32459 28033 32493 28067
rect 32597 28033 32631 28067
rect 32873 28033 32907 28067
rect 33333 28033 33367 28067
rect 33609 28033 33643 28067
rect 34253 28033 34287 28067
rect 34989 28033 35023 28067
rect 35173 28033 35207 28067
rect 36001 28033 36035 28067
rect 37841 28033 37875 28067
rect 39497 28033 39531 28067
rect 7205 27965 7239 27999
rect 17785 27965 17819 27999
rect 17969 27965 18003 27999
rect 21373 27965 21407 27999
rect 23305 27965 23339 27999
rect 23397 27965 23431 27999
rect 24041 27965 24075 27999
rect 24501 27965 24535 27999
rect 28365 27965 28399 27999
rect 28457 27965 28491 27999
rect 28549 27965 28583 27999
rect 28641 27965 28675 27999
rect 35265 27965 35299 27999
rect 37565 27965 37599 27999
rect 37933 27965 37967 27999
rect 43269 27965 43303 27999
rect 13829 27897 13863 27931
rect 6561 27829 6595 27863
rect 8217 27829 8251 27863
rect 12541 27829 12575 27863
rect 20729 27829 20763 27863
rect 28825 27829 28859 27863
rect 30665 27829 30699 27863
rect 32321 27829 32355 27863
rect 33333 27829 33367 27863
rect 25973 27625 26007 27659
rect 17693 27557 17727 27591
rect 23489 27557 23523 27591
rect 27169 27557 27203 27591
rect 32505 27557 32539 27591
rect 40233 27557 40267 27591
rect 7941 27489 7975 27523
rect 11713 27489 11747 27523
rect 25881 27489 25915 27523
rect 37933 27489 37967 27523
rect 43177 27489 43211 27523
rect 5273 27421 5307 27455
rect 8033 27421 8067 27455
rect 8309 27421 8343 27455
rect 9781 27421 9815 27455
rect 16589 27421 16623 27455
rect 17601 27421 17635 27455
rect 20637 27421 20671 27455
rect 20904 27421 20938 27455
rect 23213 27421 23247 27455
rect 23305 27421 23339 27455
rect 23581 27421 23615 27455
rect 24593 27421 24627 27455
rect 24777 27421 24811 27455
rect 25053 27421 25087 27455
rect 25973 27421 26007 27455
rect 27301 27421 27335 27455
rect 27445 27421 27479 27455
rect 27537 27421 27571 27455
rect 27721 27421 27755 27455
rect 29883 27421 29917 27455
rect 30021 27421 30055 27455
rect 30297 27421 30331 27455
rect 30941 27421 30975 27455
rect 31125 27421 31159 27455
rect 32689 27421 32723 27455
rect 32781 27421 32815 27455
rect 33057 27421 33091 27455
rect 34989 27421 35023 27455
rect 35081 27421 35115 27455
rect 35265 27421 35299 27455
rect 35357 27421 35391 27455
rect 36093 27421 36127 27455
rect 36369 27421 36403 27455
rect 36461 27421 36495 27455
rect 37105 27421 37139 27455
rect 38669 27421 38703 27455
rect 38761 27421 38795 27455
rect 39037 27421 39071 27455
rect 40417 27421 40451 27455
rect 42901 27421 42935 27455
rect 5540 27353 5574 27387
rect 8401 27353 8435 27387
rect 10048 27353 10082 27387
rect 11980 27353 12014 27387
rect 25697 27353 25731 27387
rect 30113 27353 30147 27387
rect 32873 27353 32907 27387
rect 36277 27353 36311 27387
rect 38853 27353 38887 27387
rect 40601 27353 40635 27387
rect 6653 27285 6687 27319
rect 7757 27285 7791 27319
rect 11161 27285 11195 27319
rect 13093 27285 13127 27319
rect 16681 27285 16715 27319
rect 22017 27285 22051 27319
rect 23029 27285 23063 27319
rect 25237 27285 25271 27319
rect 26157 27285 26191 27319
rect 29745 27285 29779 27319
rect 31033 27285 31067 27319
rect 35541 27285 35575 27319
rect 36645 27285 36679 27319
rect 38485 27285 38519 27319
rect 10333 27081 10367 27115
rect 10701 27081 10735 27115
rect 10793 27081 10827 27115
rect 13461 27081 13495 27115
rect 17233 27081 17267 27115
rect 22017 27081 22051 27115
rect 23213 27081 23247 27115
rect 25053 27081 25087 27115
rect 25789 27081 25823 27115
rect 26249 27081 26283 27115
rect 28365 27081 28399 27115
rect 36093 27081 36127 27115
rect 12348 27013 12382 27047
rect 24961 27013 24995 27047
rect 28733 27013 28767 27047
rect 30205 27013 30239 27047
rect 36737 27013 36771 27047
rect 37473 27013 37507 27047
rect 7205 26945 7239 26979
rect 7472 26945 7506 26979
rect 9045 26945 9079 26979
rect 9229 26945 9263 26979
rect 12081 26945 12115 26979
rect 15853 26945 15887 26979
rect 16129 26945 16163 26979
rect 18061 26945 18095 26979
rect 18245 26945 18279 26979
rect 19349 26945 19383 26979
rect 19809 26945 19843 26979
rect 21097 26945 21131 26979
rect 21189 26945 21223 26979
rect 21373 26945 21407 26979
rect 21465 26945 21499 26979
rect 22201 26945 22235 26979
rect 23397 26945 23431 26979
rect 23581 26945 23615 26979
rect 26157 26945 26191 26979
rect 28549 26945 28583 26979
rect 28825 26945 28859 26979
rect 29285 26945 29319 26979
rect 29377 26945 29411 26979
rect 29469 26945 29503 26979
rect 30849 26945 30883 26979
rect 30941 26945 30975 26979
rect 31217 26945 31251 26979
rect 32873 26945 32907 26979
rect 33057 26945 33091 26979
rect 34161 26945 34195 26979
rect 34345 26945 34379 26979
rect 36369 26945 36403 26979
rect 38853 26945 38887 26979
rect 39001 26945 39035 26979
rect 39129 26945 39163 26979
rect 39221 26945 39255 26979
rect 39318 26945 39352 26979
rect 41806 26945 41840 26979
rect 42073 26945 42107 26979
rect 42993 26945 43027 26979
rect 10885 26877 10919 26911
rect 15945 26877 15979 26911
rect 17325 26877 17359 26911
rect 17417 26877 17451 26911
rect 20913 26877 20947 26911
rect 22385 26877 22419 26911
rect 22477 26877 22511 26911
rect 23673 26877 23707 26911
rect 25237 26877 25271 26911
rect 26341 26877 26375 26911
rect 31309 26877 31343 26911
rect 36277 26877 36311 26911
rect 36645 26877 36679 26911
rect 38209 26877 38243 26911
rect 43085 26877 43119 26911
rect 43269 26877 43303 26911
rect 8585 26809 8619 26843
rect 16313 26809 16347 26843
rect 19533 26809 19567 26843
rect 9229 26741 9263 26775
rect 15853 26741 15887 26775
rect 16865 26741 16899 26775
rect 18061 26741 18095 26775
rect 19073 26741 19107 26775
rect 19441 26741 19475 26775
rect 19625 26741 19659 26775
rect 24593 26741 24627 26775
rect 33057 26741 33091 26775
rect 34069 26741 34103 26775
rect 39497 26741 39531 26775
rect 40693 26741 40727 26775
rect 42625 26741 42659 26775
rect 12173 26537 12207 26571
rect 24869 26537 24903 26571
rect 32597 26537 32631 26571
rect 34989 26537 35023 26571
rect 40785 26537 40819 26571
rect 43361 26537 43395 26571
rect 9137 26469 9171 26503
rect 14381 26469 14415 26503
rect 18337 26469 18371 26503
rect 27629 26469 27663 26503
rect 29745 26469 29779 26503
rect 34345 26469 34379 26503
rect 10977 26401 11011 26435
rect 16957 26401 16991 26435
rect 23489 26401 23523 26435
rect 27721 26401 27755 26435
rect 40325 26401 40359 26435
rect 41981 26401 42015 26435
rect 9321 26333 9355 26367
rect 9505 26333 9539 26367
rect 9689 26333 9723 26367
rect 12357 26333 12391 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 15761 26333 15795 26367
rect 17141 26333 17175 26367
rect 18153 26333 18187 26367
rect 18429 26333 18463 26367
rect 19441 26333 19475 26367
rect 23305 26333 23339 26367
rect 23397 26333 23431 26367
rect 26341 26333 26375 26367
rect 27169 26333 27203 26367
rect 27353 26333 27387 26367
rect 28181 26333 28215 26367
rect 28365 26333 28399 26367
rect 28733 26333 28767 26367
rect 29745 26333 29779 26367
rect 30021 26333 30055 26367
rect 31217 26333 31251 26367
rect 31493 26333 31527 26367
rect 32776 26333 32810 26367
rect 32873 26333 32907 26367
rect 33148 26333 33182 26367
rect 33241 26333 33275 26367
rect 33793 26333 33827 26367
rect 33977 26333 34011 26367
rect 34161 26333 34195 26367
rect 34897 26333 34931 26367
rect 35173 26333 35207 26367
rect 36507 26333 36541 26367
rect 36645 26333 36679 26367
rect 36737 26333 36771 26367
rect 36865 26333 36899 26367
rect 37013 26333 37047 26367
rect 37565 26333 37599 26367
rect 37933 26333 37967 26367
rect 38025 26333 38059 26367
rect 38669 26333 38703 26367
rect 38817 26333 38851 26367
rect 39175 26333 39209 26367
rect 40417 26333 40451 26367
rect 42248 26333 42282 26367
rect 9413 26265 9447 26299
rect 11713 26265 11747 26299
rect 12449 26265 12483 26299
rect 15516 26265 15550 26299
rect 17049 26265 17083 26299
rect 17969 26265 18003 26299
rect 19686 26265 19720 26299
rect 29929 26265 29963 26299
rect 31033 26265 31067 26299
rect 31401 26265 31435 26299
rect 32965 26265 32999 26299
rect 34069 26265 34103 26299
rect 35357 26265 35391 26299
rect 37657 26265 37691 26299
rect 38945 26265 38979 26299
rect 39037 26265 39071 26299
rect 17509 26197 17543 26231
rect 20821 26197 20855 26231
rect 22937 26197 22971 26231
rect 28641 26197 28675 26231
rect 36369 26197 36403 26231
rect 38209 26197 38243 26231
rect 39313 26197 39347 26231
rect 15853 25993 15887 26027
rect 19533 25993 19567 26027
rect 25237 25993 25271 26027
rect 27261 25993 27295 26027
rect 28365 25993 28399 26027
rect 32781 25993 32815 26027
rect 36645 25993 36679 26027
rect 40049 25993 40083 26027
rect 12633 25925 12667 25959
rect 17417 25925 17451 25959
rect 18153 25925 18187 25959
rect 19165 25925 19199 25959
rect 22836 25925 22870 25959
rect 30757 25925 30791 25959
rect 31493 25925 31527 25959
rect 33057 25925 33091 25959
rect 33149 25925 33183 25959
rect 35265 25925 35299 25959
rect 39865 25925 39899 25959
rect 43177 25925 43211 25959
rect 15485 25857 15519 25891
rect 19993 25857 20027 25891
rect 20177 25857 20211 25891
rect 22569 25857 22603 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 25973 25857 26007 25891
rect 26249 25857 26283 25891
rect 26433 25857 26467 25891
rect 27175 25857 27209 25891
rect 27365 25857 27399 25891
rect 27997 25857 28031 25891
rect 32919 25857 32953 25891
rect 33277 25857 33311 25891
rect 33425 25857 33459 25891
rect 34529 25857 34563 25891
rect 34989 25857 35023 25891
rect 36185 25857 36219 25891
rect 36647 25857 36681 25891
rect 38761 25857 38795 25891
rect 39037 25857 39071 25891
rect 39129 25857 39163 25891
rect 40141 25857 40175 25891
rect 42901 25857 42935 25891
rect 11897 25789 11931 25823
rect 15301 25789 15335 25823
rect 15393 25789 15427 25823
rect 18981 25789 19015 25823
rect 19073 25789 19107 25823
rect 28089 25789 28123 25823
rect 31125 25789 31159 25823
rect 39313 25789 39347 25823
rect 31217 25721 31251 25755
rect 36277 25721 36311 25755
rect 39865 25721 39899 25755
rect 20361 25653 20395 25687
rect 23949 25653 23983 25687
rect 31328 25653 31362 25687
rect 36829 25653 36863 25687
rect 38853 25653 38887 25687
rect 11069 25449 11103 25483
rect 18337 25449 18371 25483
rect 18705 25449 18739 25483
rect 25513 25449 25547 25483
rect 25973 25449 26007 25483
rect 32873 25449 32907 25483
rect 36553 25449 36587 25483
rect 40693 25449 40727 25483
rect 12265 25381 12299 25415
rect 17785 25381 17819 25415
rect 26985 25381 27019 25415
rect 30021 25381 30055 25415
rect 31861 25381 31895 25415
rect 13185 25313 13219 25347
rect 20637 25313 20671 25347
rect 36645 25313 36679 25347
rect 37565 25313 37599 25347
rect 39037 25313 39071 25347
rect 9689 25245 9723 25279
rect 11838 25245 11872 25279
rect 12357 25245 12391 25279
rect 13001 25245 13035 25279
rect 13277 25245 13311 25279
rect 14841 25245 14875 25279
rect 15025 25245 15059 25279
rect 15209 25245 15243 25279
rect 17141 25245 17175 25279
rect 17234 25245 17268 25279
rect 17606 25245 17640 25279
rect 18245 25245 18279 25279
rect 18521 25245 18555 25279
rect 20893 25245 20927 25279
rect 25697 25245 25731 25279
rect 25789 25245 25823 25279
rect 27117 25245 27151 25279
rect 27353 25245 27387 25279
rect 27537 25245 27571 25279
rect 29745 25245 29779 25279
rect 30941 25245 30975 25279
rect 31585 25245 31619 25279
rect 31861 25245 31895 25279
rect 32689 25245 32723 25279
rect 32873 25245 32907 25279
rect 35449 25245 35483 25279
rect 35597 25245 35631 25279
rect 35914 25245 35948 25279
rect 36553 25245 36587 25279
rect 37473 25245 37507 25279
rect 37657 25245 37691 25279
rect 38945 25245 38979 25279
rect 39221 25245 39255 25279
rect 39313 25245 39347 25279
rect 39497 25245 39531 25279
rect 42901 25245 42935 25279
rect 9956 25177 9990 25211
rect 14933 25177 14967 25211
rect 17417 25177 17451 25211
rect 17509 25177 17543 25211
rect 25513 25177 25547 25211
rect 27261 25177 27295 25211
rect 30021 25177 30055 25211
rect 30665 25177 30699 25211
rect 35725 25177 35759 25211
rect 35817 25177 35851 25211
rect 40325 25177 40359 25211
rect 40509 25177 40543 25211
rect 43177 25177 43211 25211
rect 11713 25109 11747 25143
rect 11897 25109 11931 25143
rect 12817 25109 12851 25143
rect 14657 25109 14691 25143
rect 22017 25109 22051 25143
rect 29837 25109 29871 25143
rect 31677 25109 31711 25143
rect 36093 25109 36127 25143
rect 36921 25109 36955 25143
rect 10241 24905 10275 24939
rect 10609 24905 10643 24939
rect 39221 24905 39255 24939
rect 43085 24905 43119 24939
rect 12808 24837 12842 24871
rect 17785 24837 17819 24871
rect 32689 24837 32723 24871
rect 9054 24769 9088 24803
rect 10701 24769 10735 24803
rect 14740 24769 14774 24803
rect 19717 24769 19751 24803
rect 22385 24769 22419 24803
rect 22477 24769 22511 24803
rect 23213 24769 23247 24803
rect 23673 24769 23707 24803
rect 23765 24769 23799 24803
rect 23949 24769 23983 24803
rect 24777 24769 24811 24803
rect 25053 24769 25087 24803
rect 25881 24769 25915 24803
rect 28457 24769 28491 24803
rect 28641 24769 28675 24803
rect 29101 24769 29135 24803
rect 30389 24769 30423 24803
rect 30757 24769 30791 24803
rect 30869 24769 30903 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 32873 24769 32907 24803
rect 36277 24769 36311 24803
rect 36370 24769 36404 24803
rect 36553 24769 36587 24803
rect 36645 24769 36679 24803
rect 36742 24769 36776 24803
rect 38577 24769 38611 24803
rect 38725 24769 38759 24803
rect 38853 24769 38887 24803
rect 38945 24769 38979 24803
rect 39083 24769 39117 24803
rect 39681 24769 39715 24803
rect 39865 24769 39899 24803
rect 39957 24769 39991 24803
rect 41806 24769 41840 24803
rect 42073 24769 42107 24803
rect 42993 24769 43027 24803
rect 9321 24701 9355 24735
rect 10885 24701 10919 24735
rect 12541 24701 12575 24735
rect 14473 24701 14507 24735
rect 16957 24701 16991 24735
rect 19901 24701 19935 24735
rect 24961 24701 24995 24735
rect 29285 24701 29319 24735
rect 29377 24701 29411 24735
rect 29745 24701 29779 24735
rect 30481 24701 30515 24735
rect 43269 24701 43303 24735
rect 23121 24633 23155 24667
rect 28549 24633 28583 24667
rect 39681 24633 39715 24667
rect 7941 24565 7975 24599
rect 13921 24565 13955 24599
rect 15853 24565 15887 24599
rect 19533 24565 19567 24599
rect 24133 24565 24167 24599
rect 31033 24565 31067 24599
rect 32321 24565 32355 24599
rect 36921 24565 36955 24599
rect 40693 24565 40727 24599
rect 42625 24565 42659 24599
rect 14933 24361 14967 24395
rect 28457 24361 28491 24395
rect 28825 24361 28859 24395
rect 30481 24361 30515 24395
rect 38209 24361 38243 24395
rect 39497 24361 39531 24395
rect 40785 24361 40819 24395
rect 43361 24361 43395 24395
rect 23213 24293 23247 24327
rect 26893 24293 26927 24327
rect 10333 24225 10367 24259
rect 10517 24225 10551 24259
rect 14657 24225 14691 24259
rect 17325 24225 17359 24259
rect 30297 24225 30331 24259
rect 34345 24225 34379 24259
rect 37565 24225 37599 24259
rect 38025 24225 38059 24259
rect 40325 24225 40359 24259
rect 41981 24225 42015 24259
rect 11345 24157 11379 24191
rect 14749 24157 14783 24191
rect 17049 24157 17083 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 21741 24157 21775 24191
rect 22661 24157 22695 24191
rect 22845 24157 22879 24191
rect 23489 24157 23523 24191
rect 24593 24157 24627 24191
rect 24777 24157 24811 24191
rect 27072 24157 27106 24191
rect 27169 24157 27203 24191
rect 27261 24157 27295 24191
rect 27445 24157 27479 24191
rect 28365 24157 28399 24191
rect 28641 24157 28675 24191
rect 30021 24157 30055 24191
rect 30113 24157 30147 24191
rect 30205 24157 30239 24191
rect 31309 24157 31343 24191
rect 32873 24157 32907 24191
rect 33241 24157 33275 24191
rect 33977 24157 34011 24191
rect 34253 24157 34287 24191
rect 37933 24157 37967 24191
rect 38853 24157 38887 24191
rect 38946 24157 38980 24191
rect 39083 24157 39117 24191
rect 39359 24157 39393 24191
rect 40417 24157 40451 24191
rect 42248 24157 42282 24191
rect 11612 24089 11646 24123
rect 18705 24089 18739 24123
rect 30941 24089 30975 24123
rect 31125 24089 31159 24123
rect 37657 24089 37691 24123
rect 39218 24089 39252 24123
rect 9873 24021 9907 24055
rect 10241 24021 10275 24055
rect 12725 24021 12759 24055
rect 20177 24021 20211 24055
rect 21465 24021 21499 24055
rect 24685 24021 24719 24055
rect 24409 23817 24443 23851
rect 24501 23817 24535 23851
rect 27369 23817 27403 23851
rect 28089 23817 28123 23851
rect 31677 23817 31711 23851
rect 21189 23749 21223 23783
rect 22477 23749 22511 23783
rect 24685 23749 24719 23783
rect 25605 23749 25639 23783
rect 27169 23749 27203 23783
rect 32965 23749 32999 23783
rect 35173 23749 35207 23783
rect 9229 23681 9263 23715
rect 9496 23681 9530 23715
rect 15025 23681 15059 23715
rect 15209 23681 15243 23715
rect 15761 23681 15795 23715
rect 15853 23681 15887 23715
rect 19901 23681 19935 23715
rect 19993 23681 20027 23715
rect 20085 23681 20119 23715
rect 20269 23681 20303 23715
rect 21097 23681 21131 23715
rect 23489 23681 23523 23715
rect 24317 23681 24351 23715
rect 27997 23681 28031 23715
rect 28181 23681 28215 23715
rect 28825 23681 28859 23715
rect 28917 23681 28951 23715
rect 30021 23681 30055 23715
rect 30389 23681 30423 23715
rect 31527 23681 31561 23715
rect 32597 23681 32631 23715
rect 32690 23681 32724 23715
rect 32873 23681 32907 23715
rect 33103 23681 33137 23715
rect 34069 23681 34103 23715
rect 34621 23681 34655 23715
rect 34989 23681 35023 23715
rect 36553 23681 36587 23715
rect 36737 23681 36771 23715
rect 42901 23681 42935 23715
rect 15301 23613 15335 23647
rect 16313 23613 16347 23647
rect 21373 23613 21407 23647
rect 22017 23613 22051 23647
rect 31125 23613 31159 23647
rect 31217 23613 31251 23647
rect 43177 23613 43211 23647
rect 10609 23545 10643 23579
rect 20729 23545 20763 23579
rect 22201 23545 22235 23579
rect 24133 23545 24167 23579
rect 25329 23545 25363 23579
rect 29193 23545 29227 23579
rect 30573 23545 30607 23579
rect 19625 23477 19659 23511
rect 23581 23477 23615 23511
rect 25145 23477 25179 23511
rect 27353 23477 27387 23511
rect 27537 23477 27571 23511
rect 28917 23477 28951 23511
rect 30113 23477 30147 23511
rect 33241 23477 33275 23511
rect 36645 23477 36679 23511
rect 17325 23273 17359 23307
rect 24593 23273 24627 23307
rect 18889 23205 18923 23239
rect 23397 23205 23431 23239
rect 34069 23205 34103 23239
rect 37749 23205 37783 23239
rect 39497 23205 39531 23239
rect 10701 23137 10735 23171
rect 15761 23137 15795 23171
rect 19993 23137 20027 23171
rect 21005 23137 21039 23171
rect 22385 23137 22419 23171
rect 23213 23137 23247 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 27445 23137 27479 23171
rect 27537 23137 27571 23171
rect 36553 23137 36587 23171
rect 38117 23137 38151 23171
rect 40141 23137 40175 23171
rect 40601 23137 40635 23171
rect 42717 23137 42751 23171
rect 42901 23137 42935 23171
rect 16037 23069 16071 23103
rect 18613 23069 18647 23103
rect 20085 23069 20119 23103
rect 21189 23069 21223 23103
rect 21281 23069 21315 23103
rect 22477 23069 22511 23103
rect 22569 23069 22603 23103
rect 22661 23069 22695 23103
rect 23489 23069 23523 23103
rect 24961 23069 24995 23103
rect 26157 23069 26191 23103
rect 27169 23069 27203 23103
rect 30297 23071 30331 23105
rect 33517 23069 33551 23103
rect 33701 23069 33735 23103
rect 33885 23069 33919 23103
rect 35633 23069 35667 23103
rect 35725 23069 35759 23103
rect 35817 23069 35851 23103
rect 35909 23069 35943 23103
rect 36461 23069 36495 23103
rect 36737 23069 36771 23103
rect 36829 23069 36863 23103
rect 37657 23069 37691 23103
rect 37841 23069 37875 23103
rect 37933 23069 37967 23103
rect 38853 23069 38887 23103
rect 39001 23069 39035 23103
rect 39359 23069 39393 23103
rect 40049 23069 40083 23103
rect 40325 23069 40359 23103
rect 40417 23069 40451 23103
rect 10968 23001 11002 23035
rect 18889 23001 18923 23035
rect 21649 23001 21683 23035
rect 23213 23001 23247 23035
rect 25789 23001 25823 23035
rect 25973 23001 26007 23035
rect 33793 23001 33827 23035
rect 39129 23001 39163 23035
rect 39221 23001 39255 23035
rect 12081 22933 12115 22967
rect 18705 22933 18739 22967
rect 19809 22933 19843 22967
rect 20453 22933 20487 22967
rect 22201 22933 22235 22967
rect 30389 22933 30423 22967
rect 35449 22933 35483 22967
rect 37013 22933 37047 22967
rect 42257 22933 42291 22967
rect 42625 22933 42659 22967
rect 13921 22729 13955 22763
rect 16957 22729 16991 22763
rect 18337 22729 18371 22763
rect 20361 22729 20395 22763
rect 23673 22729 23707 22763
rect 24685 22729 24719 22763
rect 28565 22729 28599 22763
rect 35633 22729 35667 22763
rect 36185 22729 36219 22763
rect 38117 22729 38151 22763
rect 17141 22661 17175 22695
rect 27629 22661 27663 22695
rect 28365 22661 28399 22695
rect 33885 22661 33919 22695
rect 35265 22661 35299 22695
rect 37565 22661 37599 22695
rect 39313 22661 39347 22695
rect 13553 22593 13587 22627
rect 16865 22593 16899 22627
rect 18278 22593 18312 22627
rect 18705 22593 18739 22627
rect 18797 22593 18831 22627
rect 20269 22593 20303 22627
rect 23857 22593 23891 22627
rect 24961 22593 24995 22627
rect 27485 22593 27519 22627
rect 27721 22593 27755 22627
rect 27905 22593 27939 22627
rect 30113 22593 30147 22627
rect 30205 22593 30239 22627
rect 30849 22593 30883 22627
rect 31217 22593 31251 22627
rect 33609 22593 33643 22627
rect 33793 22593 33827 22627
rect 33977 22593 34011 22627
rect 35081 22593 35115 22627
rect 35357 22593 35391 22627
rect 35449 22593 35483 22627
rect 36093 22593 36127 22627
rect 36277 22593 36311 22627
rect 37841 22593 37875 22627
rect 38945 22593 38979 22627
rect 39038 22593 39072 22627
rect 39221 22593 39255 22627
rect 39451 22593 39485 22627
rect 13645 22525 13679 22559
rect 20545 22525 20579 22559
rect 24041 22525 24075 22559
rect 24869 22525 24903 22559
rect 25329 22525 25363 22559
rect 29745 22525 29779 22559
rect 29929 22525 29963 22559
rect 30665 22525 30699 22559
rect 37473 22525 37507 22559
rect 37933 22525 37967 22559
rect 27353 22457 27387 22491
rect 31125 22457 31159 22491
rect 34161 22457 34195 22491
rect 17141 22389 17175 22423
rect 18153 22389 18187 22423
rect 19901 22389 19935 22423
rect 28549 22389 28583 22423
rect 28733 22389 28767 22423
rect 39589 22389 39623 22423
rect 13553 22185 13587 22219
rect 20637 22185 20671 22219
rect 39497 22185 39531 22219
rect 43177 22185 43211 22219
rect 20729 22117 20763 22151
rect 21925 22117 21959 22151
rect 30205 22117 30239 22151
rect 34897 22117 34931 22151
rect 13369 22049 13403 22083
rect 18797 22049 18831 22083
rect 21097 22049 21131 22083
rect 30021 22049 30055 22083
rect 32689 22049 32723 22083
rect 40509 22049 40543 22083
rect 10793 21981 10827 22015
rect 13277 21981 13311 22015
rect 14657 21981 14691 22015
rect 15301 21981 15335 22015
rect 19809 21981 19843 22015
rect 19901 21981 19935 22015
rect 19993 21981 20027 22015
rect 20177 21981 20211 22015
rect 22109 21981 22143 22015
rect 22201 21981 22235 22015
rect 22385 21981 22419 22015
rect 22477 21981 22511 22015
rect 24869 21981 24903 22015
rect 25237 21981 25271 22015
rect 27169 21981 27203 22015
rect 27261 21981 27295 22015
rect 27537 21981 27571 22015
rect 27997 21981 28031 22015
rect 28181 21981 28215 22015
rect 29837 21981 29871 22015
rect 30297 21981 30331 22015
rect 35173 21981 35207 22015
rect 39221 21981 39255 22015
rect 39313 21981 39347 22015
rect 41797 21981 41831 22015
rect 42064 21981 42098 22015
rect 11060 21913 11094 21947
rect 14381 21913 14415 21947
rect 15485 21913 15519 21947
rect 18521 21913 18555 21947
rect 24961 21913 24995 21947
rect 25053 21913 25087 21947
rect 27353 21913 27387 21947
rect 32422 21913 32456 21947
rect 33333 21913 33367 21947
rect 33517 21913 33551 21947
rect 34897 21913 34931 21947
rect 39497 21913 39531 21947
rect 40141 21913 40175 21947
rect 40325 21913 40359 21947
rect 12173 21845 12207 21879
rect 14479 21845 14513 21879
rect 14565 21845 14599 21879
rect 15117 21845 15151 21879
rect 18153 21845 18187 21879
rect 18613 21845 18647 21879
rect 19533 21845 19567 21879
rect 24685 21845 24719 21879
rect 26985 21845 27019 21879
rect 28273 21845 28307 21879
rect 31309 21845 31343 21879
rect 33701 21845 33735 21879
rect 35081 21845 35115 21879
rect 24961 21641 24995 21675
rect 25605 21641 25639 21675
rect 40693 21641 40727 21675
rect 15209 21573 15243 21607
rect 20177 21573 20211 21607
rect 20361 21573 20395 21607
rect 21189 21573 21223 21607
rect 31217 21573 31251 21607
rect 31401 21573 31435 21607
rect 33977 21573 34011 21607
rect 35725 21573 35759 21607
rect 37749 21573 37783 21607
rect 38945 21573 38979 21607
rect 43177 21573 43211 21607
rect 12081 21505 12115 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 15669 21505 15703 21539
rect 15853 21505 15887 21539
rect 21373 21505 21407 21539
rect 21465 21505 21499 21539
rect 22109 21505 22143 21539
rect 22385 21505 22419 21539
rect 22661 21505 22695 21539
rect 22937 21505 22971 21539
rect 23029 21505 23063 21539
rect 25789 21505 25823 21539
rect 25881 21505 25915 21539
rect 27445 21505 27479 21539
rect 27721 21505 27755 21539
rect 28181 21505 28215 21539
rect 28641 21505 28675 21539
rect 32689 21505 32723 21539
rect 33793 21505 33827 21539
rect 34069 21505 34103 21539
rect 34161 21505 34195 21539
rect 35449 21505 35483 21539
rect 37473 21505 37507 21539
rect 37657 21505 37691 21539
rect 37841 21505 37875 21539
rect 38669 21505 38703 21539
rect 38762 21505 38796 21539
rect 39037 21505 39071 21539
rect 39175 21505 39209 21539
rect 41806 21505 41840 21539
rect 42073 21505 42107 21539
rect 42901 21505 42935 21539
rect 12173 21437 12207 21471
rect 12449 21437 12483 21471
rect 15209 21437 15243 21471
rect 16865 21437 16899 21471
rect 17141 21437 17175 21471
rect 21189 21437 21223 21471
rect 24483 21437 24517 21471
rect 24961 21437 24995 21471
rect 25053 21437 25087 21471
rect 25605 21437 25639 21471
rect 31125 21437 31159 21471
rect 32321 21437 32355 21471
rect 32781 21437 32815 21471
rect 35357 21437 35391 21471
rect 35817 21437 35851 21471
rect 27261 21369 27295 21403
rect 34345 21369 34379 21403
rect 38025 21369 38059 21403
rect 15761 21301 15795 21335
rect 18429 21301 18463 21335
rect 20085 21301 20119 21335
rect 23397 21301 23431 21335
rect 31677 21301 31711 21335
rect 35173 21301 35207 21335
rect 39313 21301 39347 21335
rect 13369 21097 13403 21131
rect 16957 21097 16991 21131
rect 24961 21097 24995 21131
rect 25145 21097 25179 21131
rect 25697 21097 25731 21131
rect 29745 21097 29779 21131
rect 30113 21097 30147 21131
rect 40601 21097 40635 21131
rect 19533 21029 19567 21063
rect 21005 21029 21039 21063
rect 27537 21029 27571 21063
rect 38393 21029 38427 21063
rect 16037 20961 16071 20995
rect 17141 20961 17175 20995
rect 19441 20961 19475 20995
rect 21557 20961 21591 20995
rect 31217 20961 31251 20995
rect 31401 20961 31435 20995
rect 32413 20961 32447 20995
rect 32597 20961 32631 20995
rect 37105 20961 37139 20995
rect 37841 20961 37875 20995
rect 38853 20961 38887 20995
rect 39405 20961 39439 20995
rect 40141 20961 40175 20995
rect 43177 20961 43211 20995
rect 11989 20893 12023 20927
rect 12265 20893 12299 20927
rect 14933 20893 14967 20927
rect 15025 20893 15059 20927
rect 15209 20893 15243 20927
rect 15301 20893 15335 20927
rect 16221 20893 16255 20927
rect 17233 20893 17267 20927
rect 21281 20893 21315 20927
rect 22845 20893 22879 20927
rect 23029 20893 23063 20927
rect 24593 20893 24627 20927
rect 24961 20893 24995 20927
rect 25605 20893 25639 20927
rect 25789 20893 25823 20927
rect 29745 20893 29779 20927
rect 29929 20893 29963 20927
rect 31585 20893 31619 20927
rect 31677 20893 31711 20927
rect 32689 20893 32723 20927
rect 33793 20893 33827 20927
rect 34161 20893 34195 20927
rect 35081 20893 35115 20927
rect 35449 20893 35483 20927
rect 37013 20893 37047 20927
rect 38117 20893 38151 20927
rect 38209 20893 38243 20927
rect 39037 20893 39071 20927
rect 40233 20893 40267 20927
rect 19901 20825 19935 20859
rect 27813 20825 27847 20859
rect 28089 20825 28123 20859
rect 32229 20825 32263 20859
rect 33977 20825 34011 20859
rect 34069 20825 34103 20859
rect 35173 20825 35207 20859
rect 35265 20825 35299 20859
rect 36645 20825 36679 20859
rect 36737 20825 36771 20859
rect 37749 20825 37783 20859
rect 42993 20825 43027 20859
rect 14749 20757 14783 20791
rect 21465 20757 21499 20791
rect 22937 20757 22971 20791
rect 27997 20757 28031 20791
rect 34345 20757 34379 20791
rect 34897 20757 34931 20791
rect 37289 20757 37323 20791
rect 39313 20757 39347 20791
rect 42533 20757 42567 20791
rect 42901 20757 42935 20791
rect 13921 20553 13955 20587
rect 14289 20553 14323 20587
rect 17693 20553 17727 20587
rect 39681 20553 39715 20587
rect 40693 20553 40727 20587
rect 14841 20485 14875 20519
rect 18797 20485 18831 20519
rect 23305 20485 23339 20519
rect 27537 20485 27571 20519
rect 30113 20485 30147 20519
rect 30205 20485 30239 20519
rect 35357 20485 35391 20519
rect 39313 20485 39347 20519
rect 14105 20417 14139 20451
rect 14381 20417 14415 20451
rect 15025 20417 15059 20451
rect 15301 20417 15335 20451
rect 17693 20417 17727 20451
rect 17877 20417 17911 20451
rect 19165 20417 19199 20451
rect 19257 20417 19291 20451
rect 20269 20417 20303 20451
rect 20637 20417 20671 20451
rect 20913 20417 20947 20451
rect 21373 20417 21407 20451
rect 23121 20417 23155 20451
rect 23397 20417 23431 20451
rect 24869 20417 24903 20451
rect 25053 20417 25087 20451
rect 27393 20417 27427 20451
rect 27629 20417 27663 20451
rect 27813 20417 27847 20451
rect 28544 20417 28578 20451
rect 28641 20417 28675 20451
rect 28733 20417 28767 20451
rect 28917 20417 28951 20451
rect 30016 20417 30050 20451
rect 30389 20417 30423 20451
rect 34161 20417 34195 20451
rect 34253 20417 34287 20451
rect 34437 20417 34471 20451
rect 34529 20417 34563 20451
rect 34989 20417 35023 20451
rect 35265 20417 35299 20451
rect 35541 20417 35575 20451
rect 35725 20417 35759 20451
rect 39037 20417 39071 20451
rect 39130 20417 39164 20451
rect 39405 20417 39439 20451
rect 39502 20417 39536 20451
rect 40141 20417 40175 20451
rect 40417 20417 40451 20451
rect 40509 20417 40543 20451
rect 42901 20417 42935 20451
rect 14933 20349 14967 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 43177 20349 43211 20383
rect 15209 20281 15243 20315
rect 18521 20281 18555 20315
rect 22937 20213 22971 20247
rect 25053 20213 25087 20247
rect 27261 20213 27295 20247
rect 28365 20213 28399 20247
rect 29837 20213 29871 20247
rect 33977 20213 34011 20247
rect 40233 20213 40267 20247
rect 14657 20009 14691 20043
rect 15301 20009 15335 20043
rect 18153 20009 18187 20043
rect 23213 20009 23247 20043
rect 29837 20009 29871 20043
rect 30665 20009 30699 20043
rect 43269 20009 43303 20043
rect 25237 19941 25271 19975
rect 15393 19873 15427 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 23765 19873 23799 19907
rect 29745 19873 29779 19907
rect 40141 19873 40175 19907
rect 14933 19805 14967 19839
rect 17969 19805 18003 19839
rect 18153 19805 18187 19839
rect 20177 19805 20211 19839
rect 22937 19805 22971 19839
rect 23029 19805 23063 19839
rect 23305 19805 23339 19839
rect 23949 19805 23983 19839
rect 24041 19805 24075 19839
rect 24961 19805 24995 19839
rect 25697 19805 25731 19839
rect 25881 19805 25915 19839
rect 28069 19805 28103 19839
rect 28181 19805 28215 19839
rect 29009 19805 29043 19839
rect 29193 19805 29227 19839
rect 30021 19805 30055 19839
rect 30205 19805 30239 19839
rect 30665 19805 30699 19839
rect 30849 19805 30883 19839
rect 31769 19805 31803 19839
rect 31861 19805 31895 19839
rect 32045 19805 32079 19839
rect 33880 19805 33914 19839
rect 34069 19805 34103 19839
rect 34252 19805 34286 19839
rect 34345 19805 34379 19839
rect 37105 19805 37139 19839
rect 37198 19805 37232 19839
rect 37381 19805 37415 19839
rect 37473 19805 37507 19839
rect 37570 19805 37604 19839
rect 38853 19805 38887 19839
rect 38946 19805 38980 19839
rect 39129 19805 39163 19839
rect 39221 19805 39255 19839
rect 39318 19805 39352 19839
rect 40049 19805 40083 19839
rect 40325 19805 40359 19839
rect 40417 19805 40451 19839
rect 41889 19805 41923 19839
rect 42156 19805 42190 19839
rect 15117 19737 15151 19771
rect 25053 19737 25087 19771
rect 25237 19737 25271 19771
rect 28457 19737 28491 19771
rect 28549 19737 28583 19771
rect 32505 19737 32539 19771
rect 33977 19737 34011 19771
rect 15025 19669 15059 19703
rect 20177 19669 20211 19703
rect 22753 19669 22787 19703
rect 23765 19669 23799 19703
rect 25789 19669 25823 19703
rect 27905 19669 27939 19703
rect 29009 19669 29043 19703
rect 33701 19669 33735 19703
rect 37749 19669 37783 19703
rect 39497 19669 39531 19703
rect 40601 19669 40635 19703
rect 14841 19465 14875 19499
rect 16313 19465 16347 19499
rect 16957 19465 16991 19499
rect 22937 19465 22971 19499
rect 23949 19465 23983 19499
rect 28733 19465 28767 19499
rect 31769 19465 31803 19499
rect 32321 19465 32355 19499
rect 34161 19465 34195 19499
rect 39773 19465 39807 19499
rect 41613 19465 41647 19499
rect 41705 19465 41739 19499
rect 42993 19465 43027 19499
rect 25605 19397 25639 19431
rect 25973 19397 26007 19431
rect 28273 19397 28307 19431
rect 33456 19397 33490 19431
rect 39405 19397 39439 19431
rect 43085 19397 43119 19431
rect 12173 19329 12207 19363
rect 14657 19329 14691 19363
rect 14933 19329 14967 19363
rect 15945 19329 15979 19363
rect 17325 19329 17359 19363
rect 18245 19329 18279 19363
rect 18337 19329 18371 19363
rect 19441 19329 19475 19363
rect 23121 19329 23155 19363
rect 23305 19329 23339 19363
rect 23857 19329 23891 19363
rect 24041 19329 24075 19363
rect 24777 19329 24811 19363
rect 24869 19329 24903 19363
rect 25145 19329 25179 19363
rect 25789 19329 25823 19363
rect 26065 19329 26099 19363
rect 28089 19329 28123 19363
rect 29193 19329 29227 19363
rect 30389 19329 30423 19363
rect 31401 19329 31435 19363
rect 33701 19329 33735 19363
rect 34529 19329 34563 19363
rect 37473 19329 37507 19363
rect 37749 19329 37783 19363
rect 37841 19329 37875 19363
rect 39589 19329 39623 19363
rect 12449 19261 12483 19295
rect 15853 19261 15887 19295
rect 17233 19261 17267 19295
rect 18521 19261 18555 19295
rect 23397 19261 23431 19295
rect 27905 19261 27939 19295
rect 29101 19261 29135 19295
rect 30297 19261 30331 19295
rect 31309 19261 31343 19295
rect 34621 19261 34655 19295
rect 34805 19261 34839 19295
rect 41797 19261 41831 19295
rect 43177 19261 43211 19295
rect 13737 19193 13771 19227
rect 17877 19193 17911 19227
rect 24593 19193 24627 19227
rect 25053 19193 25087 19227
rect 29377 19193 29411 19227
rect 30757 19193 30791 19227
rect 38025 19193 38059 19227
rect 14473 19125 14507 19159
rect 15669 19125 15703 19159
rect 17233 19125 17267 19159
rect 19533 19125 19567 19159
rect 37565 19125 37599 19159
rect 41245 19125 41279 19159
rect 42625 19125 42659 19159
rect 14289 18921 14323 18955
rect 16497 18921 16531 18955
rect 25237 18921 25271 18955
rect 25605 18921 25639 18955
rect 28457 18921 28491 18955
rect 35357 18921 35391 18955
rect 43177 18921 43211 18955
rect 18613 18785 18647 18819
rect 21465 18785 21499 18819
rect 21649 18785 21683 18819
rect 23305 18785 23339 18819
rect 28641 18785 28675 18819
rect 35357 18785 35391 18819
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 15117 18717 15151 18751
rect 15393 18717 15427 18751
rect 16865 18717 16899 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 19533 18717 19567 18751
rect 19717 18717 19751 18751
rect 20361 18717 20395 18751
rect 20545 18717 20579 18751
rect 25421 18717 25455 18751
rect 25697 18717 25731 18751
rect 28733 18717 28767 18751
rect 28825 18717 28859 18751
rect 28917 18717 28951 18751
rect 34989 18717 35023 18751
rect 36277 18717 36311 18751
rect 36461 18717 36495 18751
rect 41797 18717 41831 18751
rect 42064 18717 42098 18751
rect 15209 18649 15243 18683
rect 16681 18649 16715 18683
rect 17417 18649 17451 18683
rect 18337 18649 18371 18683
rect 19441 18649 19475 18683
rect 23121 18649 23155 18683
rect 15117 18581 15151 18615
rect 17969 18581 18003 18615
rect 18429 18581 18463 18615
rect 20453 18581 20487 18615
rect 21005 18581 21039 18615
rect 21373 18581 21407 18615
rect 22753 18581 22787 18615
rect 23213 18581 23247 18615
rect 35173 18581 35207 18615
rect 36369 18581 36403 18615
rect 15393 18377 15427 18411
rect 18705 18377 18739 18411
rect 19901 18377 19935 18411
rect 22937 18377 22971 18411
rect 28641 18377 28675 18411
rect 38853 18377 38887 18411
rect 42073 18377 42107 18411
rect 17325 18309 17359 18343
rect 22753 18309 22787 18343
rect 23029 18309 23063 18343
rect 28457 18309 28491 18343
rect 30205 18309 30239 18343
rect 34805 18309 34839 18343
rect 40960 18309 40994 18343
rect 43177 18309 43211 18343
rect 15025 18241 15059 18275
rect 15209 18241 15243 18275
rect 17509 18241 17543 18275
rect 18429 18241 18463 18275
rect 18613 18241 18647 18275
rect 19809 18241 19843 18275
rect 20729 18241 20763 18275
rect 20821 18241 20855 18275
rect 28733 18241 28767 18275
rect 33885 18241 33919 18275
rect 35633 18241 35667 18275
rect 36369 18241 36403 18275
rect 37473 18241 37507 18275
rect 37729 18241 37763 18275
rect 39589 18241 39623 18275
rect 40693 18241 40727 18275
rect 42901 18241 42935 18275
rect 20085 18173 20119 18207
rect 29377 18173 29411 18207
rect 36277 18173 36311 18207
rect 39497 18173 39531 18207
rect 17141 18105 17175 18139
rect 28457 18105 28491 18139
rect 34161 18105 34195 18139
rect 34345 18105 34379 18139
rect 19441 18037 19475 18071
rect 22477 18037 22511 18071
rect 36645 18037 36679 18071
rect 39957 18037 39991 18071
rect 14657 17833 14691 17867
rect 22385 17833 22419 17867
rect 37657 17833 37691 17867
rect 41429 17833 41463 17867
rect 15117 17765 15151 17799
rect 28365 17765 28399 17799
rect 33793 17765 33827 17799
rect 16681 17697 16715 17731
rect 18797 17697 18831 17731
rect 22477 17697 22511 17731
rect 29745 17697 29779 17731
rect 32965 17697 32999 17731
rect 36277 17697 36311 17731
rect 14565 17629 14599 17663
rect 14657 17629 14691 17663
rect 15301 17629 15335 17663
rect 15577 17629 15611 17663
rect 16957 17629 16991 17663
rect 18705 17629 18739 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 19993 17629 20027 17663
rect 20085 17629 20119 17663
rect 22201 17629 22235 17663
rect 23029 17629 23063 17663
rect 23213 17629 23247 17663
rect 26525 17629 26559 17663
rect 28641 17629 28675 17663
rect 33425 17629 33459 17663
rect 33793 17629 33827 17663
rect 33977 17629 34011 17663
rect 35817 17629 35851 17663
rect 36544 17629 36578 17663
rect 40049 17629 40083 17663
rect 40305 17629 40339 17663
rect 42901 17629 42935 17663
rect 14381 17561 14415 17595
rect 15485 17561 15519 17595
rect 16773 17561 16807 17595
rect 26792 17561 26826 17595
rect 28365 17561 28399 17595
rect 30012 17561 30046 17595
rect 32698 17561 32732 17595
rect 35081 17561 35115 17595
rect 43177 17561 43211 17595
rect 19533 17493 19567 17527
rect 22017 17493 22051 17527
rect 23029 17493 23063 17527
rect 27905 17493 27939 17527
rect 28549 17493 28583 17527
rect 31125 17493 31159 17527
rect 31585 17493 31619 17527
rect 15301 17289 15335 17323
rect 27169 17289 27203 17323
rect 27537 17289 27571 17323
rect 31309 17289 31343 17323
rect 31769 17289 31803 17323
rect 35725 17289 35759 17323
rect 21097 17221 21131 17255
rect 22017 17221 22051 17255
rect 22201 17221 22235 17255
rect 25605 17221 25639 17255
rect 27629 17221 27663 17255
rect 35265 17221 35299 17255
rect 15025 17153 15059 17187
rect 15117 17153 15151 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 16313 17153 16347 17187
rect 17141 17153 17175 17187
rect 17877 17153 17911 17187
rect 18245 17153 18279 17187
rect 19349 17153 19383 17187
rect 19533 17153 19567 17187
rect 19625 17153 19659 17187
rect 20913 17153 20947 17187
rect 22845 17153 22879 17187
rect 23029 17153 23063 17187
rect 24225 17153 24259 17187
rect 30389 17153 30423 17187
rect 31401 17153 31435 17187
rect 33517 17153 33551 17187
rect 34345 17153 34379 17187
rect 17417 17085 17451 17119
rect 20545 17085 20579 17119
rect 23949 17085 23983 17119
rect 27813 17085 27847 17119
rect 31217 17085 31251 17119
rect 34805 17085 34839 17119
rect 16865 17017 16899 17051
rect 35541 17017 35575 17051
rect 19165 16949 19199 16983
rect 22293 16949 22327 16983
rect 22937 16949 22971 16983
rect 29101 16949 29135 16983
rect 33701 16949 33735 16983
rect 16497 16745 16531 16779
rect 17601 16745 17635 16779
rect 23581 16745 23615 16779
rect 27353 16745 27387 16779
rect 27537 16745 27571 16779
rect 28641 16745 28675 16779
rect 22109 16677 22143 16711
rect 18429 16609 18463 16643
rect 18521 16609 18555 16643
rect 20729 16609 20763 16643
rect 24869 16609 24903 16643
rect 28273 16609 28307 16643
rect 29837 16609 29871 16643
rect 31861 16609 31895 16643
rect 32321 16609 32355 16643
rect 38301 16609 38335 16643
rect 38393 16609 38427 16643
rect 41521 16609 41555 16643
rect 16957 16541 16991 16575
rect 17785 16541 17819 16575
rect 18797 16541 18831 16575
rect 20545 16541 20579 16575
rect 22017 16541 22051 16575
rect 22385 16541 22419 16575
rect 22661 16541 22695 16575
rect 23397 16541 23431 16575
rect 23581 16541 23615 16575
rect 25125 16541 25159 16575
rect 30665 16541 30699 16575
rect 31309 16541 31343 16575
rect 32045 16541 32079 16575
rect 32413 16541 32447 16575
rect 35633 16541 35667 16575
rect 35817 16541 35851 16575
rect 35909 16541 35943 16575
rect 36001 16541 36035 16575
rect 20821 16473 20855 16507
rect 20913 16473 20947 16507
rect 27169 16473 27203 16507
rect 28089 16473 28123 16507
rect 31401 16473 31435 16507
rect 38209 16473 38243 16507
rect 41254 16473 41288 16507
rect 26249 16405 26283 16439
rect 27369 16405 27403 16439
rect 28181 16405 28215 16439
rect 36277 16405 36311 16439
rect 37841 16405 37875 16439
rect 40141 16405 40175 16439
rect 22569 16201 22603 16235
rect 27629 16201 27663 16235
rect 29929 16201 29963 16235
rect 30297 16201 30331 16235
rect 31769 16201 31803 16235
rect 37565 16201 37599 16235
rect 40049 16201 40083 16235
rect 40509 16201 40543 16235
rect 22201 16133 22235 16167
rect 22401 16133 22435 16167
rect 23213 16133 23247 16167
rect 23397 16133 23431 16167
rect 25513 16133 25547 16167
rect 18337 16065 18371 16099
rect 18521 16065 18555 16099
rect 20545 16065 20579 16099
rect 20913 16065 20947 16099
rect 27537 16065 27571 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 31401 16065 31435 16099
rect 31493 16065 31527 16099
rect 33324 16065 33358 16099
rect 34989 16065 35023 16099
rect 35256 16065 35290 16099
rect 37473 16065 37507 16099
rect 38301 16065 38335 16099
rect 38945 16065 38979 16099
rect 40141 16065 40175 16099
rect 23857 15997 23891 16031
rect 24133 15997 24167 16031
rect 27813 15997 27847 16031
rect 30389 15997 30423 16031
rect 30481 15997 30515 16031
rect 33057 15997 33091 16031
rect 38485 15997 38519 16031
rect 38669 15997 38703 16031
rect 39865 15997 39899 16031
rect 19993 15861 20027 15895
rect 21097 15861 21131 15895
rect 22385 15861 22419 15895
rect 23029 15861 23063 15895
rect 27169 15861 27203 15895
rect 34437 15861 34471 15895
rect 36369 15861 36403 15895
rect 43361 15861 43395 15895
rect 27629 15657 27663 15691
rect 34345 15657 34379 15691
rect 35449 15657 35483 15691
rect 38853 15657 38887 15691
rect 20729 15589 20763 15623
rect 18061 15521 18095 15555
rect 22845 15521 22879 15555
rect 23673 15521 23707 15555
rect 30205 15521 30239 15555
rect 30297 15521 30331 15555
rect 36001 15521 36035 15555
rect 18337 15453 18371 15487
rect 18797 15453 18831 15487
rect 20269 15453 20303 15487
rect 20545 15453 20579 15487
rect 20913 15453 20947 15487
rect 21281 15453 21315 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 23581 15453 23615 15487
rect 26249 15453 26283 15487
rect 30113 15453 30147 15487
rect 32597 15453 32631 15487
rect 32965 15453 32999 15487
rect 34161 15453 34195 15487
rect 37473 15453 37507 15487
rect 37740 15453 37774 15487
rect 22109 15385 22143 15419
rect 26516 15385 26550 15419
rect 33977 15385 34011 15419
rect 35817 15385 35851 15419
rect 18797 15317 18831 15351
rect 29745 15317 29779 15351
rect 32045 15317 32079 15351
rect 35909 15317 35943 15351
rect 18245 15113 18279 15147
rect 22109 15113 22143 15147
rect 29929 15113 29963 15147
rect 30757 15113 30791 15147
rect 41153 15113 41187 15147
rect 28816 15045 28850 15079
rect 33701 15045 33735 15079
rect 16865 14977 16899 15011
rect 18981 14977 19015 15011
rect 19165 14977 19199 15011
rect 19993 14977 20027 15011
rect 20361 14977 20395 15011
rect 20637 14977 20671 15011
rect 22293 14977 22327 15011
rect 22385 14977 22419 15011
rect 22661 14977 22695 15011
rect 23857 14977 23891 15011
rect 24041 14977 24075 15011
rect 28549 14977 28583 15011
rect 30389 14977 30423 15011
rect 30573 14977 30607 15011
rect 32413 14977 32447 15011
rect 33793 14977 33827 15011
rect 35633 14977 35667 15011
rect 35817 14977 35851 15011
rect 35909 14977 35943 15011
rect 36001 14977 36035 15011
rect 37473 14977 37507 15011
rect 38025 14977 38059 15011
rect 38301 14977 38335 15011
rect 38669 14977 38703 15011
rect 38945 14977 38979 15011
rect 40029 14977 40063 15011
rect 17141 14909 17175 14943
rect 20453 14909 20487 14943
rect 32321 14909 32355 14943
rect 33885 14909 33919 14943
rect 36277 14909 36311 14943
rect 38485 14909 38519 14943
rect 39773 14909 39807 14943
rect 20361 14841 20395 14875
rect 22569 14841 22603 14875
rect 33333 14841 33367 14875
rect 18981 14773 19015 14807
rect 23949 14773 23983 14807
rect 32597 14773 32631 14807
rect 18429 14569 18463 14603
rect 23581 14569 23615 14603
rect 31585 14569 31619 14603
rect 33701 14569 33735 14603
rect 39497 14569 39531 14603
rect 18613 14501 18647 14535
rect 18889 14433 18923 14467
rect 22017 14433 22051 14467
rect 28549 14433 28583 14467
rect 36093 14433 36127 14467
rect 38853 14433 38887 14467
rect 19717 14365 19751 14399
rect 20545 14365 20579 14399
rect 22293 14365 22327 14399
rect 24593 14365 24627 14399
rect 27077 14365 27111 14399
rect 27353 14365 27387 14399
rect 28825 14365 28859 14399
rect 29745 14365 29779 14399
rect 30021 14365 30055 14399
rect 31217 14365 31251 14399
rect 31421 14365 31455 14399
rect 32321 14365 32355 14399
rect 39129 14365 39163 14399
rect 40049 14365 40083 14399
rect 43361 14365 43395 14399
rect 24860 14297 24894 14331
rect 27261 14297 27295 14331
rect 28733 14297 28767 14331
rect 29929 14297 29963 14331
rect 30481 14297 30515 14331
rect 31309 14297 31343 14331
rect 32588 14297 32622 14331
rect 39037 14297 39071 14331
rect 40316 14297 40350 14331
rect 25973 14229 26007 14263
rect 26893 14229 26927 14263
rect 29193 14229 29227 14263
rect 35541 14229 35575 14263
rect 35909 14229 35943 14263
rect 36001 14229 36035 14263
rect 41429 14229 41463 14263
rect 19717 14025 19751 14059
rect 25145 14025 25179 14059
rect 25513 14025 25547 14059
rect 27537 14025 27571 14059
rect 30113 14025 30147 14059
rect 32781 14025 32815 14059
rect 33241 14025 33275 14059
rect 34529 14025 34563 14059
rect 36553 14025 36587 14059
rect 40049 14025 40083 14059
rect 40417 14025 40451 14059
rect 23673 13957 23707 13991
rect 25605 13957 25639 13991
rect 26617 13957 26651 13991
rect 29000 13957 29034 13991
rect 31217 13957 31251 13991
rect 33149 13957 33183 13991
rect 34345 13957 34379 13991
rect 39957 13957 39991 13991
rect 19901 13889 19935 13923
rect 20085 13889 20119 13923
rect 23489 13889 23523 13923
rect 23765 13889 23799 13923
rect 26341 13889 26375 13923
rect 27629 13889 27663 13923
rect 31677 13889 31711 13923
rect 31769 13889 31803 13923
rect 34161 13889 34195 13923
rect 35173 13889 35207 13923
rect 35440 13889 35474 13923
rect 20177 13821 20211 13855
rect 25697 13821 25731 13855
rect 26617 13821 26651 13855
rect 27721 13821 27755 13855
rect 28733 13821 28767 13855
rect 33333 13821 33367 13855
rect 39865 13821 39899 13855
rect 26433 13753 26467 13787
rect 23489 13685 23523 13719
rect 27169 13685 27203 13719
rect 23397 13481 23431 13515
rect 23581 13481 23615 13515
rect 27537 13481 27571 13515
rect 25329 13345 25363 13379
rect 37473 13345 37507 13379
rect 38393 13345 38427 13379
rect 38761 13345 38795 13379
rect 40601 13345 40635 13379
rect 24593 13277 24627 13311
rect 26157 13277 26191 13311
rect 32597 13277 32631 13311
rect 33057 13277 33091 13311
rect 35633 13277 35667 13311
rect 35817 13277 35851 13311
rect 35909 13277 35943 13311
rect 36001 13277 36035 13311
rect 37381 13277 37415 13311
rect 38301 13277 38335 13311
rect 38853 13277 38887 13311
rect 40417 13277 40451 13311
rect 23213 13209 23247 13243
rect 26424 13209 26458 13243
rect 36277 13209 36311 13243
rect 40509 13209 40543 13243
rect 23413 13141 23447 13175
rect 32229 13141 32263 13175
rect 40049 13141 40083 13175
rect 23397 12937 23431 12971
rect 34713 12937 34747 12971
rect 37565 12937 37599 12971
rect 41153 12937 41187 12971
rect 25421 12869 25455 12903
rect 28273 12869 28307 12903
rect 31309 12869 31343 12903
rect 40040 12869 40074 12903
rect 22017 12801 22051 12835
rect 22284 12801 22318 12835
rect 24685 12801 24719 12835
rect 24777 12801 24811 12835
rect 24961 12801 24995 12835
rect 27721 12801 27755 12835
rect 27813 12801 27847 12835
rect 30665 12801 30699 12835
rect 30849 12801 30883 12835
rect 32505 12801 32539 12835
rect 32772 12801 32806 12835
rect 34345 12801 34379 12835
rect 34529 12801 34563 12835
rect 35265 12801 35299 12835
rect 35449 12801 35483 12835
rect 35541 12801 35575 12835
rect 35633 12801 35667 12835
rect 37473 12801 37507 12835
rect 38301 12801 38335 12835
rect 38669 12801 38703 12835
rect 38945 12801 38979 12835
rect 42901 12801 42935 12835
rect 30573 12733 30607 12767
rect 35909 12733 35943 12767
rect 38485 12733 38519 12767
rect 39773 12733 39807 12767
rect 43177 12733 43211 12767
rect 33885 12597 33919 12631
rect 22661 12393 22695 12427
rect 26617 12393 26651 12427
rect 29193 12393 29227 12427
rect 30849 12393 30883 12427
rect 32965 12393 32999 12427
rect 41429 12393 41463 12427
rect 23305 12257 23339 12291
rect 26065 12257 26099 12291
rect 26525 12257 26559 12291
rect 26709 12257 26743 12291
rect 28641 12257 28675 12291
rect 31401 12257 31435 12291
rect 33425 12257 33459 12291
rect 33517 12257 33551 12291
rect 36093 12257 36127 12291
rect 23029 12189 23063 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 25605 12189 25639 12223
rect 25697 12189 25731 12223
rect 25881 12189 25915 12223
rect 26801 12189 26835 12223
rect 33333 12189 33367 12223
rect 40049 12189 40083 12223
rect 28733 12121 28767 12155
rect 36001 12121 36035 12155
rect 40316 12121 40350 12155
rect 23121 12053 23155 12087
rect 28825 12053 28859 12087
rect 31217 12053 31251 12087
rect 31309 12053 31343 12087
rect 35541 12053 35575 12087
rect 35909 12053 35943 12087
rect 23121 11849 23155 11883
rect 24961 11849 24995 11883
rect 26341 11849 26375 11883
rect 28457 11849 28491 11883
rect 30941 11849 30975 11883
rect 34161 11849 34195 11883
rect 36553 11849 36587 11883
rect 40233 11849 40267 11883
rect 40601 11849 40635 11883
rect 24869 11781 24903 11815
rect 28549 11781 28583 11815
rect 33793 11781 33827 11815
rect 35440 11781 35474 11815
rect 38209 11781 38243 11815
rect 40141 11781 40175 11815
rect 23213 11713 23247 11747
rect 26249 11713 26283 11747
rect 30849 11713 30883 11747
rect 33977 11713 34011 11747
rect 35173 11713 35207 11747
rect 38117 11713 38151 11747
rect 42901 11713 42935 11747
rect 23397 11645 23431 11679
rect 25145 11645 25179 11679
rect 26525 11645 26559 11679
rect 28733 11645 28767 11679
rect 31033 11645 31067 11679
rect 38393 11645 38427 11679
rect 39957 11645 39991 11679
rect 43177 11645 43211 11679
rect 22753 11509 22787 11543
rect 24501 11509 24535 11543
rect 25881 11509 25915 11543
rect 28089 11509 28123 11543
rect 30481 11509 30515 11543
rect 37749 11509 37783 11543
rect 23213 11305 23247 11339
rect 25973 11305 26007 11339
rect 28733 11305 28767 11339
rect 31493 11305 31527 11339
rect 33793 11305 33827 11339
rect 36277 11305 36311 11339
rect 38945 11305 38979 11339
rect 27353 11169 27387 11203
rect 30113 11169 30147 11203
rect 32413 11169 32447 11203
rect 34897 11169 34931 11203
rect 21833 11101 21867 11135
rect 24593 11101 24627 11135
rect 24849 11101 24883 11135
rect 27620 11101 27654 11135
rect 30380 11101 30414 11135
rect 37565 11101 37599 11135
rect 37832 11101 37866 11135
rect 22100 11033 22134 11067
rect 32680 11033 32714 11067
rect 35164 11033 35198 11067
rect 26617 10761 26651 10795
rect 29009 10761 29043 10795
rect 31493 10761 31527 10795
rect 32873 10761 32907 10795
rect 33241 10761 33275 10795
rect 35081 10761 35115 10795
rect 35449 10761 35483 10795
rect 38945 10761 38979 10795
rect 33333 10693 33367 10727
rect 35541 10693 35575 10727
rect 25237 10625 25271 10659
rect 25504 10625 25538 10659
rect 27629 10625 27663 10659
rect 27896 10625 27930 10659
rect 30113 10625 30147 10659
rect 30380 10625 30414 10659
rect 37565 10625 37599 10659
rect 37832 10625 37866 10659
rect 33425 10557 33459 10591
rect 35633 10557 35667 10591
rect 28273 10217 28307 10251
rect 30481 10217 30515 10251
rect 37841 10217 37875 10251
rect 28733 10081 28767 10115
rect 28825 10081 28859 10115
rect 30941 10081 30975 10115
rect 31033 10081 31067 10115
rect 38301 10081 38335 10115
rect 38485 10081 38519 10115
rect 28641 10013 28675 10047
rect 30849 10013 30883 10047
rect 38209 10013 38243 10047
rect 42901 10013 42935 10047
rect 43177 9945 43211 9979
rect 42901 8449 42935 8483
rect 43177 8381 43211 8415
rect 42901 6749 42935 6783
rect 43177 6681 43211 6715
rect 42901 5661 42935 5695
rect 43177 5593 43211 5627
rect 42901 4097 42935 4131
rect 43177 4029 43211 4063
rect 42901 2397 42935 2431
rect 43177 2329 43211 2363
<< metal1 >>
rect 16942 44072 16948 44124
rect 17000 44112 17006 44124
rect 18138 44112 18144 44124
rect 17000 44084 18144 44112
rect 17000 44072 17006 44084
rect 18138 44072 18144 44084
rect 18196 44072 18202 44124
rect 1104 42458 43884 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 43884 42458
rect 1104 42384 43884 42406
rect 23382 42304 23388 42356
rect 23440 42344 23446 42356
rect 23440 42316 31616 42344
rect 23440 42304 23446 42316
rect 2961 42279 3019 42285
rect 2961 42245 2973 42279
rect 3007 42276 3019 42279
rect 6917 42279 6975 42285
rect 6917 42276 6929 42279
rect 3007 42248 6929 42276
rect 3007 42245 3019 42248
rect 2961 42239 3019 42245
rect 6917 42245 6929 42248
rect 6963 42276 6975 42279
rect 7190 42276 7196 42288
rect 6963 42248 7196 42276
rect 6963 42245 6975 42248
rect 6917 42239 6975 42245
rect 7190 42236 7196 42248
rect 7248 42236 7254 42288
rect 13357 42279 13415 42285
rect 13357 42245 13369 42279
rect 13403 42276 13415 42279
rect 14366 42276 14372 42288
rect 13403 42248 14372 42276
rect 13403 42245 13415 42248
rect 13357 42239 13415 42245
rect 14366 42236 14372 42248
rect 14424 42276 14430 42288
rect 28350 42276 28356 42288
rect 14424 42248 28356 42276
rect 14424 42236 14430 42248
rect 28350 42236 28356 42248
rect 28408 42276 28414 42288
rect 28537 42279 28595 42285
rect 28537 42276 28549 42279
rect 28408 42248 28549 42276
rect 28408 42236 28414 42248
rect 28537 42245 28549 42248
rect 28583 42245 28595 42279
rect 28537 42239 28595 42245
rect 2222 42168 2228 42220
rect 2280 42208 2286 42220
rect 2409 42211 2467 42217
rect 2409 42208 2421 42211
rect 2280 42180 2421 42208
rect 2280 42168 2286 42180
rect 2409 42177 2421 42180
rect 2455 42177 2467 42211
rect 2409 42171 2467 42177
rect 5902 42168 5908 42220
rect 5960 42168 5966 42220
rect 9674 42168 9680 42220
rect 9732 42208 9738 42220
rect 9769 42211 9827 42217
rect 9769 42208 9781 42211
rect 9732 42180 9781 42208
rect 9732 42168 9738 42180
rect 9769 42177 9781 42180
rect 9815 42177 9827 42211
rect 9769 42171 9827 42177
rect 12437 42211 12495 42217
rect 12437 42177 12449 42211
rect 12483 42208 12495 42211
rect 13262 42208 13268 42220
rect 12483 42180 13268 42208
rect 12483 42177 12495 42180
rect 12437 42171 12495 42177
rect 13262 42168 13268 42180
rect 13320 42168 13326 42220
rect 13449 42211 13507 42217
rect 13449 42177 13461 42211
rect 13495 42208 13507 42211
rect 13722 42208 13728 42220
rect 13495 42180 13728 42208
rect 13495 42177 13507 42180
rect 13449 42171 13507 42177
rect 13722 42168 13728 42180
rect 13780 42168 13786 42220
rect 14550 42168 14556 42220
rect 14608 42208 14614 42220
rect 14645 42211 14703 42217
rect 14645 42208 14657 42211
rect 14608 42180 14657 42208
rect 14608 42168 14614 42180
rect 14645 42177 14657 42180
rect 14691 42177 14703 42211
rect 14645 42171 14703 42177
rect 14737 42211 14795 42217
rect 14737 42177 14749 42211
rect 14783 42208 14795 42211
rect 15102 42208 15108 42220
rect 14783 42180 15108 42208
rect 14783 42177 14795 42180
rect 14737 42171 14795 42177
rect 15102 42168 15108 42180
rect 15160 42168 15166 42220
rect 17218 42168 17224 42220
rect 17276 42208 17282 42220
rect 17276 42180 18092 42208
rect 17276 42168 17282 42180
rect 5626 42100 5632 42152
rect 5684 42100 5690 42152
rect 7006 42100 7012 42152
rect 7064 42100 7070 42152
rect 7193 42143 7251 42149
rect 7193 42109 7205 42143
rect 7239 42140 7251 42143
rect 9214 42140 9220 42152
rect 7239 42112 9220 42140
rect 7239 42109 7251 42112
rect 7193 42103 7251 42109
rect 9214 42100 9220 42112
rect 9272 42100 9278 42152
rect 10318 42100 10324 42152
rect 10376 42100 10382 42152
rect 12161 42143 12219 42149
rect 12161 42109 12173 42143
rect 12207 42109 12219 42143
rect 12161 42103 12219 42109
rect 12176 42072 12204 42103
rect 13630 42100 13636 42152
rect 13688 42140 13694 42152
rect 14921 42143 14979 42149
rect 14921 42140 14933 42143
rect 13688 42112 14933 42140
rect 13688 42100 13694 42112
rect 14921 42109 14933 42112
rect 14967 42109 14979 42143
rect 14921 42103 14979 42109
rect 14550 42072 14556 42084
rect 12176 42044 14556 42072
rect 14550 42032 14556 42044
rect 14608 42032 14614 42084
rect 14936 42072 14964 42103
rect 17310 42100 17316 42152
rect 17368 42100 17374 42152
rect 17497 42143 17555 42149
rect 17497 42109 17509 42143
rect 17543 42140 17555 42143
rect 17770 42140 17776 42152
rect 17543 42112 17776 42140
rect 17543 42109 17555 42112
rect 17497 42103 17555 42109
rect 17512 42072 17540 42103
rect 17770 42100 17776 42112
rect 17828 42100 17834 42152
rect 14936 42044 17540 42072
rect 18064 42072 18092 42180
rect 18138 42168 18144 42220
rect 18196 42168 18202 42220
rect 20714 42168 20720 42220
rect 20772 42208 20778 42220
rect 20809 42211 20867 42217
rect 20809 42208 20821 42211
rect 20772 42180 20821 42208
rect 20772 42168 20778 42180
rect 20809 42177 20821 42180
rect 20855 42177 20867 42211
rect 20809 42171 20867 42177
rect 24302 42168 24308 42220
rect 24360 42208 24366 42220
rect 24581 42211 24639 42217
rect 24581 42208 24593 42211
rect 24360 42180 24593 42208
rect 24360 42168 24366 42180
rect 24581 42177 24593 42180
rect 24627 42177 24639 42211
rect 24581 42171 24639 42177
rect 27246 42168 27252 42220
rect 27304 42168 27310 42220
rect 27982 42168 27988 42220
rect 28040 42208 28046 42220
rect 28169 42211 28227 42217
rect 28169 42208 28181 42211
rect 28040 42180 28181 42208
rect 28040 42168 28046 42180
rect 28169 42177 28181 42180
rect 28215 42177 28227 42211
rect 28169 42171 28227 42177
rect 30558 42168 30564 42220
rect 30616 42168 30622 42220
rect 31588 42217 31616 42316
rect 31754 42236 31760 42288
rect 31812 42276 31818 42288
rect 32401 42279 32459 42285
rect 32401 42276 32413 42279
rect 31812 42248 32413 42276
rect 31812 42236 31818 42248
rect 32401 42245 32413 42248
rect 32447 42245 32459 42279
rect 32401 42239 32459 42245
rect 35342 42236 35348 42288
rect 35400 42276 35406 42288
rect 35529 42279 35587 42285
rect 35529 42276 35541 42279
rect 35400 42248 35541 42276
rect 35400 42236 35406 42248
rect 35529 42245 35541 42248
rect 35575 42245 35587 42279
rect 35529 42239 35587 42245
rect 41877 42279 41935 42285
rect 41877 42245 41889 42279
rect 41923 42276 41935 42279
rect 43990 42276 43996 42288
rect 41923 42248 43996 42276
rect 41923 42245 41935 42248
rect 41877 42239 41935 42245
rect 43990 42236 43996 42248
rect 44048 42236 44054 42288
rect 31573 42211 31631 42217
rect 31573 42177 31585 42211
rect 31619 42208 31631 42211
rect 34146 42208 34152 42220
rect 31619 42180 34152 42208
rect 31619 42177 31631 42180
rect 31573 42171 31631 42177
rect 34146 42168 34152 42180
rect 34204 42208 34210 42220
rect 34204 42180 35894 42208
rect 34204 42168 34210 42180
rect 18690 42100 18696 42152
rect 18748 42100 18754 42152
rect 21361 42143 21419 42149
rect 21361 42109 21373 42143
rect 21407 42109 21419 42143
rect 21361 42103 21419 42109
rect 21376 42072 21404 42103
rect 24946 42100 24952 42152
rect 25004 42100 25010 42152
rect 30377 42143 30435 42149
rect 30377 42109 30389 42143
rect 30423 42109 30435 42143
rect 30377 42103 30435 42109
rect 30006 42072 30012 42084
rect 18064 42044 30012 42072
rect 30006 42032 30012 42044
rect 30064 42032 30070 42084
rect 30392 42072 30420 42103
rect 31570 42072 31576 42084
rect 30392 42044 31576 42072
rect 31570 42032 31576 42044
rect 31628 42032 31634 42084
rect 32582 42032 32588 42084
rect 32640 42032 32646 42084
rect 35866 42072 35894 42180
rect 41598 42168 41604 42220
rect 41656 42168 41662 42220
rect 42702 42168 42708 42220
rect 42760 42168 42766 42220
rect 42981 42143 43039 42149
rect 42981 42109 42993 42143
rect 43027 42109 43039 42143
rect 42981 42103 43039 42109
rect 42996 42072 43024 42103
rect 35866 42044 43024 42072
rect 6546 41964 6552 42016
rect 6604 41964 6610 42016
rect 12986 41964 12992 42016
rect 13044 41964 13050 42016
rect 14274 41964 14280 42016
rect 14332 41964 14338 42016
rect 16574 41964 16580 42016
rect 16632 42004 16638 42016
rect 16853 42007 16911 42013
rect 16853 42004 16865 42007
rect 16632 41976 16865 42004
rect 16632 41964 16638 41976
rect 16853 41973 16865 41976
rect 16899 41973 16911 42007
rect 16853 41967 16911 41973
rect 27522 41964 27528 42016
rect 27580 41964 27586 42016
rect 31662 41964 31668 42016
rect 31720 41964 31726 42016
rect 35618 41964 35624 42016
rect 35676 41964 35682 42016
rect 1104 41914 43884 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 43884 41914
rect 1104 41840 43884 41862
rect 6917 41803 6975 41809
rect 6917 41769 6929 41803
rect 6963 41800 6975 41803
rect 7006 41800 7012 41812
rect 6963 41772 7012 41800
rect 6963 41769 6975 41772
rect 6917 41763 6975 41769
rect 7006 41760 7012 41772
rect 7064 41760 7070 41812
rect 26329 41803 26387 41809
rect 26329 41769 26341 41803
rect 26375 41800 26387 41803
rect 27246 41800 27252 41812
rect 26375 41772 27252 41800
rect 26375 41769 26387 41772
rect 26329 41763 26387 41769
rect 27246 41760 27252 41772
rect 27304 41760 27310 41812
rect 24581 41667 24639 41673
rect 24581 41664 24593 41667
rect 21284 41636 24593 41664
rect 5534 41556 5540 41608
rect 5592 41556 5598 41608
rect 5804 41599 5862 41605
rect 5804 41565 5816 41599
rect 5850 41596 5862 41599
rect 6546 41596 6552 41608
rect 5850 41568 6552 41596
rect 5850 41565 5862 41568
rect 5804 41559 5862 41565
rect 6546 41556 6552 41568
rect 6604 41556 6610 41608
rect 9122 41556 9128 41608
rect 9180 41556 9186 41608
rect 12066 41556 12072 41608
rect 12124 41596 12130 41608
rect 12345 41599 12403 41605
rect 12345 41596 12357 41599
rect 12124 41568 12357 41596
rect 12124 41556 12130 41568
rect 12345 41565 12357 41568
rect 12391 41565 12403 41599
rect 12345 41559 12403 41565
rect 12612 41599 12670 41605
rect 12612 41565 12624 41599
rect 12658 41596 12670 41599
rect 12986 41596 12992 41608
rect 12658 41568 12992 41596
rect 12658 41565 12670 41568
rect 12612 41559 12670 41565
rect 12986 41556 12992 41568
rect 13044 41556 13050 41608
rect 16413 41599 16471 41605
rect 16413 41565 16425 41599
rect 16459 41596 16471 41599
rect 16574 41596 16580 41608
rect 16459 41568 16580 41596
rect 16459 41565 16471 41568
rect 16413 41559 16471 41565
rect 16574 41556 16580 41568
rect 16632 41556 16638 41608
rect 16669 41599 16727 41605
rect 16669 41565 16681 41599
rect 16715 41596 16727 41599
rect 17126 41596 17132 41608
rect 16715 41568 17132 41596
rect 16715 41565 16727 41568
rect 16669 41559 16727 41565
rect 17126 41556 17132 41568
rect 17184 41556 17190 41608
rect 19613 41599 19671 41605
rect 19613 41565 19625 41599
rect 19659 41596 19671 41599
rect 20254 41596 20260 41608
rect 19659 41568 20260 41596
rect 19659 41565 19671 41568
rect 19613 41559 19671 41565
rect 20254 41556 20260 41568
rect 20312 41556 20318 41608
rect 21082 41556 21088 41608
rect 21140 41596 21146 41608
rect 21284 41605 21312 41636
rect 24581 41633 24593 41636
rect 24627 41633 24639 41667
rect 24581 41627 24639 41633
rect 27338 41624 27344 41676
rect 27396 41664 27402 41676
rect 27522 41664 27528 41676
rect 27396 41636 27528 41664
rect 27396 41624 27402 41636
rect 27522 41624 27528 41636
rect 27580 41664 27586 41676
rect 27617 41667 27675 41673
rect 27617 41664 27629 41667
rect 27580 41636 27629 41664
rect 27580 41624 27586 41636
rect 27617 41633 27629 41636
rect 27663 41633 27675 41667
rect 27617 41627 27675 41633
rect 30466 41624 30472 41676
rect 30524 41664 30530 41676
rect 32125 41667 32183 41673
rect 32125 41664 32137 41667
rect 30524 41636 32137 41664
rect 30524 41624 30530 41636
rect 32125 41633 32137 41636
rect 32171 41633 32183 41667
rect 32125 41627 32183 41633
rect 32401 41667 32459 41673
rect 32401 41633 32413 41667
rect 32447 41664 32459 41667
rect 34606 41664 34612 41676
rect 32447 41636 34612 41664
rect 32447 41633 32459 41636
rect 32401 41627 32459 41633
rect 34606 41624 34612 41636
rect 34664 41664 34670 41676
rect 34885 41667 34943 41673
rect 34885 41664 34897 41667
rect 34664 41636 34897 41664
rect 34664 41624 34670 41636
rect 34885 41633 34897 41636
rect 34931 41633 34943 41667
rect 34885 41627 34943 41633
rect 21269 41599 21327 41605
rect 21269 41596 21281 41599
rect 21140 41568 21281 41596
rect 21140 41556 21146 41568
rect 21269 41565 21281 41568
rect 21315 41565 21327 41599
rect 21269 41559 21327 41565
rect 22830 41556 22836 41608
rect 22888 41596 22894 41608
rect 23382 41596 23388 41608
rect 22888 41568 23388 41596
rect 22888 41556 22894 41568
rect 23382 41556 23388 41568
rect 23440 41596 23446 41608
rect 23845 41599 23903 41605
rect 23845 41596 23857 41599
rect 23440 41568 23857 41596
rect 23440 41556 23446 41568
rect 23845 41565 23857 41568
rect 23891 41565 23903 41599
rect 23845 41559 23903 41565
rect 9392 41531 9450 41537
rect 9392 41497 9404 41531
rect 9438 41528 9450 41531
rect 9582 41528 9588 41540
rect 9438 41500 9588 41528
rect 9438 41497 9450 41500
rect 9392 41491 9450 41497
rect 9582 41488 9588 41500
rect 9640 41488 9646 41540
rect 17402 41488 17408 41540
rect 17460 41488 17466 41540
rect 19521 41531 19579 41537
rect 19521 41528 19533 41531
rect 18630 41500 19533 41528
rect 19521 41497 19533 41500
rect 19567 41497 19579 41531
rect 19521 41491 19579 41497
rect 21174 41488 21180 41540
rect 21232 41528 21238 41540
rect 21545 41531 21603 41537
rect 21545 41528 21557 41531
rect 21232 41500 21557 41528
rect 21232 41488 21238 41500
rect 21545 41497 21557 41500
rect 21591 41497 21603 41531
rect 21545 41491 21603 41497
rect 22278 41488 22284 41540
rect 22336 41488 22342 41540
rect 24026 41488 24032 41540
rect 24084 41528 24090 41540
rect 24857 41531 24915 41537
rect 24857 41528 24869 41531
rect 24084 41500 24869 41528
rect 24084 41488 24090 41500
rect 24857 41497 24869 41500
rect 24903 41497 24915 41531
rect 24857 41491 24915 41497
rect 24964 41500 25346 41528
rect 10042 41420 10048 41472
rect 10100 41460 10106 41472
rect 10505 41463 10563 41469
rect 10505 41460 10517 41463
rect 10100 41432 10517 41460
rect 10100 41420 10106 41432
rect 10505 41429 10517 41432
rect 10551 41429 10563 41463
rect 10505 41423 10563 41429
rect 13722 41420 13728 41472
rect 13780 41420 13786 41472
rect 15289 41463 15347 41469
rect 15289 41429 15301 41463
rect 15335 41460 15347 41463
rect 17310 41460 17316 41472
rect 15335 41432 17316 41460
rect 15335 41429 15347 41432
rect 15289 41423 15347 41429
rect 17310 41420 17316 41432
rect 17368 41460 17374 41472
rect 17586 41460 17592 41472
rect 17368 41432 17592 41460
rect 17368 41420 17374 41432
rect 17586 41420 17592 41432
rect 17644 41420 17650 41472
rect 18877 41463 18935 41469
rect 18877 41429 18889 41463
rect 18923 41460 18935 41463
rect 22554 41460 22560 41472
rect 18923 41432 22560 41460
rect 18923 41429 18935 41432
rect 18877 41423 18935 41429
rect 22554 41420 22560 41432
rect 22612 41420 22618 41472
rect 23017 41463 23075 41469
rect 23017 41429 23029 41463
rect 23063 41460 23075 41463
rect 23842 41460 23848 41472
rect 23063 41432 23848 41460
rect 23063 41429 23075 41432
rect 23017 41423 23075 41429
rect 23842 41420 23848 41432
rect 23900 41420 23906 41472
rect 23937 41463 23995 41469
rect 23937 41429 23949 41463
rect 23983 41460 23995 41463
rect 24964 41460 24992 41500
rect 26970 41488 26976 41540
rect 27028 41528 27034 41540
rect 27065 41531 27123 41537
rect 27065 41528 27077 41531
rect 27028 41500 27077 41528
rect 27028 41488 27034 41500
rect 27065 41497 27077 41500
rect 27111 41497 27123 41531
rect 27065 41491 27123 41497
rect 23983 41432 24992 41460
rect 27724 41460 27752 41582
rect 28534 41556 28540 41608
rect 28592 41596 28598 41608
rect 28721 41599 28779 41605
rect 28721 41596 28733 41599
rect 28592 41568 28733 41596
rect 28592 41556 28598 41568
rect 28721 41565 28733 41568
rect 28767 41596 28779 41599
rect 28902 41596 28908 41608
rect 28767 41568 28908 41596
rect 28767 41565 28779 41568
rect 28721 41559 28779 41565
rect 28902 41556 28908 41568
rect 28960 41556 28966 41608
rect 32861 41599 32919 41605
rect 32861 41596 32873 41599
rect 32416 41568 32873 41596
rect 28997 41531 29055 41537
rect 28997 41497 29009 41531
rect 29043 41528 29055 41531
rect 29914 41528 29920 41540
rect 29043 41500 29920 41528
rect 29043 41497 29055 41500
rect 28997 41491 29055 41497
rect 29914 41488 29920 41500
rect 29972 41488 29978 41540
rect 31662 41488 31668 41540
rect 31720 41488 31726 41540
rect 27890 41460 27896 41472
rect 27724 41432 27896 41460
rect 23983 41429 23995 41432
rect 23937 41423 23995 41429
rect 27890 41420 27896 41432
rect 27948 41460 27954 41472
rect 30653 41463 30711 41469
rect 30653 41460 30665 41463
rect 27948 41432 30665 41460
rect 27948 41420 27954 41432
rect 30653 41429 30665 41432
rect 30699 41460 30711 41463
rect 30834 41460 30840 41472
rect 30699 41432 30840 41460
rect 30699 41429 30711 41432
rect 30653 41423 30711 41429
rect 30834 41420 30840 41432
rect 30892 41420 30898 41472
rect 31110 41420 31116 41472
rect 31168 41460 31174 41472
rect 32416 41460 32444 41568
rect 32861 41565 32873 41568
rect 32907 41565 32919 41599
rect 32861 41559 32919 41565
rect 33962 41556 33968 41608
rect 34020 41605 34026 41608
rect 34020 41599 34053 41605
rect 34041 41565 34053 41599
rect 34020 41559 34053 41565
rect 34149 41599 34207 41605
rect 34149 41565 34161 41599
rect 34195 41596 34207 41599
rect 34238 41596 34244 41608
rect 34195 41568 34244 41596
rect 34195 41565 34207 41568
rect 34149 41559 34207 41565
rect 34020 41556 34026 41559
rect 34238 41556 34244 41568
rect 34296 41556 34302 41608
rect 34900 41596 34928 41627
rect 41598 41624 41604 41676
rect 41656 41664 41662 41676
rect 41656 41636 42288 41664
rect 41656 41624 41662 41636
rect 35526 41596 35532 41608
rect 34900 41568 35532 41596
rect 35526 41556 35532 41568
rect 35584 41596 35590 41608
rect 37921 41599 37979 41605
rect 37921 41596 37933 41599
rect 35584 41568 37933 41596
rect 35584 41556 35590 41568
rect 37921 41565 37933 41568
rect 37967 41596 37979 41599
rect 40037 41599 40095 41605
rect 40037 41596 40049 41599
rect 37967 41568 40049 41596
rect 37967 41565 37979 41568
rect 37921 41559 37979 41565
rect 40037 41565 40049 41568
rect 40083 41596 40095 41599
rect 41874 41596 41880 41608
rect 40083 41568 41880 41596
rect 40083 41565 40095 41568
rect 40037 41559 40095 41565
rect 41874 41556 41880 41568
rect 41932 41556 41938 41608
rect 42260 41605 42288 41636
rect 42245 41599 42303 41605
rect 42245 41565 42257 41599
rect 42291 41565 42303 41599
rect 42245 41559 42303 41565
rect 42337 41599 42395 41605
rect 42337 41565 42349 41599
rect 42383 41596 42395 41599
rect 42889 41599 42947 41605
rect 42889 41596 42901 41599
rect 42383 41568 42901 41596
rect 42383 41565 42395 41568
rect 42337 41559 42395 41565
rect 42889 41565 42901 41568
rect 42935 41565 42947 41599
rect 42889 41559 42947 41565
rect 32490 41488 32496 41540
rect 32548 41528 32554 41540
rect 33137 41531 33195 41537
rect 33137 41528 33149 41531
rect 32548 41500 33149 41528
rect 32548 41488 32554 41500
rect 33137 41497 33149 41500
rect 33183 41497 33195 41531
rect 33137 41491 33195 41497
rect 35152 41531 35210 41537
rect 35152 41497 35164 41531
rect 35198 41528 35210 41531
rect 35342 41528 35348 41540
rect 35198 41500 35348 41528
rect 35198 41497 35210 41500
rect 35152 41491 35210 41497
rect 35342 41488 35348 41500
rect 35400 41488 35406 41540
rect 38010 41488 38016 41540
rect 38068 41528 38074 41540
rect 38166 41531 38224 41537
rect 38166 41528 38178 41531
rect 38068 41500 38178 41528
rect 38068 41488 38074 41500
rect 38166 41497 38178 41500
rect 38212 41497 38224 41531
rect 38166 41491 38224 41497
rect 40126 41488 40132 41540
rect 40184 41528 40190 41540
rect 40282 41531 40340 41537
rect 40282 41528 40294 41531
rect 40184 41500 40294 41528
rect 40184 41488 40190 41500
rect 40282 41497 40294 41500
rect 40328 41497 40340 41531
rect 40282 41491 40340 41497
rect 43165 41531 43223 41537
rect 43165 41497 43177 41531
rect 43211 41528 43223 41531
rect 43990 41528 43996 41540
rect 43211 41500 43996 41528
rect 43211 41497 43223 41500
rect 43165 41491 43223 41497
rect 43990 41488 43996 41500
rect 44048 41488 44054 41540
rect 31168 41432 32444 41460
rect 33781 41463 33839 41469
rect 31168 41420 31174 41432
rect 33781 41429 33793 41463
rect 33827 41460 33839 41463
rect 33870 41460 33876 41472
rect 33827 41432 33876 41460
rect 33827 41429 33839 41432
rect 33781 41423 33839 41429
rect 33870 41420 33876 41432
rect 33928 41420 33934 41472
rect 35894 41420 35900 41472
rect 35952 41460 35958 41472
rect 36265 41463 36323 41469
rect 36265 41460 36277 41463
rect 35952 41432 36277 41460
rect 35952 41420 35958 41432
rect 36265 41429 36277 41432
rect 36311 41429 36323 41463
rect 36265 41423 36323 41429
rect 39298 41420 39304 41472
rect 39356 41420 39362 41472
rect 41414 41420 41420 41472
rect 41472 41420 41478 41472
rect 1104 41370 43884 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 43884 41370
rect 1104 41296 43884 41318
rect 6822 41216 6828 41268
rect 6880 41256 6886 41268
rect 6880 41228 9260 41256
rect 6880 41216 6886 41228
rect 5534 41148 5540 41200
rect 5592 41188 5598 41200
rect 9122 41188 9128 41200
rect 5592 41160 9128 41188
rect 5592 41148 5598 41160
rect 7668 41129 7696 41160
rect 9122 41148 9128 41160
rect 9180 41148 9186 41200
rect 9232 41188 9260 41228
rect 9582 41216 9588 41268
rect 9640 41216 9646 41268
rect 12158 41216 12164 41268
rect 12216 41216 12222 41268
rect 17405 41259 17463 41265
rect 12406 41228 17356 41256
rect 12406 41188 12434 41228
rect 9232 41160 12434 41188
rect 14176 41191 14234 41197
rect 14176 41157 14188 41191
rect 14222 41188 14234 41191
rect 14274 41188 14280 41200
rect 14222 41160 14280 41188
rect 14222 41157 14234 41160
rect 14176 41151 14234 41157
rect 14274 41148 14280 41160
rect 14332 41148 14338 41200
rect 14550 41148 14556 41200
rect 14608 41188 14614 41200
rect 14608 41160 15976 41188
rect 14608 41148 14614 41160
rect 7653 41123 7711 41129
rect 7653 41089 7665 41123
rect 7699 41089 7711 41123
rect 7653 41083 7711 41089
rect 7920 41123 7978 41129
rect 7920 41089 7932 41123
rect 7966 41120 7978 41123
rect 8386 41120 8392 41132
rect 7966 41092 8392 41120
rect 7966 41089 7978 41092
rect 7920 41083 7978 41089
rect 8386 41080 8392 41092
rect 8444 41080 8450 41132
rect 9953 41123 10011 41129
rect 9953 41089 9965 41123
rect 9999 41120 10011 41123
rect 10318 41120 10324 41132
rect 9999 41092 10324 41120
rect 9999 41089 10011 41092
rect 9953 41083 10011 41089
rect 10318 41080 10324 41092
rect 10376 41080 10382 41132
rect 11974 41080 11980 41132
rect 12032 41120 12038 41132
rect 12069 41123 12127 41129
rect 12069 41120 12081 41123
rect 12032 41092 12081 41120
rect 12032 41080 12038 41092
rect 12069 41089 12081 41092
rect 12115 41120 12127 41123
rect 12115 41092 15792 41120
rect 12115 41089 12127 41092
rect 12069 41083 12127 41089
rect 10042 41012 10048 41064
rect 10100 41012 10106 41064
rect 10137 41055 10195 41061
rect 10137 41021 10149 41055
rect 10183 41052 10195 41055
rect 12253 41055 12311 41061
rect 12253 41052 12265 41055
rect 10183 41024 12265 41052
rect 10183 41021 10195 41024
rect 10137 41015 10195 41021
rect 12253 41021 12265 41024
rect 12299 41052 12311 41055
rect 13630 41052 13636 41064
rect 12299 41024 13636 41052
rect 12299 41021 12311 41024
rect 12253 41015 12311 41021
rect 9214 40944 9220 40996
rect 9272 40984 9278 40996
rect 10152 40984 10180 41015
rect 13630 41012 13636 41024
rect 13688 41012 13694 41064
rect 13909 41055 13967 41061
rect 13909 41021 13921 41055
rect 13955 41021 13967 41055
rect 13909 41015 13967 41021
rect 9272 40956 10180 40984
rect 9272 40944 9278 40956
rect 12066 40944 12072 40996
rect 12124 40984 12130 40996
rect 13924 40984 13952 41015
rect 12124 40956 13952 40984
rect 12124 40944 12130 40956
rect 15010 40944 15016 40996
rect 15068 40984 15074 40996
rect 15764 40984 15792 41092
rect 15838 41080 15844 41132
rect 15896 41080 15902 41132
rect 15948 41120 15976 41160
rect 17218 41148 17224 41200
rect 17276 41148 17282 41200
rect 17328 41188 17356 41228
rect 17405 41225 17417 41259
rect 17451 41256 17463 41259
rect 17586 41256 17592 41268
rect 17451 41228 17592 41256
rect 17451 41225 17463 41228
rect 17405 41219 17463 41225
rect 17586 41216 17592 41228
rect 17644 41216 17650 41268
rect 17696 41228 22094 41256
rect 17696 41188 17724 41228
rect 17328 41160 17724 41188
rect 19705 41191 19763 41197
rect 19705 41157 19717 41191
rect 19751 41188 19763 41191
rect 19978 41188 19984 41200
rect 19751 41160 19984 41188
rect 19751 41157 19763 41160
rect 19705 41151 19763 41157
rect 19978 41148 19984 41160
rect 20036 41148 20042 41200
rect 20346 41148 20352 41200
rect 20404 41148 20410 41200
rect 22066 41188 22094 41228
rect 22278 41216 22284 41268
rect 22336 41256 22342 41268
rect 22373 41259 22431 41265
rect 22373 41256 22385 41259
rect 22336 41228 22385 41256
rect 22336 41216 22342 41228
rect 22373 41225 22385 41228
rect 22419 41225 22431 41259
rect 24394 41256 24400 41268
rect 22373 41219 22431 41225
rect 22480 41228 24400 41256
rect 22480 41188 22508 41228
rect 24394 41216 24400 41228
rect 24452 41216 24458 41268
rect 28626 41256 28632 41268
rect 28276 41228 28632 41256
rect 22066 41160 22508 41188
rect 17497 41123 17555 41129
rect 17497 41120 17509 41123
rect 15948 41092 17509 41120
rect 17497 41089 17509 41092
rect 17543 41120 17555 41123
rect 17954 41120 17960 41132
rect 17543 41092 17960 41120
rect 17543 41089 17555 41092
rect 17497 41083 17555 41089
rect 17954 41080 17960 41092
rect 18012 41080 18018 41132
rect 18046 41080 18052 41132
rect 18104 41080 18110 41132
rect 22278 41080 22284 41132
rect 22336 41120 22342 41132
rect 22830 41120 22836 41132
rect 22336 41092 22836 41120
rect 22336 41080 22342 41092
rect 22830 41080 22836 41092
rect 22888 41080 22894 41132
rect 23201 41123 23259 41129
rect 23201 41089 23213 41123
rect 23247 41089 23259 41123
rect 23201 41083 23259 41089
rect 16117 41055 16175 41061
rect 16117 41021 16129 41055
rect 16163 41052 16175 41055
rect 16482 41052 16488 41064
rect 16163 41024 16488 41052
rect 16163 41021 16175 41024
rect 16117 41015 16175 41021
rect 16482 41012 16488 41024
rect 16540 41012 16546 41064
rect 18325 41055 18383 41061
rect 18325 41021 18337 41055
rect 18371 41052 18383 41055
rect 18414 41052 18420 41064
rect 18371 41024 18420 41052
rect 18371 41021 18383 41024
rect 18325 41015 18383 41021
rect 18414 41012 18420 41024
rect 18472 41012 18478 41064
rect 19429 41055 19487 41061
rect 19429 41021 19441 41055
rect 19475 41021 19487 41055
rect 19429 41015 19487 41021
rect 21177 41055 21235 41061
rect 21177 41021 21189 41055
rect 21223 41052 21235 41055
rect 23216 41052 23244 41083
rect 23842 41080 23848 41132
rect 23900 41120 23906 41132
rect 24118 41120 24124 41132
rect 23900 41092 24124 41120
rect 23900 41080 23906 41092
rect 24118 41080 24124 41092
rect 24176 41080 24182 41132
rect 25222 41080 25228 41132
rect 25280 41080 25286 41132
rect 25501 41123 25559 41129
rect 25501 41089 25513 41123
rect 25547 41120 25559 41123
rect 25958 41120 25964 41132
rect 25547 41092 25964 41120
rect 25547 41089 25559 41092
rect 25501 41083 25559 41089
rect 25958 41080 25964 41092
rect 26016 41120 26022 41132
rect 26421 41123 26479 41129
rect 26421 41120 26433 41123
rect 26016 41092 26433 41120
rect 26016 41080 26022 41092
rect 26421 41089 26433 41092
rect 26467 41089 26479 41123
rect 26421 41083 26479 41089
rect 21223 41024 23244 41052
rect 21223 41021 21235 41024
rect 21177 41015 21235 41021
rect 15068 40956 15424 40984
rect 15764 40956 17080 40984
rect 15068 40944 15074 40956
rect 9030 40876 9036 40928
rect 9088 40876 9094 40928
rect 11698 40876 11704 40928
rect 11756 40876 11762 40928
rect 14642 40876 14648 40928
rect 14700 40916 14706 40928
rect 15102 40916 15108 40928
rect 14700 40888 15108 40916
rect 14700 40876 14706 40888
rect 15102 40876 15108 40888
rect 15160 40916 15166 40928
rect 15289 40919 15347 40925
rect 15289 40916 15301 40919
rect 15160 40888 15301 40916
rect 15160 40876 15166 40888
rect 15289 40885 15301 40888
rect 15335 40885 15347 40919
rect 15396 40916 15424 40956
rect 16945 40919 17003 40925
rect 16945 40916 16957 40919
rect 15396 40888 16957 40916
rect 15289 40879 15347 40885
rect 16945 40885 16957 40888
rect 16991 40885 17003 40919
rect 17052 40916 17080 40956
rect 17126 40944 17132 40996
rect 17184 40984 17190 40996
rect 19444 40984 19472 41015
rect 24670 41012 24676 41064
rect 24728 41052 24734 41064
rect 26234 41052 26240 41064
rect 24728 41024 26240 41052
rect 24728 41012 24734 41024
rect 26234 41012 26240 41024
rect 26292 41012 26298 41064
rect 17184 40956 19472 40984
rect 26436 40984 26464 41083
rect 27246 41080 27252 41132
rect 27304 41080 27310 41132
rect 28276 41118 28304 41228
rect 28626 41216 28632 41228
rect 28684 41216 28690 41268
rect 28810 41216 28816 41268
rect 28868 41256 28874 41268
rect 28994 41256 29000 41268
rect 28868 41228 29000 41256
rect 28868 41216 28874 41228
rect 28994 41216 29000 41228
rect 29052 41216 29058 41268
rect 29086 41216 29092 41268
rect 29144 41256 29150 41268
rect 29144 41228 30512 41256
rect 29144 41216 29150 41228
rect 28644 41160 28856 41188
rect 28644 41129 28672 41160
rect 28353 41123 28411 41129
rect 28353 41118 28365 41123
rect 28276 41090 28365 41118
rect 28353 41089 28365 41090
rect 28399 41089 28411 41123
rect 28353 41083 28411 41089
rect 28537 41123 28595 41129
rect 28537 41089 28549 41123
rect 28583 41089 28595 41123
rect 28537 41083 28595 41089
rect 28629 41123 28687 41129
rect 28629 41089 28641 41123
rect 28675 41089 28687 41123
rect 28629 41083 28687 41089
rect 28721 41123 28779 41129
rect 28721 41089 28733 41123
rect 28767 41089 28779 41123
rect 28828 41120 28856 41160
rect 28902 41148 28908 41200
rect 28960 41188 28966 41200
rect 30484 41188 30512 41228
rect 30834 41216 30840 41268
rect 30892 41256 30898 41268
rect 30892 41228 33640 41256
rect 30892 41216 30898 41228
rect 32309 41191 32367 41197
rect 32309 41188 32321 41191
rect 28960 41160 30420 41188
rect 30484 41160 32321 41188
rect 28960 41148 28966 41160
rect 30098 41120 30104 41132
rect 28828 41092 30104 41120
rect 28721 41083 28779 41089
rect 27801 41055 27859 41061
rect 27801 41021 27813 41055
rect 27847 41052 27859 41055
rect 28074 41052 28080 41064
rect 27847 41024 28080 41052
rect 27847 41021 27859 41024
rect 27801 41015 27859 41021
rect 28074 41012 28080 41024
rect 28132 41012 28138 41064
rect 28442 41012 28448 41064
rect 28500 41052 28506 41064
rect 28552 41052 28580 41083
rect 28736 41052 28764 41083
rect 30098 41080 30104 41092
rect 30156 41080 30162 41132
rect 30190 41080 30196 41132
rect 30248 41120 30254 41132
rect 30392 41129 30420 41160
rect 32309 41157 32321 41160
rect 32355 41157 32367 41191
rect 32309 41151 32367 41157
rect 30285 41123 30343 41129
rect 30285 41120 30297 41123
rect 30248 41092 30297 41120
rect 30248 41080 30254 41092
rect 30285 41089 30297 41092
rect 30331 41089 30343 41123
rect 30285 41083 30343 41089
rect 30377 41123 30435 41129
rect 30377 41089 30389 41123
rect 30423 41120 30435 41123
rect 31018 41120 31024 41132
rect 30423 41092 31024 41120
rect 30423 41089 30435 41092
rect 30377 41083 30435 41089
rect 31018 41080 31024 41092
rect 31076 41080 31082 41132
rect 31110 41080 31116 41132
rect 31168 41126 31174 41132
rect 31168 41120 31248 41126
rect 31168 41098 31340 41120
rect 31168 41080 31174 41098
rect 31220 41092 31340 41098
rect 28500 41024 28580 41052
rect 28644 41024 28764 41052
rect 28500 41012 28506 41024
rect 28534 40984 28540 40996
rect 26436 40956 28540 40984
rect 17184 40944 17190 40956
rect 18690 40916 18696 40928
rect 17052 40888 18696 40916
rect 16945 40879 17003 40885
rect 18690 40876 18696 40888
rect 18748 40876 18754 40928
rect 19444 40916 19472 40956
rect 28534 40944 28540 40956
rect 28592 40944 28598 40996
rect 21082 40916 21088 40928
rect 19444 40888 21088 40916
rect 21082 40876 21088 40888
rect 21140 40876 21146 40928
rect 23474 40876 23480 40928
rect 23532 40876 23538 40928
rect 23842 40876 23848 40928
rect 23900 40916 23906 40928
rect 24946 40916 24952 40928
rect 23900 40888 24952 40916
rect 23900 40876 23906 40888
rect 24946 40876 24952 40888
rect 25004 40876 25010 40928
rect 26605 40919 26663 40925
rect 26605 40885 26617 40919
rect 26651 40916 26663 40919
rect 27062 40916 27068 40928
rect 26651 40888 27068 40916
rect 26651 40885 26663 40888
rect 26605 40879 26663 40885
rect 27062 40876 27068 40888
rect 27120 40876 27126 40928
rect 28442 40876 28448 40928
rect 28500 40916 28506 40928
rect 28644 40916 28672 41024
rect 28810 41012 28816 41064
rect 28868 41052 28874 41064
rect 29457 41055 29515 41061
rect 29457 41052 29469 41055
rect 28868 41024 29469 41052
rect 28868 41012 28874 41024
rect 29457 41021 29469 41024
rect 29503 41021 29515 41055
rect 29457 41015 29515 41021
rect 29825 41055 29883 41061
rect 29825 41021 29837 41055
rect 29871 41021 29883 41055
rect 31312 41052 31340 41092
rect 31662 41080 31668 41132
rect 31720 41080 31726 41132
rect 32490 41129 32496 41132
rect 32456 41123 32496 41129
rect 32456 41089 32468 41123
rect 32456 41083 32496 41089
rect 32490 41080 32496 41083
rect 32548 41080 32554 41132
rect 32030 41052 32036 41064
rect 31312 41024 32036 41052
rect 29825 41015 29883 41021
rect 28718 40944 28724 40996
rect 28776 40984 28782 40996
rect 29840 40984 29868 41015
rect 32030 41012 32036 41024
rect 32088 41052 32094 41064
rect 32677 41055 32735 41061
rect 32677 41052 32689 41055
rect 32088 41024 32689 41052
rect 32088 41012 32094 41024
rect 32677 41021 32689 41024
rect 32723 41021 32735 41055
rect 33612 41052 33640 41228
rect 38010 41216 38016 41268
rect 38068 41216 38074 41268
rect 39945 41259 40003 41265
rect 39945 41225 39957 41259
rect 39991 41256 40003 41259
rect 40126 41256 40132 41268
rect 39991 41228 40132 41256
rect 39991 41225 40003 41228
rect 39945 41219 40003 41225
rect 40126 41216 40132 41228
rect 40184 41216 40190 41268
rect 34238 41188 34244 41200
rect 33704 41160 34244 41188
rect 33704 41132 33732 41160
rect 34238 41148 34244 41160
rect 34296 41148 34302 41200
rect 35618 41148 35624 41200
rect 35676 41188 35682 41200
rect 35774 41191 35832 41197
rect 35774 41188 35786 41191
rect 35676 41160 35786 41188
rect 35676 41148 35682 41160
rect 35774 41157 35786 41160
rect 35820 41157 35832 41191
rect 35774 41151 35832 41157
rect 38378 41148 38384 41200
rect 38436 41188 38442 41200
rect 38749 41191 38807 41197
rect 38749 41188 38761 41191
rect 38436 41160 38761 41188
rect 38436 41148 38442 41160
rect 38749 41157 38761 41160
rect 38795 41157 38807 41191
rect 38749 41151 38807 41157
rect 33686 41080 33692 41132
rect 33744 41080 33750 41132
rect 33873 41123 33931 41129
rect 33873 41089 33885 41123
rect 33919 41120 33931 41123
rect 33962 41120 33968 41132
rect 33919 41092 33968 41120
rect 33919 41089 33931 41092
rect 33873 41083 33931 41089
rect 33888 41052 33916 41083
rect 33962 41080 33968 41092
rect 34020 41080 34026 41132
rect 34256 41120 34284 41148
rect 34547 41123 34605 41129
rect 34547 41120 34559 41123
rect 34256 41092 34559 41120
rect 34547 41089 34559 41092
rect 34593 41089 34605 41123
rect 34547 41083 34605 41089
rect 34701 41123 34759 41129
rect 34701 41089 34713 41123
rect 34747 41089 34759 41123
rect 34701 41083 34759 41089
rect 34716 41052 34744 41083
rect 35526 41080 35532 41132
rect 35584 41080 35590 41132
rect 37645 41123 37703 41129
rect 37645 41089 37657 41123
rect 37691 41120 37703 41123
rect 37691 41092 38516 41120
rect 37691 41089 37703 41092
rect 37645 41083 37703 41089
rect 38488 41064 38516 41092
rect 38562 41080 38568 41132
rect 38620 41120 38626 41132
rect 38933 41123 38991 41129
rect 38933 41120 38945 41123
rect 38620 41092 38945 41120
rect 38620 41080 38626 41092
rect 38933 41089 38945 41092
rect 38979 41089 38991 41123
rect 38933 41083 38991 41089
rect 39117 41123 39175 41129
rect 39117 41089 39129 41123
rect 39163 41120 39175 41123
rect 39761 41123 39819 41129
rect 39761 41120 39773 41123
rect 39163 41092 39773 41120
rect 39163 41089 39175 41092
rect 39117 41083 39175 41089
rect 39761 41089 39773 41092
rect 39807 41089 39819 41123
rect 39761 41083 39819 41089
rect 40678 41080 40684 41132
rect 40736 41120 40742 41132
rect 40845 41123 40903 41129
rect 40845 41120 40857 41123
rect 40736 41092 40857 41120
rect 40736 41080 40742 41092
rect 40845 41089 40857 41092
rect 40891 41089 40903 41123
rect 40845 41083 40903 41089
rect 42889 41123 42947 41129
rect 42889 41089 42901 41123
rect 42935 41120 42947 41123
rect 43070 41120 43076 41132
rect 42935 41092 43076 41120
rect 42935 41089 42947 41092
rect 42889 41083 42947 41089
rect 43070 41080 43076 41092
rect 43128 41080 43134 41132
rect 35434 41052 35440 41064
rect 33612 41024 35440 41052
rect 32677 41015 32735 41021
rect 35434 41012 35440 41024
rect 35492 41012 35498 41064
rect 37550 41012 37556 41064
rect 37608 41012 37614 41064
rect 38470 41012 38476 41064
rect 38528 41052 38534 41064
rect 39577 41055 39635 41061
rect 39577 41052 39589 41055
rect 38528 41024 39589 41052
rect 38528 41012 38534 41024
rect 39577 41021 39589 41024
rect 39623 41021 39635 41055
rect 39577 41015 39635 41021
rect 40034 41012 40040 41064
rect 40092 41052 40098 41064
rect 40589 41055 40647 41061
rect 40589 41052 40601 41055
rect 40092 41024 40601 41052
rect 40092 41012 40098 41024
rect 40589 41021 40601 41024
rect 40635 41021 40647 41055
rect 40589 41015 40647 41021
rect 43165 41055 43223 41061
rect 43165 41021 43177 41055
rect 43211 41052 43223 41055
rect 43990 41052 43996 41064
rect 43211 41024 43996 41052
rect 43211 41021 43223 41024
rect 43165 41015 43223 41021
rect 43990 41012 43996 41024
rect 44048 41012 44054 41064
rect 28776 40956 29868 40984
rect 28776 40944 28782 40956
rect 29914 40944 29920 40996
rect 29972 40944 29978 40996
rect 32582 40944 32588 40996
rect 32640 40944 32646 40996
rect 34238 40944 34244 40996
rect 34296 40984 34302 40996
rect 34333 40987 34391 40993
rect 34333 40984 34345 40987
rect 34296 40956 34345 40984
rect 34296 40944 34302 40956
rect 34333 40953 34345 40956
rect 34379 40953 34391 40987
rect 34333 40947 34391 40953
rect 28500 40888 28672 40916
rect 28500 40876 28506 40888
rect 28810 40876 28816 40928
rect 28868 40916 28874 40928
rect 28997 40919 29055 40925
rect 28997 40916 29009 40919
rect 28868 40888 29009 40916
rect 28868 40876 28874 40888
rect 28997 40885 29009 40888
rect 29043 40885 29055 40919
rect 28997 40879 29055 40885
rect 30098 40876 30104 40928
rect 30156 40916 30162 40928
rect 31573 40919 31631 40925
rect 31573 40916 31585 40919
rect 30156 40888 31585 40916
rect 30156 40876 30162 40888
rect 31573 40885 31585 40888
rect 31619 40885 31631 40919
rect 31573 40879 31631 40885
rect 31846 40876 31852 40928
rect 31904 40916 31910 40928
rect 32769 40919 32827 40925
rect 32769 40916 32781 40919
rect 31904 40888 32781 40916
rect 31904 40876 31910 40888
rect 32769 40885 32781 40888
rect 32815 40885 32827 40919
rect 32769 40879 32827 40885
rect 33502 40876 33508 40928
rect 33560 40876 33566 40928
rect 36906 40876 36912 40928
rect 36964 40876 36970 40928
rect 41506 40876 41512 40928
rect 41564 40916 41570 40928
rect 41969 40919 42027 40925
rect 41969 40916 41981 40919
rect 41564 40888 41981 40916
rect 41564 40876 41570 40888
rect 41969 40885 41981 40888
rect 42015 40885 42027 40919
rect 41969 40879 42027 40885
rect 1104 40826 43884 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 43884 40826
rect 1104 40752 43884 40774
rect 12158 40672 12164 40724
rect 12216 40712 12222 40724
rect 12253 40715 12311 40721
rect 12253 40712 12265 40715
rect 12216 40684 12265 40712
rect 12216 40672 12222 40684
rect 12253 40681 12265 40684
rect 12299 40681 12311 40715
rect 12253 40675 12311 40681
rect 15194 40672 15200 40724
rect 15252 40712 15258 40724
rect 15838 40712 15844 40724
rect 15252 40684 15844 40712
rect 15252 40672 15258 40684
rect 15838 40672 15844 40684
rect 15896 40712 15902 40724
rect 16209 40715 16267 40721
rect 16209 40712 16221 40715
rect 15896 40684 16221 40712
rect 15896 40672 15902 40684
rect 16209 40681 16221 40684
rect 16255 40681 16267 40715
rect 16209 40675 16267 40681
rect 16408 40684 20300 40712
rect 8938 40644 8944 40656
rect 5920 40616 8944 40644
rect 5920 40585 5948 40616
rect 8938 40604 8944 40616
rect 8996 40644 9002 40656
rect 9214 40644 9220 40656
rect 8996 40616 9220 40644
rect 8996 40604 9002 40616
rect 9214 40604 9220 40616
rect 9272 40604 9278 40656
rect 15102 40604 15108 40656
rect 15160 40604 15166 40656
rect 5905 40579 5963 40585
rect 5905 40545 5917 40579
rect 5951 40545 5963 40579
rect 5905 40539 5963 40545
rect 7098 40536 7104 40588
rect 7156 40536 7162 40588
rect 9122 40536 9128 40588
rect 9180 40576 9186 40588
rect 9180 40548 10916 40576
rect 9180 40536 9186 40548
rect 5626 40468 5632 40520
rect 5684 40508 5690 40520
rect 6822 40508 6828 40520
rect 5684 40480 6828 40508
rect 5684 40468 5690 40480
rect 6822 40468 6828 40480
rect 6880 40468 6886 40520
rect 7116 40508 7144 40536
rect 9582 40508 9588 40520
rect 7116 40480 9588 40508
rect 9582 40468 9588 40480
rect 9640 40468 9646 40520
rect 10888 40517 10916 40548
rect 9769 40511 9827 40517
rect 9769 40508 9781 40511
rect 9692 40480 9781 40508
rect 6917 40443 6975 40449
rect 6917 40409 6929 40443
rect 6963 40440 6975 40443
rect 7006 40440 7012 40452
rect 6963 40412 7012 40440
rect 6963 40409 6975 40412
rect 6917 40403 6975 40409
rect 7006 40400 7012 40412
rect 7064 40400 7070 40452
rect 8754 40400 8760 40452
rect 8812 40440 8818 40452
rect 9125 40443 9183 40449
rect 9125 40440 9137 40443
rect 8812 40412 9137 40440
rect 8812 40400 8818 40412
rect 9125 40409 9137 40412
rect 9171 40409 9183 40443
rect 9125 40403 9183 40409
rect 5258 40332 5264 40384
rect 5316 40332 5322 40384
rect 5721 40375 5779 40381
rect 5721 40341 5733 40375
rect 5767 40372 5779 40375
rect 5994 40372 6000 40384
rect 5767 40344 6000 40372
rect 5767 40341 5779 40344
rect 5721 40335 5779 40341
rect 5994 40332 6000 40344
rect 6052 40332 6058 40384
rect 6457 40375 6515 40381
rect 6457 40341 6469 40375
rect 6503 40372 6515 40375
rect 6638 40372 6644 40384
rect 6503 40344 6644 40372
rect 6503 40341 6515 40344
rect 6457 40335 6515 40341
rect 6638 40332 6644 40344
rect 6696 40332 6702 40384
rect 6825 40375 6883 40381
rect 6825 40341 6837 40375
rect 6871 40372 6883 40375
rect 7190 40372 7196 40384
rect 6871 40344 7196 40372
rect 6871 40341 6883 40344
rect 6825 40335 6883 40341
rect 7190 40332 7196 40344
rect 7248 40332 7254 40384
rect 9030 40332 9036 40384
rect 9088 40372 9094 40384
rect 9692 40372 9720 40480
rect 9769 40477 9781 40480
rect 9815 40477 9827 40511
rect 9769 40471 9827 40477
rect 9861 40511 9919 40517
rect 9861 40477 9873 40511
rect 9907 40477 9919 40511
rect 9861 40471 9919 40477
rect 10873 40511 10931 40517
rect 10873 40477 10885 40511
rect 10919 40508 10931 40511
rect 12066 40508 12072 40520
rect 10919 40480 12072 40508
rect 10919 40477 10931 40480
rect 10873 40471 10931 40477
rect 9876 40384 9904 40471
rect 12066 40468 12072 40480
rect 12124 40468 12130 40520
rect 16408 40517 16436 40684
rect 17954 40604 17960 40656
rect 18012 40644 18018 40656
rect 18233 40647 18291 40653
rect 18233 40644 18245 40647
rect 18012 40616 18245 40644
rect 18012 40604 18018 40616
rect 18233 40613 18245 40616
rect 18279 40613 18291 40647
rect 20272 40644 20300 40684
rect 20346 40672 20352 40724
rect 20404 40672 20410 40724
rect 22462 40712 22468 40724
rect 20456 40684 22468 40712
rect 20456 40644 20484 40684
rect 22462 40672 22468 40684
rect 22520 40672 22526 40724
rect 22971 40715 23029 40721
rect 22971 40681 22983 40715
rect 23017 40712 23029 40715
rect 25222 40712 25228 40724
rect 23017 40684 25228 40712
rect 23017 40681 23029 40684
rect 22971 40675 23029 40681
rect 25222 40672 25228 40684
rect 25280 40672 25286 40724
rect 27614 40712 27620 40724
rect 26252 40684 27620 40712
rect 20272 40616 20484 40644
rect 18233 40607 18291 40613
rect 23382 40604 23388 40656
rect 23440 40644 23446 40656
rect 24854 40644 24860 40656
rect 23440 40616 24860 40644
rect 23440 40604 23446 40616
rect 24854 40604 24860 40616
rect 24912 40644 24918 40656
rect 26252 40644 26280 40684
rect 27614 40672 27620 40684
rect 27672 40672 27678 40724
rect 28902 40672 28908 40724
rect 28960 40712 28966 40724
rect 30285 40715 30343 40721
rect 30285 40712 30297 40715
rect 28960 40684 30297 40712
rect 28960 40672 28966 40684
rect 30285 40681 30297 40684
rect 30331 40681 30343 40715
rect 30285 40675 30343 40681
rect 32401 40715 32459 40721
rect 32401 40681 32413 40715
rect 32447 40712 32459 40715
rect 32490 40712 32496 40724
rect 32447 40684 32496 40712
rect 32447 40681 32459 40684
rect 32401 40675 32459 40681
rect 32490 40672 32496 40684
rect 32548 40672 32554 40724
rect 35069 40715 35127 40721
rect 35069 40681 35081 40715
rect 35115 40712 35127 40715
rect 35342 40712 35348 40724
rect 35115 40684 35348 40712
rect 35115 40681 35127 40684
rect 35069 40675 35127 40681
rect 35342 40672 35348 40684
rect 35400 40672 35406 40724
rect 36081 40715 36139 40721
rect 36081 40681 36093 40715
rect 36127 40712 36139 40715
rect 36906 40712 36912 40724
rect 36127 40684 36912 40712
rect 36127 40681 36139 40684
rect 36081 40675 36139 40681
rect 36906 40672 36912 40684
rect 36964 40672 36970 40724
rect 38470 40672 38476 40724
rect 38528 40672 38534 40724
rect 40589 40715 40647 40721
rect 40589 40681 40601 40715
rect 40635 40712 40647 40715
rect 40678 40712 40684 40724
rect 40635 40684 40684 40712
rect 40635 40681 40647 40684
rect 40589 40675 40647 40681
rect 40678 40672 40684 40684
rect 40736 40672 40742 40724
rect 24912 40616 26280 40644
rect 26329 40647 26387 40653
rect 24912 40604 24918 40616
rect 26329 40613 26341 40647
rect 26375 40613 26387 40647
rect 26329 40607 26387 40613
rect 16853 40579 16911 40585
rect 16853 40545 16865 40579
rect 16899 40576 16911 40579
rect 17218 40576 17224 40588
rect 16899 40548 17224 40576
rect 16899 40545 16911 40548
rect 16853 40539 16911 40545
rect 17218 40536 17224 40548
rect 17276 40536 17282 40588
rect 21082 40536 21088 40588
rect 21140 40576 21146 40588
rect 21177 40579 21235 40585
rect 21177 40576 21189 40579
rect 21140 40548 21189 40576
rect 21140 40536 21146 40548
rect 21177 40545 21189 40548
rect 21223 40545 21235 40579
rect 22278 40576 22284 40588
rect 21177 40539 21235 40545
rect 21284 40548 22284 40576
rect 16393 40511 16451 40517
rect 12406 40480 16344 40508
rect 11140 40443 11198 40449
rect 11140 40409 11152 40443
rect 11186 40440 11198 40443
rect 11698 40440 11704 40452
rect 11186 40412 11704 40440
rect 11186 40409 11198 40412
rect 11140 40403 11198 40409
rect 11698 40400 11704 40412
rect 11756 40400 11762 40452
rect 9088 40344 9720 40372
rect 9088 40332 9094 40344
rect 9858 40332 9864 40384
rect 9916 40372 9922 40384
rect 12406 40372 12434 40480
rect 14274 40400 14280 40452
rect 14332 40440 14338 40452
rect 14550 40440 14556 40452
rect 14332 40412 14556 40440
rect 14332 40400 14338 40412
rect 14550 40400 14556 40412
rect 14608 40400 14614 40452
rect 14642 40400 14648 40452
rect 14700 40400 14706 40452
rect 14734 40400 14740 40452
rect 14792 40440 14798 40452
rect 14829 40443 14887 40449
rect 14829 40440 14841 40443
rect 14792 40412 14841 40440
rect 14792 40400 14798 40412
rect 14829 40409 14841 40412
rect 14875 40440 14887 40443
rect 14918 40440 14924 40452
rect 14875 40412 14924 40440
rect 14875 40409 14887 40412
rect 14829 40403 14887 40409
rect 14918 40400 14924 40412
rect 14976 40400 14982 40452
rect 9916 40344 12434 40372
rect 16316 40372 16344 40480
rect 16393 40477 16405 40511
rect 16439 40477 16451 40511
rect 16393 40471 16451 40477
rect 17126 40468 17132 40520
rect 17184 40468 17190 40520
rect 20254 40468 20260 40520
rect 20312 40508 20318 40520
rect 21284 40508 21312 40548
rect 22278 40536 22284 40548
rect 22336 40536 22342 40588
rect 22554 40536 22560 40588
rect 22612 40576 22618 40588
rect 26234 40576 26240 40588
rect 22612 40548 24624 40576
rect 22612 40536 22618 40548
rect 20312 40480 21312 40508
rect 20312 40468 20318 40480
rect 21542 40468 21548 40520
rect 21600 40468 21606 40520
rect 23382 40468 23388 40520
rect 23440 40508 23446 40520
rect 24596 40517 24624 40548
rect 25700 40548 26240 40576
rect 23845 40511 23903 40517
rect 23845 40508 23857 40511
rect 23440 40480 23857 40508
rect 23440 40468 23446 40480
rect 23845 40477 23857 40480
rect 23891 40477 23903 40511
rect 23845 40471 23903 40477
rect 24029 40511 24087 40517
rect 24029 40477 24041 40511
rect 24075 40477 24087 40511
rect 24029 40471 24087 40477
rect 24581 40511 24639 40517
rect 24581 40477 24593 40511
rect 24627 40477 24639 40511
rect 24581 40471 24639 40477
rect 17788 40412 18368 40440
rect 17788 40372 17816 40412
rect 16316 40344 17816 40372
rect 18340 40372 18368 40412
rect 22278 40400 22284 40452
rect 22336 40400 22342 40452
rect 23474 40400 23480 40452
rect 23532 40440 23538 40452
rect 24044 40440 24072 40471
rect 24854 40468 24860 40520
rect 24912 40468 24918 40520
rect 25700 40517 25728 40548
rect 26234 40536 26240 40548
rect 26292 40536 26298 40588
rect 26344 40576 26372 40607
rect 28718 40604 28724 40656
rect 28776 40604 28782 40656
rect 30193 40647 30251 40653
rect 30193 40644 30205 40647
rect 28966 40616 30205 40644
rect 26510 40576 26516 40588
rect 26344 40548 26516 40576
rect 26510 40536 26516 40548
rect 26568 40576 26574 40588
rect 27433 40579 27491 40585
rect 27433 40576 27445 40579
rect 26568 40548 27445 40576
rect 26568 40536 26574 40548
rect 27433 40545 27445 40548
rect 27479 40545 27491 40579
rect 28736 40576 28764 40604
rect 28966 40588 28994 40616
rect 30193 40613 30205 40616
rect 30239 40644 30251 40647
rect 30558 40644 30564 40656
rect 30239 40616 30564 40644
rect 30239 40613 30251 40616
rect 30193 40607 30251 40613
rect 30558 40604 30564 40616
rect 30616 40644 30622 40656
rect 32582 40644 32588 40656
rect 30616 40616 32588 40644
rect 30616 40604 30622 40616
rect 32582 40604 32588 40616
rect 32640 40604 32646 40656
rect 35621 40647 35679 40653
rect 35621 40613 35633 40647
rect 35667 40613 35679 40647
rect 35621 40607 35679 40613
rect 28902 40576 28908 40588
rect 27433 40539 27491 40545
rect 28184 40548 28908 40576
rect 25685 40511 25743 40517
rect 25685 40477 25697 40511
rect 25731 40477 25743 40511
rect 25685 40471 25743 40477
rect 25958 40468 25964 40520
rect 26016 40468 26022 40520
rect 26970 40468 26976 40520
rect 27028 40468 27034 40520
rect 27062 40468 27068 40520
rect 27120 40468 27126 40520
rect 27890 40468 27896 40520
rect 27948 40468 27954 40520
rect 28074 40468 28080 40520
rect 28132 40468 28138 40520
rect 24762 40440 24768 40452
rect 23532 40412 24768 40440
rect 23532 40400 23538 40412
rect 24762 40400 24768 40412
rect 24820 40400 24826 40452
rect 24872 40440 24900 40468
rect 26053 40443 26111 40449
rect 26053 40440 26065 40443
rect 24872 40412 26065 40440
rect 26053 40409 26065 40412
rect 26099 40409 26111 40443
rect 26053 40403 26111 40409
rect 26142 40400 26148 40452
rect 26200 40449 26206 40452
rect 26200 40443 26228 40449
rect 26216 40440 26228 40443
rect 26216 40412 26924 40440
rect 26216 40409 26228 40412
rect 26200 40403 26228 40409
rect 26200 40400 26206 40403
rect 23842 40372 23848 40384
rect 18340 40344 23848 40372
rect 9916 40332 9922 40344
rect 23842 40332 23848 40344
rect 23900 40332 23906 40384
rect 23937 40375 23995 40381
rect 23937 40341 23949 40375
rect 23983 40372 23995 40375
rect 24118 40372 24124 40384
rect 23983 40344 24124 40372
rect 23983 40341 23995 40344
rect 23937 40335 23995 40341
rect 24118 40332 24124 40344
rect 24176 40332 24182 40384
rect 24210 40332 24216 40384
rect 24268 40372 24274 40384
rect 25958 40372 25964 40384
rect 24268 40344 25964 40372
rect 24268 40332 24274 40344
rect 25958 40332 25964 40344
rect 26016 40332 26022 40384
rect 26786 40332 26792 40384
rect 26844 40332 26850 40384
rect 26896 40372 26924 40412
rect 27154 40400 27160 40452
rect 27212 40400 27218 40452
rect 27246 40400 27252 40452
rect 27304 40449 27310 40452
rect 27304 40443 27353 40449
rect 27304 40409 27307 40443
rect 27341 40440 27353 40443
rect 27985 40443 28043 40449
rect 27985 40440 27997 40443
rect 27341 40412 27997 40440
rect 27341 40409 27353 40412
rect 27304 40403 27353 40409
rect 27985 40409 27997 40412
rect 28031 40409 28043 40443
rect 27985 40403 28043 40409
rect 27304 40400 27310 40403
rect 28184 40372 28212 40548
rect 28902 40536 28908 40548
rect 28960 40548 28994 40588
rect 30101 40579 30159 40585
rect 28960 40536 28966 40548
rect 30101 40545 30113 40579
rect 30147 40576 30159 40579
rect 30282 40576 30288 40588
rect 30147 40548 30288 40576
rect 30147 40545 30159 40548
rect 30101 40539 30159 40545
rect 30282 40536 30288 40548
rect 30340 40576 30346 40588
rect 31110 40576 31116 40588
rect 30340 40548 31116 40576
rect 30340 40536 30346 40548
rect 31110 40536 31116 40548
rect 31168 40536 31174 40588
rect 31662 40536 31668 40588
rect 31720 40576 31726 40588
rect 32493 40579 32551 40585
rect 32493 40576 32505 40579
rect 31720 40548 32505 40576
rect 31720 40536 31726 40548
rect 32493 40545 32505 40548
rect 32539 40545 32551 40579
rect 35161 40579 35219 40585
rect 32493 40539 32551 40545
rect 34164 40548 35112 40576
rect 28718 40468 28724 40520
rect 28776 40468 28782 40520
rect 28810 40468 28816 40520
rect 28868 40468 28874 40520
rect 29914 40468 29920 40520
rect 29972 40508 29978 40520
rect 30650 40508 30656 40520
rect 29972 40480 30656 40508
rect 29972 40468 29978 40480
rect 30650 40468 30656 40480
rect 30708 40468 30714 40520
rect 31297 40511 31355 40517
rect 31297 40477 31309 40511
rect 31343 40508 31355 40511
rect 31846 40508 31852 40520
rect 31343 40480 31852 40508
rect 31343 40477 31355 40480
rect 31297 40471 31355 40477
rect 31846 40468 31852 40480
rect 31904 40468 31910 40520
rect 31941 40511 31999 40517
rect 31941 40477 31953 40511
rect 31987 40477 31999 40511
rect 31941 40471 31999 40477
rect 29086 40400 29092 40452
rect 29144 40400 29150 40452
rect 29178 40400 29184 40452
rect 29236 40440 29242 40452
rect 31205 40443 31263 40449
rect 31205 40440 31217 40443
rect 29236 40412 31217 40440
rect 29236 40400 29242 40412
rect 31205 40409 31217 40412
rect 31251 40409 31263 40443
rect 31205 40403 31263 40409
rect 26896 40344 28212 40372
rect 28534 40332 28540 40384
rect 28592 40332 28598 40384
rect 29822 40332 29828 40384
rect 29880 40332 29886 40384
rect 30650 40332 30656 40384
rect 30708 40372 30714 40384
rect 31478 40372 31484 40384
rect 30708 40344 31484 40372
rect 30708 40332 30714 40344
rect 31478 40332 31484 40344
rect 31536 40372 31542 40384
rect 31956 40372 31984 40471
rect 32030 40468 32036 40520
rect 32088 40468 32094 40520
rect 33042 40468 33048 40520
rect 33100 40508 33106 40520
rect 33321 40511 33379 40517
rect 33321 40508 33333 40511
rect 33100 40480 33333 40508
rect 33100 40468 33106 40480
rect 33321 40477 33333 40480
rect 33367 40477 33379 40511
rect 33321 40471 33379 40477
rect 33505 40511 33563 40517
rect 33505 40477 33517 40511
rect 33551 40477 33563 40511
rect 33505 40471 33563 40477
rect 33520 40440 33548 40471
rect 33594 40468 33600 40520
rect 33652 40508 33658 40520
rect 34164 40517 34192 40548
rect 34149 40511 34207 40517
rect 34149 40508 34161 40511
rect 33652 40480 34161 40508
rect 33652 40468 33658 40480
rect 34149 40477 34161 40480
rect 34195 40477 34207 40511
rect 34149 40471 34207 40477
rect 34241 40511 34299 40517
rect 34241 40477 34253 40511
rect 34287 40508 34299 40511
rect 34790 40508 34796 40520
rect 34287 40480 34796 40508
rect 34287 40477 34299 40480
rect 34241 40471 34299 40477
rect 34790 40468 34796 40480
rect 34848 40508 34854 40520
rect 34885 40511 34943 40517
rect 34885 40508 34897 40511
rect 34848 40480 34897 40508
rect 34848 40468 34854 40480
rect 34885 40477 34897 40480
rect 34931 40477 34943 40511
rect 34885 40471 34943 40477
rect 34974 40468 34980 40520
rect 35032 40468 35038 40520
rect 35084 40508 35112 40548
rect 35161 40545 35173 40579
rect 35207 40576 35219 40579
rect 35636 40576 35664 40607
rect 35207 40548 35664 40576
rect 35207 40545 35219 40548
rect 35161 40539 35219 40545
rect 40126 40536 40132 40588
rect 40184 40536 40190 40588
rect 35894 40508 35900 40520
rect 35084 40480 35900 40508
rect 35894 40468 35900 40480
rect 35952 40468 35958 40520
rect 36173 40511 36231 40517
rect 36173 40477 36185 40511
rect 36219 40477 36231 40511
rect 36173 40471 36231 40477
rect 32784 40412 33548 40440
rect 33689 40443 33747 40449
rect 31536 40344 31984 40372
rect 31536 40332 31542 40344
rect 32122 40332 32128 40384
rect 32180 40372 32186 40384
rect 32784 40381 32812 40412
rect 33689 40409 33701 40443
rect 33735 40440 33747 40443
rect 33778 40440 33784 40452
rect 33735 40412 33784 40440
rect 33735 40409 33747 40412
rect 33689 40403 33747 40409
rect 33778 40400 33784 40412
rect 33836 40400 33842 40452
rect 35618 40400 35624 40452
rect 35676 40440 35682 40452
rect 36188 40440 36216 40471
rect 38378 40468 38384 40520
rect 38436 40468 38442 40520
rect 38562 40468 38568 40520
rect 38620 40468 38626 40520
rect 38838 40468 38844 40520
rect 38896 40508 38902 40520
rect 40221 40511 40279 40517
rect 40221 40508 40233 40511
rect 38896 40480 40233 40508
rect 38896 40468 38902 40480
rect 40221 40477 40233 40480
rect 40267 40477 40279 40511
rect 40221 40471 40279 40477
rect 41874 40468 41880 40520
rect 41932 40468 41938 40520
rect 35676 40412 36216 40440
rect 42144 40443 42202 40449
rect 35676 40400 35682 40412
rect 42144 40409 42156 40443
rect 42190 40440 42202 40443
rect 42610 40440 42616 40452
rect 42190 40412 42616 40440
rect 42190 40409 42202 40412
rect 42144 40403 42202 40409
rect 42610 40400 42616 40412
rect 42668 40400 42674 40452
rect 32769 40375 32827 40381
rect 32769 40372 32781 40375
rect 32180 40344 32781 40372
rect 32180 40332 32186 40344
rect 32769 40341 32781 40344
rect 32815 40341 32827 40375
rect 32769 40335 32827 40341
rect 42886 40332 42892 40384
rect 42944 40372 42950 40384
rect 43257 40375 43315 40381
rect 43257 40372 43269 40375
rect 42944 40344 43269 40372
rect 42944 40332 42950 40344
rect 43257 40341 43269 40344
rect 43303 40341 43315 40375
rect 43257 40335 43315 40341
rect 1104 40282 43884 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 43884 40282
rect 1104 40208 43884 40230
rect 5994 40128 6000 40180
rect 6052 40168 6058 40180
rect 7009 40171 7067 40177
rect 7009 40168 7021 40171
rect 6052 40140 7021 40168
rect 6052 40128 6058 40140
rect 7009 40137 7021 40140
rect 7055 40137 7067 40171
rect 7009 40131 7067 40137
rect 8386 40128 8392 40180
rect 8444 40128 8450 40180
rect 8849 40171 8907 40177
rect 8849 40137 8861 40171
rect 8895 40168 8907 40171
rect 9030 40168 9036 40180
rect 8895 40140 9036 40168
rect 8895 40137 8907 40140
rect 8849 40131 8907 40137
rect 9030 40128 9036 40140
rect 9088 40128 9094 40180
rect 11974 40128 11980 40180
rect 12032 40168 12038 40180
rect 12069 40171 12127 40177
rect 12069 40168 12081 40171
rect 12032 40140 12081 40168
rect 12032 40128 12038 40140
rect 12069 40137 12081 40140
rect 12115 40137 12127 40171
rect 12069 40131 12127 40137
rect 12158 40128 12164 40180
rect 12216 40128 12222 40180
rect 14277 40171 14335 40177
rect 14277 40137 14289 40171
rect 14323 40168 14335 40171
rect 14366 40168 14372 40180
rect 14323 40140 14372 40168
rect 14323 40137 14335 40140
rect 14277 40131 14335 40137
rect 14366 40128 14372 40140
rect 14424 40128 14430 40180
rect 23842 40168 23848 40180
rect 18340 40140 23848 40168
rect 4884 40103 4942 40109
rect 4884 40069 4896 40103
rect 4930 40100 4942 40103
rect 5258 40100 5264 40112
rect 4930 40072 5264 40100
rect 4930 40069 4942 40072
rect 4884 40063 4942 40069
rect 5258 40060 5264 40072
rect 5316 40060 5322 40112
rect 6822 40060 6828 40112
rect 6880 40100 6886 40112
rect 6917 40103 6975 40109
rect 6917 40100 6929 40103
rect 6880 40072 6929 40100
rect 6880 40060 6886 40072
rect 6917 40069 6929 40072
rect 6963 40069 6975 40103
rect 6917 40063 6975 40069
rect 8757 40103 8815 40109
rect 8757 40069 8769 40103
rect 8803 40100 8815 40103
rect 9858 40100 9864 40112
rect 8803 40072 9864 40100
rect 8803 40069 8815 40072
rect 8757 40063 8815 40069
rect 9858 40060 9864 40072
rect 9916 40060 9922 40112
rect 10042 40060 10048 40112
rect 10100 40100 10106 40112
rect 17037 40103 17095 40109
rect 10100 40072 10640 40100
rect 10100 40060 10106 40072
rect 9674 39992 9680 40044
rect 9732 40032 9738 40044
rect 10612 40041 10640 40072
rect 17037 40069 17049 40103
rect 17083 40100 17095 40103
rect 17083 40072 18092 40100
rect 17083 40069 17095 40072
rect 17037 40063 17095 40069
rect 10413 40035 10471 40041
rect 10413 40032 10425 40035
rect 9732 40004 10425 40032
rect 9732 39992 9738 40004
rect 10413 40001 10425 40004
rect 10459 40001 10471 40035
rect 10413 39995 10471 40001
rect 10597 40035 10655 40041
rect 10597 40001 10609 40035
rect 10643 40001 10655 40035
rect 10597 39995 10655 40001
rect 4617 39967 4675 39973
rect 4617 39933 4629 39967
rect 4663 39933 4675 39967
rect 4617 39927 4675 39933
rect 4632 39840 4660 39927
rect 7098 39924 7104 39976
rect 7156 39924 7162 39976
rect 8938 39924 8944 39976
rect 8996 39924 9002 39976
rect 9950 39924 9956 39976
rect 10008 39924 10014 39976
rect 10428 39896 10456 39995
rect 13722 39992 13728 40044
rect 13780 40032 13786 40044
rect 17221 40035 17279 40041
rect 13780 40004 14030 40032
rect 13780 39992 13786 40004
rect 17221 40001 17233 40035
rect 17267 40001 17279 40035
rect 17221 39995 17279 40001
rect 17313 40035 17371 40041
rect 17313 40001 17325 40035
rect 17359 40001 17371 40035
rect 17313 39995 17371 40001
rect 10686 39924 10692 39976
rect 10744 39924 10750 39976
rect 12253 39967 12311 39973
rect 12253 39933 12265 39967
rect 12299 39933 12311 39967
rect 12253 39927 12311 39933
rect 12268 39896 12296 39927
rect 12434 39924 12440 39976
rect 12492 39964 12498 39976
rect 13265 39967 13323 39973
rect 13265 39964 13277 39967
rect 12492 39936 13277 39964
rect 12492 39924 12498 39936
rect 13265 39933 13277 39936
rect 13311 39933 13323 39967
rect 13265 39927 13323 39933
rect 14274 39924 14280 39976
rect 14332 39924 14338 39976
rect 14292 39896 14320 39924
rect 10428 39868 14320 39896
rect 17037 39899 17095 39905
rect 17037 39865 17049 39899
rect 17083 39896 17095 39899
rect 17126 39896 17132 39908
rect 17083 39868 17132 39896
rect 17083 39865 17095 39868
rect 17037 39859 17095 39865
rect 17126 39856 17132 39868
rect 17184 39856 17190 39908
rect 17236 39896 17264 39995
rect 17328 39964 17356 39995
rect 17770 39992 17776 40044
rect 17828 39992 17834 40044
rect 18064 40032 18092 40072
rect 18230 40060 18236 40112
rect 18288 40100 18294 40112
rect 18340 40109 18368 40140
rect 23842 40128 23848 40140
rect 23900 40128 23906 40180
rect 24118 40128 24124 40180
rect 24176 40128 24182 40180
rect 24946 40128 24952 40180
rect 25004 40168 25010 40180
rect 26234 40168 26240 40180
rect 25004 40140 26240 40168
rect 25004 40128 25010 40140
rect 26234 40128 26240 40140
rect 26292 40128 26298 40180
rect 26405 40171 26463 40177
rect 26405 40137 26417 40171
rect 26451 40168 26463 40171
rect 27062 40168 27068 40180
rect 26451 40140 27068 40168
rect 26451 40137 26463 40140
rect 26405 40131 26463 40137
rect 27062 40128 27068 40140
rect 27120 40128 27126 40180
rect 27430 40128 27436 40180
rect 27488 40168 27494 40180
rect 28074 40168 28080 40180
rect 27488 40140 28080 40168
rect 27488 40128 27494 40140
rect 28074 40128 28080 40140
rect 28132 40168 28138 40180
rect 33686 40168 33692 40180
rect 28132 40140 33692 40168
rect 28132 40128 28138 40140
rect 33686 40128 33692 40140
rect 33744 40128 33750 40180
rect 34698 40128 34704 40180
rect 34756 40168 34762 40180
rect 35621 40171 35679 40177
rect 35621 40168 35633 40171
rect 34756 40140 35633 40168
rect 34756 40128 34762 40140
rect 35621 40137 35633 40140
rect 35667 40137 35679 40171
rect 35621 40131 35679 40137
rect 42610 40128 42616 40180
rect 42668 40128 42674 40180
rect 18325 40103 18383 40109
rect 18325 40100 18337 40103
rect 18288 40072 18337 40100
rect 18288 40060 18294 40072
rect 18325 40069 18337 40072
rect 18371 40069 18383 40103
rect 20254 40100 20260 40112
rect 18325 40063 18383 40069
rect 19306 40072 20260 40100
rect 18141 40035 18199 40041
rect 18141 40032 18153 40035
rect 18064 40004 18153 40032
rect 18141 40001 18153 40004
rect 18187 40032 18199 40035
rect 19306 40032 19334 40072
rect 20254 40060 20260 40072
rect 20312 40060 20318 40112
rect 24136 40100 24164 40128
rect 26605 40103 26663 40109
rect 24136 40072 26372 40100
rect 18187 40004 19334 40032
rect 18187 40001 18199 40004
rect 18141 39995 18199 40001
rect 22278 39992 22284 40044
rect 22336 39992 22342 40044
rect 22370 39992 22376 40044
rect 22428 39992 22434 40044
rect 22830 39992 22836 40044
rect 22888 40032 22894 40044
rect 23382 40032 23388 40044
rect 22888 40004 23388 40032
rect 22888 39992 22894 40004
rect 23382 39992 23388 40004
rect 23440 39992 23446 40044
rect 23845 40035 23903 40041
rect 23845 40001 23857 40035
rect 23891 40032 23903 40035
rect 24210 40032 24216 40044
rect 23891 40004 24216 40032
rect 23891 40001 23903 40004
rect 23845 39995 23903 40001
rect 24210 39992 24216 40004
rect 24268 39992 24274 40044
rect 24397 40035 24455 40041
rect 24397 40001 24409 40035
rect 24443 40032 24455 40035
rect 24670 40032 24676 40044
rect 24443 40004 24676 40032
rect 24443 40001 24455 40004
rect 24397 39995 24455 40001
rect 24670 39992 24676 40004
rect 24728 39992 24734 40044
rect 24762 39992 24768 40044
rect 24820 40032 24826 40044
rect 24949 40035 25007 40041
rect 24949 40032 24961 40035
rect 24820 40004 24961 40032
rect 24820 39992 24826 40004
rect 24949 40001 24961 40004
rect 24995 40032 25007 40035
rect 26142 40032 26148 40044
rect 24995 40004 26148 40032
rect 24995 40001 25007 40004
rect 24949 39995 25007 40001
rect 26142 39992 26148 40004
rect 26200 39992 26206 40044
rect 26344 40032 26372 40072
rect 26605 40069 26617 40103
rect 26651 40100 26663 40103
rect 27246 40100 27252 40112
rect 26651 40072 27252 40100
rect 26651 40069 26663 40072
rect 26605 40063 26663 40069
rect 27246 40060 27252 40072
rect 27304 40060 27310 40112
rect 28994 40100 29000 40112
rect 27540 40072 29000 40100
rect 27154 40032 27160 40044
rect 26344 40004 27160 40032
rect 18322 39964 18328 39976
rect 17328 39936 18328 39964
rect 18322 39924 18328 39936
rect 18380 39924 18386 39976
rect 23934 39924 23940 39976
rect 23992 39924 23998 39976
rect 24688 39964 24716 39992
rect 25038 39964 25044 39976
rect 24688 39936 25044 39964
rect 25038 39924 25044 39936
rect 25096 39924 25102 39976
rect 18230 39896 18236 39908
rect 17236 39868 18236 39896
rect 18230 39856 18236 39868
rect 18288 39856 18294 39908
rect 24578 39896 24584 39908
rect 22066 39868 24584 39896
rect 4614 39788 4620 39840
rect 4672 39828 4678 39840
rect 5534 39828 5540 39840
rect 4672 39800 5540 39828
rect 4672 39788 4678 39800
rect 5534 39788 5540 39800
rect 5592 39788 5598 39840
rect 6546 39788 6552 39840
rect 6604 39788 6610 39840
rect 11701 39831 11759 39837
rect 11701 39797 11713 39831
rect 11747 39828 11759 39831
rect 11790 39828 11796 39840
rect 11747 39800 11796 39828
rect 11747 39797 11759 39800
rect 11701 39791 11759 39797
rect 11790 39788 11796 39800
rect 11848 39788 11854 39840
rect 18874 39788 18880 39840
rect 18932 39828 18938 39840
rect 22066 39828 22094 39868
rect 24578 39856 24584 39868
rect 24636 39856 24642 39908
rect 18932 39800 22094 39828
rect 18932 39788 18938 39800
rect 25314 39788 25320 39840
rect 25372 39828 25378 39840
rect 26237 39831 26295 39837
rect 26237 39828 26249 39831
rect 25372 39800 26249 39828
rect 25372 39788 25378 39800
rect 26237 39797 26249 39800
rect 26283 39797 26295 39831
rect 26344 39828 26372 40004
rect 27154 39992 27160 40004
rect 27212 39992 27218 40044
rect 27062 39924 27068 39976
rect 27120 39964 27126 39976
rect 27540 39973 27568 40072
rect 28994 40060 29000 40072
rect 29052 40100 29058 40112
rect 29822 40100 29828 40112
rect 29052 40072 29828 40100
rect 29052 40060 29058 40072
rect 29822 40060 29828 40072
rect 29880 40060 29886 40112
rect 29917 40103 29975 40109
rect 29917 40069 29929 40103
rect 29963 40100 29975 40103
rect 30282 40100 30288 40112
rect 29963 40072 30288 40100
rect 29963 40069 29975 40072
rect 29917 40063 29975 40069
rect 30282 40060 30288 40072
rect 30340 40060 30346 40112
rect 33502 40100 33508 40112
rect 33428 40072 33508 40100
rect 27614 39992 27620 40044
rect 27672 39992 27678 40044
rect 27985 40035 28043 40041
rect 27985 40001 27997 40035
rect 28031 40032 28043 40035
rect 29178 40032 29184 40044
rect 28031 40004 29184 40032
rect 28031 40001 28043 40004
rect 27985 39995 28043 40001
rect 29178 39992 29184 40004
rect 29236 39992 29242 40044
rect 30190 39992 30196 40044
rect 30248 39992 30254 40044
rect 31018 39992 31024 40044
rect 31076 39992 31082 40044
rect 31478 39992 31484 40044
rect 31536 39992 31542 40044
rect 33428 40041 33456 40072
rect 33502 40060 33508 40072
rect 33560 40060 33566 40112
rect 34606 40100 34612 40112
rect 34440 40072 34612 40100
rect 33413 40035 33471 40041
rect 33413 40001 33425 40035
rect 33459 40001 33471 40035
rect 33413 39995 33471 40001
rect 34241 40035 34299 40041
rect 34241 40001 34253 40035
rect 34287 40032 34299 40035
rect 34440 40032 34468 40072
rect 34606 40060 34612 40072
rect 34664 40060 34670 40112
rect 38654 40060 38660 40112
rect 38712 40109 38718 40112
rect 38712 40103 38775 40109
rect 38712 40069 38729 40103
rect 38763 40069 38775 40103
rect 38712 40063 38775 40069
rect 38712 40060 38718 40063
rect 38838 40060 38844 40112
rect 38896 40100 38902 40112
rect 38933 40103 38991 40109
rect 38933 40100 38945 40103
rect 38896 40072 38945 40100
rect 38896 40060 38902 40072
rect 38933 40069 38945 40072
rect 38979 40069 38991 40103
rect 38933 40063 38991 40069
rect 42886 40060 42892 40112
rect 42944 40100 42950 40112
rect 42981 40103 43039 40109
rect 42981 40100 42993 40103
rect 42944 40072 42993 40100
rect 42944 40060 42950 40072
rect 42981 40069 42993 40072
rect 43027 40069 43039 40103
rect 42981 40063 43039 40069
rect 34514 40041 34520 40044
rect 34287 40004 34468 40032
rect 34287 40001 34299 40004
rect 34241 39995 34299 40001
rect 34508 39995 34520 40041
rect 34514 39992 34520 39995
rect 34572 39992 34578 40044
rect 27525 39967 27583 39973
rect 27525 39964 27537 39967
rect 27120 39936 27537 39964
rect 27120 39924 27126 39936
rect 27525 39933 27537 39936
rect 27571 39933 27583 39967
rect 27525 39927 27583 39933
rect 27893 39967 27951 39973
rect 27893 39933 27905 39967
rect 27939 39964 27951 39967
rect 28166 39964 28172 39976
rect 27939 39936 28172 39964
rect 27939 39933 27951 39936
rect 27893 39927 27951 39933
rect 28166 39924 28172 39936
rect 28224 39924 28230 39976
rect 28810 39924 28816 39976
rect 28868 39964 28874 39976
rect 32766 39964 32772 39976
rect 28868 39936 32772 39964
rect 28868 39924 28874 39936
rect 32766 39924 32772 39936
rect 32824 39924 32830 39976
rect 32858 39924 32864 39976
rect 32916 39924 32922 39976
rect 43070 39924 43076 39976
rect 43128 39924 43134 39976
rect 43162 39924 43168 39976
rect 43220 39924 43226 39976
rect 27246 39856 27252 39908
rect 27304 39896 27310 39908
rect 27304 39868 34284 39896
rect 27304 39856 27310 39868
rect 26421 39831 26479 39837
rect 26421 39828 26433 39831
rect 26344 39800 26433 39828
rect 26237 39791 26295 39797
rect 26421 39797 26433 39800
rect 26467 39797 26479 39831
rect 26421 39791 26479 39797
rect 26602 39788 26608 39840
rect 26660 39828 26666 39840
rect 27341 39831 27399 39837
rect 27341 39828 27353 39831
rect 26660 39800 27353 39828
rect 26660 39788 26666 39800
rect 27341 39797 27353 39800
rect 27387 39797 27399 39831
rect 27341 39791 27399 39797
rect 31665 39831 31723 39837
rect 31665 39797 31677 39831
rect 31711 39828 31723 39831
rect 31754 39828 31760 39840
rect 31711 39800 31760 39828
rect 31711 39797 31723 39800
rect 31665 39791 31723 39797
rect 31754 39788 31760 39800
rect 31812 39788 31818 39840
rect 34256 39828 34284 39868
rect 36446 39856 36452 39908
rect 36504 39896 36510 39908
rect 39298 39896 39304 39908
rect 36504 39868 39304 39896
rect 36504 39856 36510 39868
rect 39298 39856 39304 39868
rect 39356 39896 39362 39908
rect 40402 39896 40408 39908
rect 39356 39868 40408 39896
rect 39356 39856 39362 39868
rect 40402 39856 40408 39868
rect 40460 39856 40466 39908
rect 34422 39828 34428 39840
rect 34256 39800 34428 39828
rect 34422 39788 34428 39800
rect 34480 39788 34486 39840
rect 34606 39788 34612 39840
rect 34664 39828 34670 39840
rect 34974 39828 34980 39840
rect 34664 39800 34980 39828
rect 34664 39788 34670 39800
rect 34974 39788 34980 39800
rect 35032 39788 35038 39840
rect 38562 39788 38568 39840
rect 38620 39788 38626 39840
rect 38749 39831 38807 39837
rect 38749 39797 38761 39831
rect 38795 39828 38807 39831
rect 38930 39828 38936 39840
rect 38795 39800 38936 39828
rect 38795 39797 38807 39800
rect 38749 39791 38807 39797
rect 38930 39788 38936 39800
rect 38988 39828 38994 39840
rect 40126 39828 40132 39840
rect 38988 39800 40132 39828
rect 38988 39788 38994 39800
rect 40126 39788 40132 39800
rect 40184 39788 40190 39840
rect 1104 39738 43884 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 43884 39738
rect 1104 39664 43884 39686
rect 18322 39584 18328 39636
rect 18380 39584 18386 39636
rect 20993 39627 21051 39633
rect 20993 39624 21005 39627
rect 20088 39596 21005 39624
rect 6549 39491 6607 39497
rect 6549 39457 6561 39491
rect 6595 39488 6607 39491
rect 6730 39488 6736 39500
rect 6595 39460 6736 39488
rect 6595 39457 6607 39460
rect 6549 39451 6607 39457
rect 6730 39448 6736 39460
rect 6788 39448 6794 39500
rect 9950 39448 9956 39500
rect 10008 39488 10014 39500
rect 10008 39460 10640 39488
rect 10008 39448 10014 39460
rect 6638 39380 6644 39432
rect 6696 39380 6702 39432
rect 7374 39380 7380 39432
rect 7432 39420 7438 39432
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 7432 39392 9137 39420
rect 7432 39380 7438 39392
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9401 39423 9459 39429
rect 9401 39389 9413 39423
rect 9447 39420 9459 39423
rect 10410 39420 10416 39432
rect 9447 39392 10416 39420
rect 9447 39389 9459 39392
rect 9401 39383 9459 39389
rect 10410 39380 10416 39392
rect 10468 39380 10474 39432
rect 10612 39429 10640 39460
rect 16850 39448 16856 39500
rect 16908 39488 16914 39500
rect 17678 39488 17684 39500
rect 16908 39460 17684 39488
rect 16908 39448 16914 39460
rect 17678 39448 17684 39460
rect 17736 39488 17742 39500
rect 20088 39488 20116 39596
rect 20993 39593 21005 39596
rect 21039 39593 21051 39627
rect 20993 39587 21051 39593
rect 20162 39516 20168 39568
rect 20220 39556 20226 39568
rect 21008 39556 21036 39587
rect 21174 39584 21180 39636
rect 21232 39584 21238 39636
rect 23845 39627 23903 39633
rect 23845 39593 23857 39627
rect 23891 39593 23903 39627
rect 23845 39587 23903 39593
rect 23860 39556 23888 39587
rect 24026 39584 24032 39636
rect 24084 39584 24090 39636
rect 27614 39584 27620 39636
rect 27672 39584 27678 39636
rect 31662 39584 31668 39636
rect 31720 39624 31726 39636
rect 31757 39627 31815 39633
rect 31757 39624 31769 39627
rect 31720 39596 31769 39624
rect 31720 39584 31726 39596
rect 31757 39593 31769 39596
rect 31803 39593 31815 39627
rect 33042 39624 33048 39636
rect 31757 39587 31815 39593
rect 31956 39596 33048 39624
rect 28534 39556 28540 39568
rect 20220 39528 20944 39556
rect 21008 39528 22094 39556
rect 23860 39528 28540 39556
rect 20220 39516 20226 39528
rect 17736 39460 18460 39488
rect 20088 39460 20392 39488
rect 17736 39448 17742 39460
rect 18432 39432 18460 39460
rect 10597 39423 10655 39429
rect 10597 39389 10609 39423
rect 10643 39389 10655 39423
rect 10597 39383 10655 39389
rect 11330 39380 11336 39432
rect 11388 39420 11394 39432
rect 11609 39423 11667 39429
rect 11609 39420 11621 39423
rect 11388 39392 11621 39420
rect 11388 39380 11394 39392
rect 11609 39389 11621 39392
rect 11655 39389 11667 39423
rect 11609 39383 11667 39389
rect 15746 39380 15752 39432
rect 15804 39420 15810 39432
rect 16209 39423 16267 39429
rect 16209 39420 16221 39423
rect 15804 39392 16221 39420
rect 15804 39380 15810 39392
rect 16209 39389 16221 39392
rect 16255 39389 16267 39423
rect 16209 39383 16267 39389
rect 16393 39423 16451 39429
rect 16393 39389 16405 39423
rect 16439 39389 16451 39423
rect 16393 39383 16451 39389
rect 7098 39312 7104 39364
rect 7156 39312 7162 39364
rect 9493 39355 9551 39361
rect 9493 39321 9505 39355
rect 9539 39352 9551 39355
rect 10226 39352 10232 39364
rect 9539 39324 10232 39352
rect 9539 39321 9551 39324
rect 9493 39315 9551 39321
rect 10226 39312 10232 39324
rect 10284 39312 10290 39364
rect 11882 39312 11888 39364
rect 11940 39312 11946 39364
rect 14734 39312 14740 39364
rect 14792 39352 14798 39364
rect 16408 39352 16436 39383
rect 16482 39380 16488 39432
rect 16540 39420 16546 39432
rect 17497 39423 17555 39429
rect 17497 39420 17509 39423
rect 16540 39392 17509 39420
rect 16540 39380 16546 39392
rect 17497 39389 17509 39392
rect 17543 39389 17555 39423
rect 17497 39383 17555 39389
rect 17954 39380 17960 39432
rect 18012 39420 18018 39432
rect 18233 39423 18291 39429
rect 18233 39420 18245 39423
rect 18012 39392 18245 39420
rect 18012 39380 18018 39392
rect 18233 39389 18245 39392
rect 18279 39389 18291 39423
rect 18233 39383 18291 39389
rect 18414 39380 18420 39432
rect 18472 39380 18478 39432
rect 20070 39380 20076 39432
rect 20128 39420 20134 39432
rect 20364 39429 20392 39460
rect 20165 39423 20223 39429
rect 20165 39420 20177 39423
rect 20128 39392 20177 39420
rect 20128 39380 20134 39392
rect 20165 39389 20177 39392
rect 20211 39389 20223 39423
rect 20165 39383 20223 39389
rect 20349 39423 20407 39429
rect 20349 39389 20361 39423
rect 20395 39389 20407 39423
rect 20349 39383 20407 39389
rect 20806 39380 20812 39432
rect 20864 39380 20870 39432
rect 20916 39429 20944 39528
rect 22066 39488 22094 39528
rect 28534 39516 28540 39528
rect 28592 39516 28598 39568
rect 31956 39500 31984 39596
rect 33042 39584 33048 39596
rect 33100 39584 33106 39636
rect 34333 39627 34391 39633
rect 34333 39593 34345 39627
rect 34379 39624 34391 39627
rect 34514 39624 34520 39636
rect 34379 39596 34520 39624
rect 34379 39593 34391 39596
rect 34333 39587 34391 39593
rect 34514 39584 34520 39596
rect 34572 39584 34578 39636
rect 34882 39584 34888 39636
rect 34940 39624 34946 39636
rect 37737 39627 37795 39633
rect 34940 39596 37504 39624
rect 34940 39584 34946 39596
rect 32217 39559 32275 39565
rect 32217 39525 32229 39559
rect 32263 39525 32275 39559
rect 32217 39519 32275 39525
rect 27154 39488 27160 39500
rect 22066 39460 27160 39488
rect 27154 39448 27160 39460
rect 27212 39448 27218 39500
rect 27249 39491 27307 39497
rect 27249 39457 27261 39491
rect 27295 39488 27307 39491
rect 27338 39488 27344 39500
rect 27295 39460 27344 39488
rect 27295 39457 27307 39460
rect 27249 39451 27307 39457
rect 27338 39448 27344 39460
rect 27396 39488 27402 39500
rect 29086 39488 29092 39500
rect 27396 39460 29092 39488
rect 27396 39448 27402 39460
rect 29086 39448 29092 39460
rect 29144 39448 29150 39500
rect 31294 39488 31300 39500
rect 30392 39460 31300 39488
rect 20901 39423 20959 39429
rect 20901 39389 20913 39423
rect 20947 39389 20959 39423
rect 20901 39383 20959 39389
rect 21082 39380 21088 39432
rect 21140 39420 21146 39432
rect 22922 39420 22928 39432
rect 21140 39392 22928 39420
rect 21140 39380 21146 39392
rect 22922 39380 22928 39392
rect 22980 39380 22986 39432
rect 23106 39380 23112 39432
rect 23164 39380 23170 39432
rect 23750 39380 23756 39432
rect 23808 39380 23814 39432
rect 23845 39423 23903 39429
rect 23845 39389 23857 39423
rect 23891 39389 23903 39423
rect 23845 39383 23903 39389
rect 27433 39423 27491 39429
rect 27433 39389 27445 39423
rect 27479 39420 27491 39423
rect 27890 39420 27896 39432
rect 27479 39392 27896 39420
rect 27479 39389 27491 39392
rect 27433 39383 27491 39389
rect 14792 39324 16436 39352
rect 14792 39312 14798 39324
rect 10781 39287 10839 39293
rect 10781 39253 10793 39287
rect 10827 39284 10839 39287
rect 11974 39284 11980 39296
rect 10827 39256 11980 39284
rect 10827 39253 10839 39256
rect 10781 39247 10839 39253
rect 11974 39244 11980 39256
rect 12032 39244 12038 39296
rect 16298 39244 16304 39296
rect 16356 39244 16362 39296
rect 16408 39284 16436 39324
rect 16942 39312 16948 39364
rect 17000 39352 17006 39364
rect 23569 39355 23627 39361
rect 23569 39352 23581 39355
rect 17000 39324 20852 39352
rect 17000 39312 17006 39324
rect 17681 39287 17739 39293
rect 17681 39284 17693 39287
rect 16408 39256 17693 39284
rect 17681 39253 17693 39256
rect 17727 39284 17739 39287
rect 18046 39284 18052 39296
rect 17727 39256 18052 39284
rect 17727 39253 17739 39256
rect 17681 39247 17739 39253
rect 18046 39244 18052 39256
rect 18104 39244 18110 39296
rect 20254 39244 20260 39296
rect 20312 39244 20318 39296
rect 20824 39284 20852 39324
rect 21100 39324 23581 39352
rect 21100 39284 21128 39324
rect 23569 39321 23581 39324
rect 23615 39321 23627 39355
rect 23860 39352 23888 39383
rect 27890 39380 27896 39392
rect 27948 39380 27954 39432
rect 30098 39380 30104 39432
rect 30156 39380 30162 39432
rect 30392 39429 30420 39460
rect 31294 39448 31300 39460
rect 31352 39448 31358 39500
rect 31938 39448 31944 39500
rect 31996 39448 32002 39500
rect 32232 39488 32260 39519
rect 33778 39516 33784 39568
rect 33836 39556 33842 39568
rect 37476 39556 37504 39596
rect 37737 39593 37749 39627
rect 37783 39624 37795 39627
rect 38378 39624 38384 39636
rect 37783 39596 38384 39624
rect 37783 39593 37795 39596
rect 37737 39587 37795 39593
rect 38378 39584 38384 39596
rect 38436 39584 38442 39636
rect 38657 39627 38715 39633
rect 38657 39593 38669 39627
rect 38703 39624 38715 39627
rect 39206 39624 39212 39636
rect 38703 39596 39212 39624
rect 38703 39593 38715 39596
rect 38657 39587 38715 39593
rect 39206 39584 39212 39596
rect 39264 39584 39270 39636
rect 40954 39584 40960 39636
rect 41012 39624 41018 39636
rect 41414 39624 41420 39636
rect 41012 39596 41420 39624
rect 41012 39584 41018 39596
rect 41414 39584 41420 39596
rect 41472 39584 41478 39636
rect 39666 39556 39672 39568
rect 33836 39528 36584 39556
rect 33836 39516 33842 39528
rect 32232 39460 35020 39488
rect 30377 39423 30435 39429
rect 30377 39389 30389 39423
rect 30423 39389 30435 39423
rect 30377 39383 30435 39389
rect 30469 39423 30527 39429
rect 30469 39389 30481 39423
rect 30515 39389 30527 39423
rect 30469 39383 30527 39389
rect 23569 39315 23627 39321
rect 23768 39324 23888 39352
rect 20824 39256 21128 39284
rect 23014 39244 23020 39296
rect 23072 39284 23078 39296
rect 23768 39284 23796 39324
rect 24946 39312 24952 39364
rect 25004 39352 25010 39364
rect 28258 39352 28264 39364
rect 25004 39324 28264 39352
rect 25004 39312 25010 39324
rect 28258 39312 28264 39324
rect 28316 39312 28322 39364
rect 30484 39352 30512 39383
rect 31570 39380 31576 39432
rect 31628 39420 31634 39432
rect 32030 39420 32036 39432
rect 31628 39392 32036 39420
rect 31628 39380 31634 39392
rect 32030 39380 32036 39392
rect 32088 39380 32094 39432
rect 33873 39423 33931 39429
rect 33873 39389 33885 39423
rect 33919 39420 33931 39423
rect 34054 39420 34060 39432
rect 33919 39392 34060 39420
rect 33919 39389 33931 39392
rect 33873 39383 33931 39389
rect 34054 39380 34060 39392
rect 34112 39380 34118 39432
rect 34146 39380 34152 39432
rect 34204 39380 34210 39432
rect 34422 39380 34428 39432
rect 34480 39420 34486 39432
rect 34882 39420 34888 39432
rect 34480 39392 34888 39420
rect 34480 39380 34486 39392
rect 34882 39380 34888 39392
rect 34940 39380 34946 39432
rect 34992 39429 35020 39460
rect 36556 39429 36584 39528
rect 37476 39528 39672 39556
rect 36630 39448 36636 39500
rect 36688 39488 36694 39500
rect 36998 39488 37004 39500
rect 36688 39460 37004 39488
rect 36688 39448 36694 39460
rect 36998 39448 37004 39460
rect 37056 39488 37062 39500
rect 37056 39460 37412 39488
rect 37056 39448 37062 39460
rect 34977 39423 35035 39429
rect 34977 39389 34989 39423
rect 35023 39389 35035 39423
rect 34977 39383 35035 39389
rect 36541 39423 36599 39429
rect 36541 39389 36553 39423
rect 36587 39389 36599 39423
rect 36541 39383 36599 39389
rect 31754 39352 31760 39364
rect 30484 39324 31760 39352
rect 31754 39312 31760 39324
rect 31812 39312 31818 39364
rect 32769 39355 32827 39361
rect 32769 39321 32781 39355
rect 32815 39352 32827 39355
rect 32858 39352 32864 39364
rect 32815 39324 32864 39352
rect 32815 39321 32827 39324
rect 32769 39315 32827 39321
rect 32858 39312 32864 39324
rect 32916 39312 32922 39364
rect 34072 39352 34100 39380
rect 35345 39355 35403 39361
rect 35345 39352 35357 39355
rect 34072 39324 35357 39352
rect 35345 39321 35357 39324
rect 35391 39321 35403 39355
rect 35345 39315 35403 39321
rect 36078 39312 36084 39364
rect 36136 39352 36142 39364
rect 36265 39355 36323 39361
rect 36265 39352 36277 39355
rect 36136 39324 36277 39352
rect 36136 39312 36142 39324
rect 36265 39321 36277 39324
rect 36311 39321 36323 39355
rect 36556 39352 36584 39383
rect 37090 39380 37096 39432
rect 37148 39380 37154 39432
rect 37182 39380 37188 39432
rect 37240 39420 37246 39432
rect 37384 39429 37412 39460
rect 37369 39423 37427 39429
rect 37240 39392 37285 39420
rect 37240 39380 37246 39392
rect 37369 39389 37381 39423
rect 37415 39389 37427 39423
rect 37369 39383 37427 39389
rect 37476 39361 37504 39528
rect 39666 39516 39672 39528
rect 39724 39516 39730 39568
rect 37734 39448 37740 39500
rect 37792 39488 37798 39500
rect 37792 39460 39068 39488
rect 37792 39448 37798 39460
rect 37599 39423 37657 39429
rect 37599 39389 37611 39423
rect 37645 39420 37657 39423
rect 37918 39420 37924 39432
rect 37645 39392 37924 39420
rect 37645 39389 37657 39392
rect 37599 39383 37657 39389
rect 37918 39380 37924 39392
rect 37976 39380 37982 39432
rect 38930 39380 38936 39432
rect 38988 39380 38994 39432
rect 37461 39355 37519 39361
rect 36556 39324 37320 39352
rect 36265 39315 36323 39321
rect 37292 39296 37320 39324
rect 37461 39321 37473 39355
rect 37507 39321 37519 39355
rect 37461 39315 37519 39321
rect 38654 39312 38660 39364
rect 38712 39312 38718 39364
rect 38838 39312 38844 39364
rect 38896 39312 38902 39364
rect 23072 39256 23796 39284
rect 23072 39244 23078 39256
rect 30558 39244 30564 39296
rect 30616 39244 30622 39296
rect 33965 39287 34023 39293
rect 33965 39253 33977 39287
rect 34011 39284 34023 39287
rect 34698 39284 34704 39296
rect 34011 39256 34704 39284
rect 34011 39253 34023 39256
rect 33965 39247 34023 39253
rect 34698 39244 34704 39256
rect 34756 39244 34762 39296
rect 37274 39244 37280 39296
rect 37332 39244 37338 39296
rect 39040 39284 39068 39460
rect 40037 39423 40095 39429
rect 40037 39389 40049 39423
rect 40083 39420 40095 39423
rect 41782 39420 41788 39432
rect 40083 39392 41788 39420
rect 40083 39389 40095 39392
rect 40037 39383 40095 39389
rect 41782 39380 41788 39392
rect 41840 39380 41846 39432
rect 42702 39380 42708 39432
rect 42760 39420 42766 39432
rect 42889 39423 42947 39429
rect 42889 39420 42901 39423
rect 42760 39392 42901 39420
rect 42760 39380 42766 39392
rect 42889 39389 42901 39392
rect 42935 39389 42947 39423
rect 42889 39383 42947 39389
rect 39114 39312 39120 39364
rect 39172 39352 39178 39364
rect 40282 39355 40340 39361
rect 40282 39352 40294 39355
rect 39172 39324 40294 39352
rect 39172 39312 39178 39324
rect 40282 39321 40294 39324
rect 40328 39321 40340 39355
rect 40282 39315 40340 39321
rect 43165 39355 43223 39361
rect 43165 39321 43177 39355
rect 43211 39352 43223 39355
rect 43990 39352 43996 39364
rect 43211 39324 43996 39352
rect 43211 39321 43223 39324
rect 43165 39315 43223 39321
rect 43990 39312 43996 39324
rect 44048 39312 44054 39364
rect 41322 39284 41328 39296
rect 39040 39256 41328 39284
rect 41322 39244 41328 39256
rect 41380 39244 41386 39296
rect 41414 39244 41420 39296
rect 41472 39244 41478 39296
rect 1104 39194 43884 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 43884 39194
rect 1104 39120 43884 39142
rect 15749 39083 15807 39089
rect 15749 39049 15761 39083
rect 15795 39049 15807 39083
rect 15749 39043 15807 39049
rect 6730 39012 6736 39024
rect 5828 38984 6736 39012
rect 5828 38956 5856 38984
rect 6730 38972 6736 38984
rect 6788 39012 6794 39024
rect 6788 38984 7512 39012
rect 6788 38972 6794 38984
rect 5810 38904 5816 38956
rect 5868 38904 5874 38956
rect 5902 38904 5908 38956
rect 5960 38944 5966 38956
rect 5997 38947 6055 38953
rect 5997 38944 6009 38947
rect 5960 38916 6009 38944
rect 5960 38904 5966 38916
rect 5997 38913 6009 38916
rect 6043 38944 6055 38947
rect 6546 38944 6552 38956
rect 6043 38916 6552 38944
rect 6043 38913 6055 38916
rect 5997 38907 6055 38913
rect 6546 38904 6552 38916
rect 6604 38904 6610 38956
rect 7374 38904 7380 38956
rect 7432 38904 7438 38956
rect 7484 38953 7512 38984
rect 8754 38972 8760 39024
rect 8812 38972 8818 39024
rect 8941 39015 8999 39021
rect 8941 38981 8953 39015
rect 8987 39012 8999 39015
rect 8987 38984 10456 39012
rect 8987 38981 8999 38984
rect 8941 38975 8999 38981
rect 7469 38947 7527 38953
rect 7469 38913 7481 38947
rect 7515 38944 7527 38947
rect 8956 38944 8984 38975
rect 10428 38956 10456 38984
rect 12986 38972 12992 39024
rect 13044 39012 13050 39024
rect 13265 39015 13323 39021
rect 13265 39012 13277 39015
rect 13044 38984 13277 39012
rect 13044 38972 13050 38984
rect 13265 38981 13277 38984
rect 13311 38981 13323 39015
rect 15289 39015 15347 39021
rect 15289 39012 15301 39015
rect 13265 38975 13323 38981
rect 13372 38984 15301 39012
rect 7515 38916 8984 38944
rect 7515 38913 7527 38916
rect 7469 38907 7527 38913
rect 9950 38904 9956 38956
rect 10008 38904 10014 38956
rect 10410 38904 10416 38956
rect 10468 38944 10474 38956
rect 10689 38947 10747 38953
rect 10689 38944 10701 38947
rect 10468 38916 10701 38944
rect 10468 38904 10474 38916
rect 10689 38913 10701 38916
rect 10735 38913 10747 38947
rect 10689 38907 10747 38913
rect 11790 38904 11796 38956
rect 11848 38944 11854 38956
rect 11885 38947 11943 38953
rect 11885 38944 11897 38947
rect 11848 38916 11897 38944
rect 11848 38904 11854 38916
rect 11885 38913 11897 38916
rect 11931 38913 11943 38947
rect 12802 38944 12808 38956
rect 11885 38907 11943 38913
rect 11992 38916 12808 38944
rect 6730 38836 6736 38888
rect 6788 38876 6794 38888
rect 6917 38879 6975 38885
rect 6917 38876 6929 38879
rect 6788 38848 6929 38876
rect 6788 38836 6794 38848
rect 6917 38845 6929 38848
rect 6963 38845 6975 38879
rect 6917 38839 6975 38845
rect 10965 38879 11023 38885
rect 10965 38845 10977 38879
rect 11011 38876 11023 38879
rect 11992 38876 12020 38916
rect 12802 38904 12808 38916
rect 12860 38944 12866 38956
rect 13173 38947 13231 38953
rect 13173 38944 13185 38947
rect 12860 38916 13185 38944
rect 12860 38904 12866 38916
rect 13173 38913 13185 38916
rect 13219 38944 13231 38947
rect 13372 38944 13400 38984
rect 15289 38981 15301 38984
rect 15335 38981 15347 39015
rect 15764 39012 15792 39043
rect 16942 39040 16948 39092
rect 17000 39040 17006 39092
rect 17402 39040 17408 39092
rect 17460 39080 17466 39092
rect 18509 39083 18567 39089
rect 18509 39080 18521 39083
rect 17460 39052 18521 39080
rect 17460 39040 17466 39052
rect 18509 39049 18521 39052
rect 18555 39049 18567 39083
rect 18509 39043 18567 39049
rect 20070 39040 20076 39092
rect 20128 39040 20134 39092
rect 21082 39080 21088 39092
rect 20180 39052 21088 39080
rect 20180 39012 20208 39052
rect 21082 39040 21088 39052
rect 21140 39040 21146 39092
rect 21453 39083 21511 39089
rect 21453 39049 21465 39083
rect 21499 39080 21511 39083
rect 21542 39080 21548 39092
rect 21499 39052 21548 39080
rect 21499 39049 21511 39052
rect 21453 39043 21511 39049
rect 21542 39040 21548 39052
rect 21600 39040 21606 39092
rect 25133 39083 25191 39089
rect 25133 39080 25145 39083
rect 22066 39052 25145 39080
rect 15764 38984 20208 39012
rect 15289 38975 15347 38981
rect 20990 38972 20996 39024
rect 21048 39012 21054 39024
rect 22066 39012 22094 39052
rect 25133 39049 25145 39052
rect 25179 39049 25191 39083
rect 25133 39043 25191 39049
rect 26510 39040 26516 39092
rect 26568 39040 26574 39092
rect 27154 39040 27160 39092
rect 27212 39040 27218 39092
rect 32122 39080 32128 39092
rect 29012 39052 32128 39080
rect 26528 39012 26556 39040
rect 27982 39012 27988 39024
rect 21048 38984 22094 39012
rect 23216 38984 26464 39012
rect 26528 38984 27476 39012
rect 21048 38972 21054 38984
rect 13219 38916 13400 38944
rect 13449 38947 13507 38953
rect 13219 38913 13231 38916
rect 13173 38907 13231 38913
rect 13449 38913 13461 38947
rect 13495 38913 13507 38947
rect 13449 38907 13507 38913
rect 11011 38848 12020 38876
rect 12069 38879 12127 38885
rect 11011 38845 11023 38848
rect 10965 38839 11023 38845
rect 12069 38845 12081 38879
rect 12115 38845 12127 38879
rect 12069 38839 12127 38845
rect 11422 38768 11428 38820
rect 11480 38808 11486 38820
rect 12084 38808 12112 38839
rect 13078 38836 13084 38888
rect 13136 38876 13142 38888
rect 13464 38876 13492 38907
rect 13998 38904 14004 38956
rect 14056 38944 14062 38956
rect 14093 38947 14151 38953
rect 14093 38944 14105 38947
rect 14056 38916 14105 38944
rect 14056 38904 14062 38916
rect 14093 38913 14105 38916
rect 14139 38913 14151 38947
rect 14093 38907 14151 38913
rect 14829 38947 14887 38953
rect 14829 38913 14841 38947
rect 14875 38944 14887 38947
rect 15102 38944 15108 38956
rect 14875 38916 15108 38944
rect 14875 38913 14887 38916
rect 14829 38907 14887 38913
rect 15102 38904 15108 38916
rect 15160 38904 15166 38956
rect 15565 38947 15623 38953
rect 15565 38913 15577 38947
rect 15611 38913 15623 38947
rect 15565 38907 15623 38913
rect 14461 38879 14519 38885
rect 14461 38876 14473 38879
rect 13136 38848 14473 38876
rect 13136 38836 13142 38848
rect 14461 38845 14473 38848
rect 14507 38845 14519 38879
rect 15120 38876 15148 38904
rect 15381 38879 15439 38885
rect 15381 38876 15393 38879
rect 15120 38848 15393 38876
rect 14461 38839 14519 38845
rect 15381 38845 15393 38848
rect 15427 38845 15439 38879
rect 15381 38839 15439 38845
rect 12434 38808 12440 38820
rect 11480 38780 12112 38808
rect 11480 38768 11486 38780
rect 12406 38768 12440 38808
rect 12492 38768 12498 38820
rect 14734 38768 14740 38820
rect 14792 38808 14798 38820
rect 15580 38808 15608 38907
rect 16850 38904 16856 38956
rect 16908 38904 16914 38956
rect 17037 38947 17095 38953
rect 17037 38913 17049 38947
rect 17083 38913 17095 38947
rect 17037 38907 17095 38913
rect 18693 38947 18751 38953
rect 18693 38913 18705 38947
rect 18739 38913 18751 38947
rect 18693 38907 18751 38913
rect 16574 38836 16580 38888
rect 16632 38876 16638 38888
rect 17052 38876 17080 38907
rect 16632 38848 17080 38876
rect 18708 38876 18736 38907
rect 18782 38904 18788 38956
rect 18840 38904 18846 38956
rect 18874 38904 18880 38956
rect 18932 38904 18938 38956
rect 19426 38904 19432 38956
rect 19484 38904 19490 38956
rect 19518 38904 19524 38956
rect 19576 38944 19582 38956
rect 19889 38947 19947 38953
rect 19889 38944 19901 38947
rect 19576 38916 19901 38944
rect 19576 38904 19582 38916
rect 19889 38913 19901 38916
rect 19935 38944 19947 38947
rect 19978 38944 19984 38956
rect 19935 38916 19984 38944
rect 19935 38913 19947 38916
rect 19889 38907 19947 38913
rect 19978 38904 19984 38916
rect 20036 38904 20042 38956
rect 20809 38947 20867 38953
rect 20809 38913 20821 38947
rect 20855 38944 20867 38947
rect 21174 38944 21180 38956
rect 20855 38916 21180 38944
rect 20855 38913 20867 38916
rect 20809 38907 20867 38913
rect 21174 38904 21180 38916
rect 21232 38904 21238 38956
rect 21269 38947 21327 38953
rect 21269 38913 21281 38947
rect 21315 38944 21327 38947
rect 23216 38944 23244 38984
rect 21315 38916 23244 38944
rect 23293 38947 23351 38953
rect 21315 38913 21327 38916
rect 21269 38907 21327 38913
rect 23293 38913 23305 38947
rect 23339 38944 23351 38947
rect 23474 38944 23480 38956
rect 23339 38916 23480 38944
rect 23339 38913 23351 38916
rect 23293 38907 23351 38913
rect 23474 38904 23480 38916
rect 23532 38904 23538 38956
rect 24486 38904 24492 38956
rect 24544 38904 24550 38956
rect 24946 38904 24952 38956
rect 25004 38904 25010 38956
rect 26050 38904 26056 38956
rect 26108 38944 26114 38956
rect 26329 38947 26387 38953
rect 26329 38944 26341 38947
rect 26108 38916 26341 38944
rect 26108 38904 26114 38916
rect 26329 38913 26341 38916
rect 26375 38913 26387 38947
rect 26436 38944 26464 38984
rect 26605 38947 26663 38953
rect 26436 38916 26556 38944
rect 26329 38907 26387 38913
rect 19444 38876 19472 38904
rect 18708 38848 19472 38876
rect 19797 38879 19855 38885
rect 16632 38836 16638 38848
rect 19797 38845 19809 38879
rect 19843 38845 19855 38879
rect 19797 38839 19855 38845
rect 14792 38780 15608 38808
rect 14792 38768 14798 38780
rect 16298 38768 16304 38820
rect 16356 38808 16362 38820
rect 19812 38808 19840 38839
rect 20898 38836 20904 38888
rect 20956 38876 20962 38888
rect 21085 38879 21143 38885
rect 21085 38876 21097 38879
rect 20956 38848 21097 38876
rect 20956 38836 20962 38848
rect 21085 38845 21097 38848
rect 21131 38845 21143 38879
rect 21085 38839 21143 38845
rect 22833 38879 22891 38885
rect 22833 38845 22845 38879
rect 22879 38876 22891 38879
rect 22879 38848 23336 38876
rect 22879 38845 22891 38848
rect 22833 38839 22891 38845
rect 21174 38808 21180 38820
rect 16356 38780 19564 38808
rect 19812 38780 21180 38808
rect 16356 38768 16362 38780
rect 5905 38743 5963 38749
rect 5905 38709 5917 38743
rect 5951 38740 5963 38743
rect 7006 38740 7012 38752
rect 5951 38712 7012 38740
rect 5951 38709 5963 38712
rect 5905 38703 5963 38709
rect 7006 38700 7012 38712
rect 7064 38700 7070 38752
rect 7282 38700 7288 38752
rect 7340 38740 7346 38752
rect 8573 38743 8631 38749
rect 8573 38740 8585 38743
rect 7340 38712 8585 38740
rect 7340 38700 7346 38712
rect 8573 38709 8585 38712
rect 8619 38709 8631 38743
rect 8573 38703 8631 38709
rect 8757 38743 8815 38749
rect 8757 38709 8769 38743
rect 8803 38740 8815 38743
rect 9030 38740 9036 38752
rect 8803 38712 9036 38740
rect 8803 38709 8815 38712
rect 8757 38703 8815 38709
rect 9030 38700 9036 38712
rect 9088 38740 9094 38752
rect 12406 38740 12434 38768
rect 9088 38712 12434 38740
rect 13633 38743 13691 38749
rect 9088 38700 9094 38712
rect 13633 38709 13645 38743
rect 13679 38740 13691 38743
rect 14182 38740 14188 38752
rect 13679 38712 14188 38740
rect 13679 38709 13691 38712
rect 13633 38703 13691 38709
rect 14182 38700 14188 38712
rect 14240 38700 14246 38752
rect 14826 38700 14832 38752
rect 14884 38740 14890 38752
rect 19536 38749 19564 38780
rect 21174 38768 21180 38780
rect 21232 38768 21238 38820
rect 22741 38811 22799 38817
rect 22741 38777 22753 38811
rect 22787 38808 22799 38811
rect 23198 38808 23204 38820
rect 22787 38780 23204 38808
rect 22787 38777 22799 38780
rect 22741 38771 22799 38777
rect 23198 38768 23204 38780
rect 23256 38768 23262 38820
rect 23308 38808 23336 38848
rect 23382 38836 23388 38888
rect 23440 38836 23446 38888
rect 24857 38879 24915 38885
rect 24857 38845 24869 38879
rect 24903 38876 24915 38879
rect 26418 38876 26424 38888
rect 24903 38848 26424 38876
rect 24903 38845 24915 38848
rect 24857 38839 24915 38845
rect 26418 38836 26424 38848
rect 26476 38836 26482 38888
rect 25038 38808 25044 38820
rect 23308 38780 25044 38808
rect 25038 38768 25044 38780
rect 25096 38768 25102 38820
rect 26050 38768 26056 38820
rect 26108 38808 26114 38820
rect 26528 38808 26556 38916
rect 26605 38913 26617 38947
rect 26651 38944 26663 38947
rect 26970 38944 26976 38956
rect 26651 38916 26976 38944
rect 26651 38913 26663 38916
rect 26605 38907 26663 38913
rect 26970 38904 26976 38916
rect 27028 38944 27034 38956
rect 27448 38953 27476 38984
rect 27632 38984 27988 39012
rect 27632 38953 27660 38984
rect 27982 38972 27988 38984
rect 28040 38972 28046 39024
rect 28810 38972 28816 39024
rect 28868 39012 28874 39024
rect 28905 39015 28963 39021
rect 28905 39012 28917 39015
rect 28868 38984 28917 39012
rect 28868 38972 28874 38984
rect 28905 38981 28917 38984
rect 28951 38981 28963 39015
rect 28905 38975 28963 38981
rect 27341 38947 27399 38953
rect 27341 38944 27353 38947
rect 27028 38916 27353 38944
rect 27028 38904 27034 38916
rect 27341 38913 27353 38916
rect 27387 38913 27399 38947
rect 27341 38907 27399 38913
rect 27433 38947 27491 38953
rect 27433 38913 27445 38947
rect 27479 38913 27491 38947
rect 27433 38907 27491 38913
rect 27617 38947 27675 38953
rect 27617 38913 27629 38947
rect 27663 38913 27675 38947
rect 27617 38907 27675 38913
rect 27709 38947 27767 38953
rect 27709 38913 27721 38947
rect 27755 38913 27767 38947
rect 27709 38907 27767 38913
rect 27632 38808 27660 38907
rect 27724 38820 27752 38907
rect 27798 38904 27804 38956
rect 27856 38944 27862 38956
rect 28169 38947 28227 38953
rect 28169 38944 28181 38947
rect 27856 38916 28181 38944
rect 27856 38904 27862 38916
rect 28169 38913 28181 38916
rect 28215 38913 28227 38947
rect 28169 38907 28227 38913
rect 28353 38947 28411 38953
rect 28353 38913 28365 38947
rect 28399 38944 28411 38947
rect 28534 38944 28540 38956
rect 28399 38916 28540 38944
rect 28399 38913 28411 38916
rect 28353 38907 28411 38913
rect 28534 38904 28540 38916
rect 28592 38944 28598 38956
rect 29012 38944 29040 39052
rect 32122 39040 32128 39052
rect 32180 39040 32186 39092
rect 32766 39040 32772 39092
rect 32824 39080 32830 39092
rect 36722 39080 36728 39092
rect 32824 39052 36728 39080
rect 32824 39040 32830 39052
rect 30024 38984 30420 39012
rect 28592 38916 29040 38944
rect 29181 38947 29239 38953
rect 28592 38904 28598 38916
rect 29181 38913 29193 38947
rect 29227 38944 29239 38947
rect 30024 38944 30052 38984
rect 30392 38953 30420 38984
rect 31294 38972 31300 39024
rect 31352 39012 31358 39024
rect 33962 39012 33968 39024
rect 31352 38984 33968 39012
rect 31352 38972 31358 38984
rect 33962 38972 33968 38984
rect 34020 39012 34026 39024
rect 34149 39015 34207 39021
rect 34149 39012 34161 39015
rect 34020 38984 34161 39012
rect 34020 38972 34026 38984
rect 34149 38981 34161 38984
rect 34195 38981 34207 39015
rect 34149 38975 34207 38981
rect 36538 38972 36544 39024
rect 36596 38972 36602 39024
rect 36648 39021 36676 39052
rect 36722 39040 36728 39052
rect 36780 39040 36786 39092
rect 36909 39083 36967 39089
rect 36909 39049 36921 39083
rect 36955 39080 36967 39083
rect 37550 39080 37556 39092
rect 36955 39052 37556 39080
rect 36955 39049 36967 39052
rect 36909 39043 36967 39049
rect 37550 39040 37556 39052
rect 37608 39040 37614 39092
rect 37918 39080 37924 39092
rect 37660 39052 37924 39080
rect 36633 39015 36691 39021
rect 36633 38981 36645 39015
rect 36679 38981 36691 39015
rect 37660 39012 37688 39052
rect 37918 39040 37924 39052
rect 37976 39040 37982 39092
rect 38105 39083 38163 39089
rect 38105 39049 38117 39083
rect 38151 39080 38163 39083
rect 38930 39080 38936 39092
rect 38151 39052 38936 39080
rect 38151 39049 38163 39052
rect 38105 39043 38163 39049
rect 38930 39040 38936 39052
rect 38988 39040 38994 39092
rect 39114 39040 39120 39092
rect 39172 39040 39178 39092
rect 36633 38975 36691 38981
rect 36924 38984 37688 39012
rect 29227 38916 30052 38944
rect 30101 38947 30159 38953
rect 29227 38913 29239 38916
rect 29181 38907 29239 38913
rect 30101 38913 30113 38947
rect 30147 38913 30159 38947
rect 30101 38907 30159 38913
rect 30377 38947 30435 38953
rect 30377 38913 30389 38947
rect 30423 38944 30435 38947
rect 30466 38944 30472 38956
rect 30423 38916 30472 38944
rect 30423 38913 30435 38916
rect 30377 38907 30435 38913
rect 29638 38836 29644 38888
rect 29696 38836 29702 38888
rect 30116 38876 30144 38907
rect 30466 38904 30472 38916
rect 30524 38944 30530 38956
rect 31389 38947 31447 38953
rect 31389 38944 31401 38947
rect 30524 38916 31401 38944
rect 30524 38904 30530 38916
rect 31389 38913 31401 38916
rect 31435 38944 31447 38947
rect 31754 38944 31760 38956
rect 31435 38916 31760 38944
rect 31435 38913 31447 38916
rect 31389 38907 31447 38913
rect 31754 38904 31760 38916
rect 31812 38944 31818 38956
rect 32306 38944 32312 38956
rect 31812 38916 32312 38944
rect 31812 38904 31818 38916
rect 32306 38904 32312 38916
rect 32364 38904 32370 38956
rect 33137 38947 33195 38953
rect 33137 38913 33149 38947
rect 33183 38944 33195 38947
rect 33778 38944 33784 38956
rect 33183 38916 33784 38944
rect 33183 38913 33195 38916
rect 33137 38907 33195 38913
rect 33778 38904 33784 38916
rect 33836 38904 33842 38956
rect 33870 38904 33876 38956
rect 33928 38904 33934 38956
rect 34790 38904 34796 38956
rect 34848 38904 34854 38956
rect 36262 38904 36268 38956
rect 36320 38904 36326 38956
rect 36446 38953 36452 38956
rect 36413 38947 36452 38953
rect 36413 38913 36425 38947
rect 36413 38907 36452 38913
rect 36446 38904 36452 38907
rect 36504 38904 36510 38956
rect 36771 38947 36829 38953
rect 36771 38913 36783 38947
rect 36817 38944 36829 38947
rect 36924 38944 36952 38984
rect 37734 38972 37740 39024
rect 37792 38972 37798 39024
rect 36817 38916 36952 38944
rect 36817 38913 36829 38916
rect 36771 38907 36829 38913
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 37642 38953 37648 38956
rect 37461 38947 37519 38953
rect 37461 38944 37473 38947
rect 37424 38916 37473 38944
rect 37424 38904 37430 38916
rect 37461 38913 37473 38916
rect 37507 38913 37519 38947
rect 37461 38907 37519 38913
rect 37609 38947 37648 38953
rect 37609 38913 37621 38947
rect 37609 38907 37648 38913
rect 37642 38904 37648 38907
rect 37700 38904 37706 38956
rect 37829 38947 37887 38953
rect 37829 38913 37841 38947
rect 37875 38913 37887 38947
rect 37829 38907 37887 38913
rect 31481 38879 31539 38885
rect 29748 38848 30420 38876
rect 26108 38780 26464 38808
rect 26528 38780 27660 38808
rect 26108 38768 26114 38780
rect 15289 38743 15347 38749
rect 15289 38740 15301 38743
rect 14884 38712 15301 38740
rect 14884 38700 14890 38712
rect 15289 38709 15301 38712
rect 15335 38709 15347 38743
rect 15289 38703 15347 38709
rect 19521 38743 19579 38749
rect 19521 38709 19533 38743
rect 19567 38709 19579 38743
rect 19521 38703 19579 38709
rect 20254 38700 20260 38752
rect 20312 38740 20318 38752
rect 20901 38743 20959 38749
rect 20901 38740 20913 38743
rect 20312 38712 20913 38740
rect 20312 38700 20318 38712
rect 20901 38709 20913 38712
rect 20947 38709 20959 38743
rect 20901 38703 20959 38709
rect 22925 38743 22983 38749
rect 22925 38709 22937 38743
rect 22971 38740 22983 38743
rect 24210 38740 24216 38752
rect 22971 38712 24216 38740
rect 22971 38709 22983 38712
rect 22925 38703 22983 38709
rect 24210 38700 24216 38712
rect 24268 38700 24274 38752
rect 24578 38700 24584 38752
rect 24636 38700 24642 38752
rect 26142 38700 26148 38752
rect 26200 38700 26206 38752
rect 26436 38740 26464 38780
rect 27706 38768 27712 38820
rect 27764 38768 27770 38820
rect 28074 38768 28080 38820
rect 28132 38808 28138 38820
rect 28718 38808 28724 38820
rect 28132 38780 28724 38808
rect 28132 38768 28138 38780
rect 28718 38768 28724 38780
rect 28776 38808 28782 38820
rect 29089 38811 29147 38817
rect 29089 38808 29101 38811
rect 28776 38780 29101 38808
rect 28776 38768 28782 38780
rect 29089 38777 29101 38780
rect 29135 38808 29147 38811
rect 29748 38808 29776 38848
rect 29135 38780 29776 38808
rect 29135 38777 29147 38780
rect 29089 38771 29147 38777
rect 30098 38768 30104 38820
rect 30156 38808 30162 38820
rect 30285 38811 30343 38817
rect 30285 38808 30297 38811
rect 30156 38780 30297 38808
rect 30156 38768 30162 38780
rect 30285 38777 30297 38780
rect 30331 38777 30343 38811
rect 30392 38808 30420 38848
rect 31481 38845 31493 38879
rect 31527 38876 31539 38879
rect 31662 38876 31668 38888
rect 31527 38848 31668 38876
rect 31527 38845 31539 38848
rect 31481 38839 31539 38845
rect 31662 38836 31668 38848
rect 31720 38836 31726 38888
rect 32861 38879 32919 38885
rect 32861 38845 32873 38879
rect 32907 38845 32919 38879
rect 32861 38839 32919 38845
rect 35069 38879 35127 38885
rect 35069 38845 35081 38879
rect 35115 38876 35127 38879
rect 36078 38876 36084 38888
rect 35115 38848 36084 38876
rect 35115 38845 35127 38848
rect 35069 38839 35127 38845
rect 32674 38808 32680 38820
rect 30392 38780 32680 38808
rect 30285 38771 30343 38777
rect 32674 38768 32680 38780
rect 32732 38808 32738 38820
rect 32876 38808 32904 38839
rect 36078 38836 36084 38848
rect 36136 38836 36142 38888
rect 36906 38836 36912 38888
rect 36964 38876 36970 38888
rect 37844 38876 37872 38907
rect 37918 38904 37924 38956
rect 37976 38953 37982 38956
rect 37976 38944 37984 38953
rect 37976 38916 38021 38944
rect 37976 38907 37984 38916
rect 37976 38904 37982 38907
rect 38562 38904 38568 38956
rect 38620 38944 38626 38956
rect 39025 38947 39083 38953
rect 39025 38944 39037 38947
rect 38620 38916 39037 38944
rect 38620 38904 38626 38916
rect 39025 38913 39037 38916
rect 39071 38913 39083 38947
rect 39025 38907 39083 38913
rect 39206 38904 39212 38956
rect 39264 38904 39270 38956
rect 42978 38904 42984 38956
rect 43036 38904 43042 38956
rect 39758 38876 39764 38888
rect 36964 38848 39764 38876
rect 36964 38836 36970 38848
rect 39758 38836 39764 38848
rect 39816 38836 39822 38888
rect 42702 38836 42708 38888
rect 42760 38876 42766 38888
rect 43073 38879 43131 38885
rect 43073 38876 43085 38879
rect 42760 38848 43085 38876
rect 42760 38836 42766 38848
rect 43073 38845 43085 38848
rect 43119 38845 43131 38879
rect 43073 38839 43131 38845
rect 43162 38836 43168 38888
rect 43220 38836 43226 38888
rect 32732 38780 32904 38808
rect 32732 38768 32738 38780
rect 34698 38768 34704 38820
rect 34756 38808 34762 38820
rect 34885 38811 34943 38817
rect 34885 38808 34897 38811
rect 34756 38780 34897 38808
rect 34756 38768 34762 38780
rect 34885 38777 34897 38780
rect 34931 38777 34943 38811
rect 34885 38771 34943 38777
rect 36722 38768 36728 38820
rect 36780 38808 36786 38820
rect 39206 38808 39212 38820
rect 36780 38780 39212 38808
rect 36780 38768 36786 38780
rect 39206 38768 39212 38780
rect 39264 38768 39270 38820
rect 28169 38743 28227 38749
rect 28169 38740 28181 38743
rect 26436 38712 28181 38740
rect 28169 38709 28181 38712
rect 28215 38709 28227 38743
rect 28169 38703 28227 38709
rect 28994 38700 29000 38752
rect 29052 38700 29058 38752
rect 31294 38700 31300 38752
rect 31352 38740 31358 38752
rect 31389 38743 31447 38749
rect 31389 38740 31401 38743
rect 31352 38712 31401 38740
rect 31352 38700 31358 38712
rect 31389 38709 31401 38712
rect 31435 38709 31447 38743
rect 31389 38703 31447 38709
rect 31757 38743 31815 38749
rect 31757 38709 31769 38743
rect 31803 38740 31815 38743
rect 33042 38740 33048 38752
rect 31803 38712 33048 38740
rect 31803 38709 31815 38712
rect 31757 38703 31815 38709
rect 33042 38700 33048 38712
rect 33100 38700 33106 38752
rect 35253 38743 35311 38749
rect 35253 38709 35265 38743
rect 35299 38740 35311 38743
rect 35526 38740 35532 38752
rect 35299 38712 35532 38740
rect 35299 38709 35311 38712
rect 35253 38703 35311 38709
rect 35526 38700 35532 38712
rect 35584 38700 35590 38752
rect 37182 38700 37188 38752
rect 37240 38740 37246 38752
rect 40954 38740 40960 38752
rect 37240 38712 40960 38740
rect 37240 38700 37246 38712
rect 40954 38700 40960 38712
rect 41012 38700 41018 38752
rect 42610 38700 42616 38752
rect 42668 38700 42674 38752
rect 1104 38650 43884 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 43884 38650
rect 1104 38576 43884 38598
rect 12342 38496 12348 38548
rect 12400 38536 12406 38548
rect 14461 38539 14519 38545
rect 14461 38536 14473 38539
rect 12400 38508 14473 38536
rect 12400 38496 12406 38508
rect 14461 38505 14473 38508
rect 14507 38505 14519 38539
rect 17681 38539 17739 38545
rect 17681 38536 17693 38539
rect 14461 38499 14519 38505
rect 14568 38508 17693 38536
rect 14274 38468 14280 38480
rect 13004 38440 14280 38468
rect 7024 38372 7604 38400
rect 7024 38344 7052 38372
rect 5810 38292 5816 38344
rect 5868 38292 5874 38344
rect 5902 38292 5908 38344
rect 5960 38292 5966 38344
rect 7006 38292 7012 38344
rect 7064 38292 7070 38344
rect 7101 38335 7159 38341
rect 7101 38301 7113 38335
rect 7147 38332 7159 38335
rect 7190 38332 7196 38344
rect 7147 38304 7196 38332
rect 7147 38301 7159 38304
rect 7101 38295 7159 38301
rect 7190 38292 7196 38304
rect 7248 38292 7254 38344
rect 7576 38341 7604 38372
rect 10134 38360 10140 38412
rect 10192 38360 10198 38412
rect 13004 38409 13032 38440
rect 14274 38428 14280 38440
rect 14332 38468 14338 38480
rect 14568 38468 14596 38508
rect 17681 38505 17693 38508
rect 17727 38536 17739 38539
rect 17954 38536 17960 38548
rect 17727 38508 17960 38536
rect 17727 38505 17739 38508
rect 17681 38499 17739 38505
rect 17954 38496 17960 38508
rect 18012 38496 18018 38548
rect 19429 38539 19487 38545
rect 19429 38505 19441 38539
rect 19475 38536 19487 38539
rect 19518 38536 19524 38548
rect 19475 38508 19524 38536
rect 19475 38505 19487 38508
rect 19429 38499 19487 38505
rect 19518 38496 19524 38508
rect 19576 38496 19582 38548
rect 19797 38539 19855 38545
rect 19797 38505 19809 38539
rect 19843 38536 19855 38539
rect 19886 38536 19892 38548
rect 19843 38508 19892 38536
rect 19843 38505 19855 38508
rect 19797 38499 19855 38505
rect 19886 38496 19892 38508
rect 19944 38496 19950 38548
rect 19978 38496 19984 38548
rect 20036 38536 20042 38548
rect 20257 38539 20315 38545
rect 20257 38536 20269 38539
rect 20036 38508 20269 38536
rect 20036 38496 20042 38508
rect 20257 38505 20269 38508
rect 20303 38505 20315 38539
rect 20717 38539 20775 38545
rect 20257 38499 20315 38505
rect 20364 38508 20668 38536
rect 14332 38440 14596 38468
rect 14921 38471 14979 38477
rect 14332 38428 14338 38440
rect 14921 38437 14933 38471
rect 14967 38468 14979 38471
rect 20364 38468 20392 38508
rect 14967 38440 20392 38468
rect 20640 38468 20668 38508
rect 20717 38505 20729 38539
rect 20763 38536 20775 38539
rect 20806 38536 20812 38548
rect 20763 38508 20812 38536
rect 20763 38505 20775 38508
rect 20717 38499 20775 38505
rect 20806 38496 20812 38508
rect 20864 38496 20870 38548
rect 21174 38496 21180 38548
rect 21232 38496 21238 38548
rect 21358 38496 21364 38548
rect 21416 38496 21422 38548
rect 23934 38496 23940 38548
rect 23992 38496 23998 38548
rect 24854 38496 24860 38548
rect 24912 38496 24918 38548
rect 36909 38539 36967 38545
rect 32140 38508 36860 38536
rect 23201 38471 23259 38477
rect 20640 38440 21496 38468
rect 14967 38437 14979 38440
rect 14921 38431 14979 38437
rect 12989 38403 13047 38409
rect 12406 38372 12848 38400
rect 7561 38335 7619 38341
rect 7561 38301 7573 38335
rect 7607 38301 7619 38335
rect 7561 38295 7619 38301
rect 7926 38292 7932 38344
rect 7984 38292 7990 38344
rect 8110 38292 8116 38344
rect 8168 38292 8174 38344
rect 8754 38292 8760 38344
rect 8812 38332 8818 38344
rect 9217 38335 9275 38341
rect 9217 38332 9229 38335
rect 8812 38304 9229 38332
rect 8812 38292 8818 38304
rect 9217 38301 9229 38304
rect 9263 38301 9275 38335
rect 9217 38295 9275 38301
rect 10321 38335 10379 38341
rect 10321 38301 10333 38335
rect 10367 38301 10379 38335
rect 10321 38295 10379 38301
rect 6178 38224 6184 38276
rect 6236 38264 6242 38276
rect 6549 38267 6607 38273
rect 6549 38264 6561 38267
rect 6236 38236 6561 38264
rect 6236 38224 6242 38236
rect 6549 38233 6561 38236
rect 6595 38233 6607 38267
rect 10336 38264 10364 38295
rect 11146 38292 11152 38344
rect 11204 38332 11210 38344
rect 11517 38335 11575 38341
rect 11517 38332 11529 38335
rect 11204 38304 11529 38332
rect 11204 38292 11210 38304
rect 11517 38301 11529 38304
rect 11563 38301 11575 38335
rect 11517 38295 11575 38301
rect 11885 38335 11943 38341
rect 11885 38301 11897 38335
rect 11931 38332 11943 38335
rect 12406 38332 12434 38372
rect 11931 38304 12434 38332
rect 11931 38301 11943 38304
rect 11885 38295 11943 38301
rect 10336 38236 11928 38264
rect 6549 38227 6607 38233
rect 6089 38199 6147 38205
rect 6089 38165 6101 38199
rect 6135 38196 6147 38199
rect 8202 38196 8208 38208
rect 6135 38168 8208 38196
rect 6135 38165 6147 38168
rect 6089 38159 6147 38165
rect 8202 38156 8208 38168
rect 8260 38156 8266 38208
rect 11900 38196 11928 38236
rect 11974 38224 11980 38276
rect 12032 38264 12038 38276
rect 12069 38267 12127 38273
rect 12069 38264 12081 38267
rect 12032 38236 12081 38264
rect 12032 38224 12038 38236
rect 12069 38233 12081 38236
rect 12115 38233 12127 38267
rect 12618 38264 12624 38276
rect 12069 38227 12127 38233
rect 12406 38236 12624 38264
rect 12406 38196 12434 38236
rect 12618 38224 12624 38236
rect 12676 38224 12682 38276
rect 11900 38168 12434 38196
rect 12820 38196 12848 38372
rect 12989 38369 13001 38403
rect 13035 38369 13047 38403
rect 12989 38363 13047 38369
rect 13081 38403 13139 38409
rect 13081 38369 13093 38403
rect 13127 38400 13139 38403
rect 14090 38400 14096 38412
rect 13127 38372 14096 38400
rect 13127 38369 13139 38372
rect 13081 38363 13139 38369
rect 14090 38360 14096 38372
rect 14148 38360 14154 38412
rect 14645 38403 14703 38409
rect 14645 38369 14657 38403
rect 14691 38400 14703 38403
rect 15102 38400 15108 38412
rect 14691 38372 15108 38400
rect 14691 38369 14703 38372
rect 14645 38363 14703 38369
rect 15102 38360 15108 38372
rect 15160 38360 15166 38412
rect 16850 38400 16856 38412
rect 16224 38372 16856 38400
rect 13446 38292 13452 38344
rect 13504 38292 13510 38344
rect 14108 38332 14136 38360
rect 14108 38304 14688 38332
rect 12894 38224 12900 38276
rect 12952 38264 12958 38276
rect 14461 38267 14519 38273
rect 14461 38264 14473 38267
rect 12952 38236 14473 38264
rect 12952 38224 12958 38236
rect 14461 38233 14473 38236
rect 14507 38233 14519 38267
rect 14660 38264 14688 38304
rect 14734 38292 14740 38344
rect 14792 38292 14798 38344
rect 16224 38341 16252 38372
rect 16850 38360 16856 38372
rect 16908 38400 16914 38412
rect 17126 38400 17132 38412
rect 16908 38372 17132 38400
rect 16908 38360 16914 38372
rect 17126 38360 17132 38372
rect 17184 38360 17190 38412
rect 18785 38403 18843 38409
rect 18785 38369 18797 38403
rect 18831 38400 18843 38403
rect 18831 38372 20208 38400
rect 18831 38369 18843 38372
rect 18785 38363 18843 38369
rect 16117 38335 16175 38341
rect 16117 38301 16129 38335
rect 16163 38301 16175 38335
rect 16117 38295 16175 38301
rect 16209 38335 16267 38341
rect 16209 38301 16221 38335
rect 16255 38301 16267 38335
rect 16209 38295 16267 38301
rect 16132 38264 16160 38295
rect 16390 38292 16396 38344
rect 16448 38292 16454 38344
rect 16482 38292 16488 38344
rect 16540 38292 16546 38344
rect 17497 38335 17555 38341
rect 17497 38332 17509 38335
rect 16868 38304 17509 38332
rect 16868 38276 16896 38304
rect 17497 38301 17509 38304
rect 17543 38301 17555 38335
rect 17497 38295 17555 38301
rect 17678 38292 17684 38344
rect 17736 38292 17742 38344
rect 18690 38292 18696 38344
rect 18748 38292 18754 38344
rect 18874 38292 18880 38344
rect 18932 38292 18938 38344
rect 19705 38335 19763 38341
rect 19705 38301 19717 38335
rect 19751 38301 19763 38335
rect 19705 38295 19763 38301
rect 16850 38264 16856 38276
rect 14660 38236 16856 38264
rect 14461 38227 14519 38233
rect 16850 38224 16856 38236
rect 16908 38224 16914 38276
rect 13078 38196 13084 38208
rect 12820 38168 13084 38196
rect 13078 38156 13084 38168
rect 13136 38156 13142 38208
rect 13262 38156 13268 38208
rect 13320 38156 13326 38208
rect 13354 38156 13360 38208
rect 13412 38156 13418 38208
rect 13725 38199 13783 38205
rect 13725 38165 13737 38199
rect 13771 38196 13783 38199
rect 13814 38196 13820 38208
rect 13771 38168 13820 38196
rect 13771 38165 13783 38168
rect 13725 38159 13783 38165
rect 13814 38156 13820 38168
rect 13872 38156 13878 38208
rect 16666 38156 16672 38208
rect 16724 38156 16730 38208
rect 17865 38199 17923 38205
rect 17865 38165 17877 38199
rect 17911 38196 17923 38199
rect 19334 38196 19340 38208
rect 17911 38168 19340 38196
rect 17911 38165 17923 38168
rect 17865 38159 17923 38165
rect 19334 38156 19340 38168
rect 19392 38156 19398 38208
rect 19720 38196 19748 38295
rect 19794 38292 19800 38344
rect 19852 38292 19858 38344
rect 19886 38224 19892 38276
rect 19944 38264 19950 38276
rect 20070 38264 20076 38276
rect 19944 38236 20076 38264
rect 19944 38224 19950 38236
rect 20070 38224 20076 38236
rect 20128 38224 20134 38276
rect 20180 38264 20208 38372
rect 20346 38360 20352 38412
rect 20404 38400 20410 38412
rect 20441 38403 20499 38409
rect 20441 38400 20453 38403
rect 20404 38372 20453 38400
rect 20404 38360 20410 38372
rect 20441 38369 20453 38372
rect 20487 38400 20499 38403
rect 20487 38372 21404 38400
rect 20487 38369 20499 38372
rect 20441 38363 20499 38369
rect 20254 38292 20260 38344
rect 20312 38292 20318 38344
rect 20533 38335 20591 38341
rect 20533 38301 20545 38335
rect 20579 38326 20591 38335
rect 20622 38326 20628 38344
rect 20579 38301 20628 38326
rect 20533 38298 20628 38301
rect 20533 38295 20591 38298
rect 20622 38292 20628 38298
rect 20680 38292 20686 38344
rect 21376 38341 21404 38372
rect 21361 38335 21419 38341
rect 21361 38301 21373 38335
rect 21407 38301 21419 38335
rect 21468 38332 21496 38440
rect 23201 38437 23213 38471
rect 23247 38468 23259 38471
rect 23247 38440 24900 38468
rect 23247 38437 23259 38440
rect 23201 38431 23259 38437
rect 21545 38403 21603 38409
rect 21545 38369 21557 38403
rect 21591 38400 21603 38403
rect 23014 38400 23020 38412
rect 21591 38372 23020 38400
rect 21591 38369 21603 38372
rect 21545 38363 21603 38369
rect 23014 38360 23020 38372
rect 23072 38360 23078 38412
rect 24872 38409 24900 38440
rect 25866 38428 25872 38480
rect 25924 38468 25930 38480
rect 28353 38471 28411 38477
rect 28353 38468 28365 38471
rect 25924 38440 28365 38468
rect 25924 38428 25930 38440
rect 28353 38437 28365 38440
rect 28399 38468 28411 38471
rect 28994 38468 29000 38480
rect 28399 38440 29000 38468
rect 28399 38437 28411 38440
rect 28353 38431 28411 38437
rect 28994 38428 29000 38440
rect 29052 38428 29058 38480
rect 30377 38471 30435 38477
rect 30377 38437 30389 38471
rect 30423 38468 30435 38471
rect 31018 38468 31024 38480
rect 30423 38440 31024 38468
rect 30423 38437 30435 38440
rect 30377 38431 30435 38437
rect 31018 38428 31024 38440
rect 31076 38468 31082 38480
rect 31938 38468 31944 38480
rect 31076 38440 31944 38468
rect 31076 38428 31082 38440
rect 31938 38428 31944 38440
rect 31996 38428 32002 38480
rect 23753 38403 23811 38409
rect 23753 38369 23765 38403
rect 23799 38369 23811 38403
rect 23753 38363 23811 38369
rect 24857 38403 24915 38409
rect 24857 38369 24869 38403
rect 24903 38369 24915 38403
rect 27249 38403 27307 38409
rect 24857 38363 24915 38369
rect 24964 38372 27016 38400
rect 21468 38304 21772 38332
rect 21361 38295 21419 38301
rect 21637 38267 21695 38273
rect 21637 38264 21649 38267
rect 20180 38236 21649 38264
rect 21637 38233 21649 38236
rect 21683 38233 21695 38267
rect 21637 38227 21695 38233
rect 20622 38196 20628 38208
rect 19720 38168 20628 38196
rect 20622 38156 20628 38168
rect 20680 38156 20686 38208
rect 21744 38196 21772 38304
rect 22922 38292 22928 38344
rect 22980 38332 22986 38344
rect 23109 38335 23167 38341
rect 23109 38332 23121 38335
rect 22980 38304 23121 38332
rect 22980 38292 22986 38304
rect 23109 38301 23121 38304
rect 23155 38301 23167 38335
rect 23109 38295 23167 38301
rect 23293 38335 23351 38341
rect 23293 38301 23305 38335
rect 23339 38332 23351 38335
rect 23768 38332 23796 38363
rect 23339 38304 23796 38332
rect 24029 38335 24087 38341
rect 23339 38301 23351 38304
rect 23293 38295 23351 38301
rect 24029 38301 24041 38335
rect 24075 38332 24087 38335
rect 24302 38332 24308 38344
rect 24075 38304 24308 38332
rect 24075 38301 24087 38304
rect 24029 38295 24087 38301
rect 23308 38264 23336 38295
rect 24302 38292 24308 38304
rect 24360 38332 24366 38344
rect 24964 38332 24992 38372
rect 24360 38304 24992 38332
rect 25041 38335 25099 38341
rect 24360 38292 24366 38304
rect 25041 38301 25053 38335
rect 25087 38332 25099 38335
rect 25958 38332 25964 38344
rect 25087 38304 25964 38332
rect 25087 38301 25099 38304
rect 25041 38295 25099 38301
rect 25958 38292 25964 38304
rect 26016 38292 26022 38344
rect 22066 38236 23336 38264
rect 24581 38267 24639 38273
rect 22066 38196 22094 38236
rect 24581 38233 24593 38267
rect 24627 38264 24639 38267
rect 24627 38236 26924 38264
rect 24627 38233 24639 38236
rect 24581 38227 24639 38233
rect 21744 38168 22094 38196
rect 23753 38199 23811 38205
rect 23753 38165 23765 38199
rect 23799 38196 23811 38199
rect 25130 38196 25136 38208
rect 23799 38168 25136 38196
rect 23799 38165 23811 38168
rect 23753 38159 23811 38165
rect 25130 38156 25136 38168
rect 25188 38156 25194 38208
rect 25222 38156 25228 38208
rect 25280 38156 25286 38208
rect 26896 38205 26924 38236
rect 26881 38199 26939 38205
rect 26881 38165 26893 38199
rect 26927 38165 26939 38199
rect 26988 38196 27016 38372
rect 27249 38369 27261 38403
rect 27295 38400 27307 38403
rect 28534 38400 28540 38412
rect 27295 38372 28540 38400
rect 27295 38369 27307 38372
rect 27249 38363 27307 38369
rect 28534 38360 28540 38372
rect 28592 38360 28598 38412
rect 28902 38360 28908 38412
rect 28960 38400 28966 38412
rect 29733 38403 29791 38409
rect 29733 38400 29745 38403
rect 28960 38372 29745 38400
rect 28960 38360 28966 38372
rect 29733 38369 29745 38372
rect 29779 38369 29791 38403
rect 29733 38363 29791 38369
rect 30006 38360 30012 38412
rect 30064 38400 30070 38412
rect 32140 38400 32168 38508
rect 36832 38468 36860 38508
rect 36909 38505 36921 38539
rect 36955 38536 36967 38539
rect 37090 38536 37096 38548
rect 36955 38508 37096 38536
rect 36955 38505 36967 38508
rect 36909 38499 36967 38505
rect 37090 38496 37096 38508
rect 37148 38496 37154 38548
rect 38105 38539 38163 38545
rect 38105 38505 38117 38539
rect 38151 38536 38163 38539
rect 38654 38536 38660 38548
rect 38151 38508 38660 38536
rect 38151 38505 38163 38508
rect 38105 38499 38163 38505
rect 38654 38496 38660 38508
rect 38712 38496 38718 38548
rect 40681 38539 40739 38545
rect 40681 38505 40693 38539
rect 40727 38536 40739 38539
rect 43070 38536 43076 38548
rect 40727 38508 43076 38536
rect 40727 38505 40739 38508
rect 40681 38499 40739 38505
rect 43070 38496 43076 38508
rect 43128 38496 43134 38548
rect 39485 38471 39543 38477
rect 36832 38440 37872 38468
rect 30064 38372 32168 38400
rect 30064 38360 30070 38372
rect 36170 38360 36176 38412
rect 36228 38400 36234 38412
rect 36228 38372 36676 38400
rect 36228 38360 36234 38372
rect 27062 38292 27068 38344
rect 27120 38292 27126 38344
rect 27154 38292 27160 38344
rect 27212 38292 27218 38344
rect 27341 38335 27399 38341
rect 27341 38301 27353 38335
rect 27387 38332 27399 38335
rect 28166 38332 28172 38344
rect 27387 38304 28172 38332
rect 27387 38301 27399 38304
rect 27341 38295 27399 38301
rect 28166 38292 28172 38304
rect 28224 38332 28230 38344
rect 28442 38332 28448 38344
rect 28224 38304 28448 38332
rect 28224 38292 28230 38304
rect 28442 38292 28448 38304
rect 28500 38292 28506 38344
rect 30098 38292 30104 38344
rect 30156 38332 30162 38344
rect 30193 38335 30251 38341
rect 30193 38332 30205 38335
rect 30156 38304 30205 38332
rect 30156 38292 30162 38304
rect 30193 38301 30205 38304
rect 30239 38301 30251 38335
rect 30193 38295 30251 38301
rect 30466 38292 30472 38344
rect 30524 38292 30530 38344
rect 31386 38292 31392 38344
rect 31444 38332 31450 38344
rect 31481 38335 31539 38341
rect 31481 38332 31493 38335
rect 31444 38304 31493 38332
rect 31444 38292 31450 38304
rect 31481 38301 31493 38304
rect 31527 38332 31539 38335
rect 31570 38332 31576 38344
rect 31527 38304 31576 38332
rect 31527 38301 31539 38304
rect 31481 38295 31539 38301
rect 31570 38292 31576 38304
rect 31628 38292 31634 38344
rect 31754 38292 31760 38344
rect 31812 38292 31818 38344
rect 32674 38292 32680 38344
rect 32732 38292 32738 38344
rect 32766 38292 32772 38344
rect 32824 38292 32830 38344
rect 32861 38335 32919 38341
rect 32861 38301 32873 38335
rect 32907 38301 32919 38335
rect 32861 38295 32919 38301
rect 27522 38224 27528 38276
rect 27580 38264 27586 38276
rect 27985 38267 28043 38273
rect 27985 38264 27997 38267
rect 27580 38236 27997 38264
rect 27580 38224 27586 38236
rect 27985 38233 27997 38236
rect 28031 38233 28043 38267
rect 27985 38227 28043 38233
rect 28092 38236 28580 38264
rect 28092 38196 28120 38236
rect 26988 38168 28120 38196
rect 26881 38159 26939 38165
rect 28258 38156 28264 38208
rect 28316 38196 28322 38208
rect 28445 38199 28503 38205
rect 28445 38196 28457 38199
rect 28316 38168 28457 38196
rect 28316 38156 28322 38168
rect 28445 38165 28457 38168
rect 28491 38165 28503 38199
rect 28552 38196 28580 38236
rect 31662 38224 31668 38276
rect 31720 38224 31726 38276
rect 32876 38264 32904 38295
rect 33042 38292 33048 38344
rect 33100 38292 33106 38344
rect 34238 38292 34244 38344
rect 34296 38292 34302 38344
rect 34422 38292 34428 38344
rect 34480 38332 34486 38344
rect 34885 38335 34943 38341
rect 34885 38332 34897 38335
rect 34480 38304 34897 38332
rect 34480 38292 34486 38304
rect 34885 38301 34897 38304
rect 34931 38301 34943 38335
rect 34885 38295 34943 38301
rect 35066 38292 35072 38344
rect 35124 38292 35130 38344
rect 36078 38292 36084 38344
rect 36136 38332 36142 38344
rect 36265 38335 36323 38341
rect 36265 38332 36277 38335
rect 36136 38304 36277 38332
rect 36136 38292 36142 38304
rect 36265 38301 36277 38304
rect 36311 38301 36323 38335
rect 36265 38295 36323 38301
rect 36354 38292 36360 38344
rect 36412 38292 36418 38344
rect 36648 38341 36676 38372
rect 36633 38335 36691 38341
rect 36633 38301 36645 38335
rect 36679 38301 36691 38335
rect 36633 38295 36691 38301
rect 36722 38292 36728 38344
rect 36780 38341 36786 38344
rect 36780 38332 36788 38341
rect 36780 38304 36825 38332
rect 36780 38295 36788 38304
rect 36780 38292 36786 38295
rect 37458 38292 37464 38344
rect 37516 38292 37522 38344
rect 37642 38341 37648 38344
rect 37609 38335 37648 38341
rect 37609 38301 37621 38335
rect 37609 38295 37648 38301
rect 37642 38292 37648 38295
rect 37700 38292 37706 38344
rect 33594 38264 33600 38276
rect 32324 38236 32536 38264
rect 32876 38236 33600 38264
rect 32324 38196 32352 38236
rect 28552 38168 32352 38196
rect 28445 38159 28503 38165
rect 32398 38156 32404 38208
rect 32456 38156 32462 38208
rect 32508 38196 32536 38236
rect 33594 38224 33600 38236
rect 33652 38224 33658 38276
rect 33778 38224 33784 38276
rect 33836 38224 33842 38276
rect 34514 38224 34520 38276
rect 34572 38264 34578 38276
rect 36373 38264 36401 38292
rect 34572 38236 36401 38264
rect 36541 38267 36599 38273
rect 34572 38224 34578 38236
rect 36541 38233 36553 38267
rect 36587 38264 36599 38267
rect 36814 38264 36820 38276
rect 36587 38236 36820 38264
rect 36587 38233 36599 38236
rect 36541 38227 36599 38233
rect 32858 38196 32864 38208
rect 32508 38168 32864 38196
rect 32858 38156 32864 38168
rect 32916 38156 32922 38208
rect 34790 38156 34796 38208
rect 34848 38196 34854 38208
rect 34977 38199 35035 38205
rect 34977 38196 34989 38199
rect 34848 38168 34989 38196
rect 34848 38156 34854 38168
rect 34977 38165 34989 38168
rect 35023 38165 35035 38199
rect 34977 38159 35035 38165
rect 35986 38156 35992 38208
rect 36044 38196 36050 38208
rect 36556 38196 36584 38227
rect 36814 38224 36820 38236
rect 36872 38224 36878 38276
rect 36998 38224 37004 38276
rect 37056 38264 37062 38276
rect 37734 38264 37740 38276
rect 37056 38236 37740 38264
rect 37056 38224 37062 38236
rect 37734 38224 37740 38236
rect 37792 38224 37798 38276
rect 37844 38273 37872 38440
rect 39485 38437 39497 38471
rect 39531 38437 39543 38471
rect 39485 38431 39543 38437
rect 38764 38372 39436 38400
rect 37918 38292 37924 38344
rect 37976 38341 37982 38344
rect 37976 38332 37984 38341
rect 37976 38304 38021 38332
rect 37976 38295 37984 38304
rect 37976 38292 37982 38295
rect 37829 38267 37887 38273
rect 37829 38233 37841 38267
rect 37875 38264 37887 38267
rect 38654 38264 38660 38276
rect 37875 38236 38660 38264
rect 37875 38233 37887 38236
rect 37829 38227 37887 38233
rect 38654 38224 38660 38236
rect 38712 38224 38718 38276
rect 36044 38168 36584 38196
rect 36044 38156 36050 38168
rect 36906 38156 36912 38208
rect 36964 38196 36970 38208
rect 38764 38196 38792 38372
rect 38933 38335 38991 38341
rect 38933 38301 38945 38335
rect 38979 38332 38991 38335
rect 38979 38304 39068 38332
rect 38979 38301 38991 38304
rect 38933 38295 38991 38301
rect 36964 38168 38792 38196
rect 39040 38196 39068 38304
rect 39206 38292 39212 38344
rect 39264 38292 39270 38344
rect 39298 38292 39304 38344
rect 39356 38292 39362 38344
rect 39114 38224 39120 38276
rect 39172 38224 39178 38276
rect 39408 38264 39436 38372
rect 39500 38332 39528 38431
rect 40297 38372 41736 38400
rect 40037 38335 40095 38341
rect 40037 38332 40049 38335
rect 39500 38304 40049 38332
rect 40037 38301 40049 38304
rect 40083 38301 40095 38335
rect 40037 38295 40095 38301
rect 40130 38335 40188 38341
rect 40130 38301 40142 38335
rect 40176 38332 40188 38335
rect 40297 38332 40325 38372
rect 40176 38304 40325 38332
rect 40176 38301 40188 38304
rect 40130 38295 40188 38301
rect 40144 38264 40172 38295
rect 40402 38292 40408 38344
rect 40460 38292 40466 38344
rect 40543 38335 40601 38341
rect 40543 38301 40555 38335
rect 40589 38332 40601 38335
rect 41138 38332 41144 38344
rect 40589 38304 41144 38332
rect 40589 38301 40601 38304
rect 40543 38295 40601 38301
rect 41138 38292 41144 38304
rect 41196 38292 41202 38344
rect 39408 38236 40172 38264
rect 40313 38267 40371 38273
rect 40313 38233 40325 38267
rect 40359 38233 40371 38267
rect 41708 38264 41736 38372
rect 41782 38360 41788 38412
rect 41840 38360 41846 38412
rect 42052 38335 42110 38341
rect 42052 38301 42064 38335
rect 42098 38332 42110 38335
rect 42610 38332 42616 38344
rect 42098 38304 42616 38332
rect 42098 38301 42110 38304
rect 42052 38295 42110 38301
rect 42610 38292 42616 38304
rect 42668 38292 42674 38344
rect 42886 38264 42892 38276
rect 41708 38236 42892 38264
rect 40313 38227 40371 38233
rect 39206 38196 39212 38208
rect 39040 38168 39212 38196
rect 36964 38156 36970 38168
rect 39206 38156 39212 38168
rect 39264 38156 39270 38208
rect 40328 38196 40356 38227
rect 42886 38224 42892 38236
rect 42944 38224 42950 38276
rect 40402 38196 40408 38208
rect 40328 38168 40408 38196
rect 40402 38156 40408 38168
rect 40460 38156 40466 38208
rect 43070 38156 43076 38208
rect 43128 38196 43134 38208
rect 43165 38199 43223 38205
rect 43165 38196 43177 38199
rect 43128 38168 43177 38196
rect 43128 38156 43134 38168
rect 43165 38165 43177 38168
rect 43211 38165 43223 38199
rect 43165 38159 43223 38165
rect 1104 38106 43884 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 43884 38106
rect 1104 38032 43884 38054
rect 9582 37992 9588 38004
rect 7944 37964 9588 37992
rect 4614 37924 4620 37936
rect 4264 37896 4620 37924
rect 4264 37865 4292 37896
rect 4614 37884 4620 37896
rect 4672 37884 4678 37936
rect 7006 37884 7012 37936
rect 7064 37924 7070 37936
rect 7101 37927 7159 37933
rect 7101 37924 7113 37927
rect 7064 37896 7113 37924
rect 7064 37884 7070 37896
rect 7101 37893 7113 37896
rect 7147 37893 7159 37927
rect 7101 37887 7159 37893
rect 4249 37859 4307 37865
rect 4249 37825 4261 37859
rect 4295 37825 4307 37859
rect 4249 37819 4307 37825
rect 4516 37859 4574 37865
rect 4516 37825 4528 37859
rect 4562 37856 4574 37859
rect 4890 37856 4896 37868
rect 4562 37828 4896 37856
rect 4562 37825 4574 37828
rect 4516 37819 4574 37825
rect 4890 37816 4896 37828
rect 4948 37816 4954 37868
rect 7190 37816 7196 37868
rect 7248 37856 7254 37868
rect 7285 37859 7343 37865
rect 7285 37856 7297 37859
rect 7248 37828 7297 37856
rect 7248 37816 7254 37828
rect 7285 37825 7297 37828
rect 7331 37856 7343 37859
rect 7834 37856 7840 37868
rect 7331 37828 7840 37856
rect 7331 37825 7343 37828
rect 7285 37819 7343 37825
rect 7834 37816 7840 37828
rect 7892 37816 7898 37868
rect 7944 37865 7972 37964
rect 9582 37952 9588 37964
rect 9640 37952 9646 38004
rect 12618 37952 12624 38004
rect 12676 37992 12682 38004
rect 13998 37992 14004 38004
rect 12676 37964 14004 37992
rect 12676 37952 12682 37964
rect 13998 37952 14004 37964
rect 14056 37952 14062 38004
rect 18233 37995 18291 38001
rect 18233 37961 18245 37995
rect 18279 37992 18291 37995
rect 18690 37992 18696 38004
rect 18279 37964 18696 37992
rect 18279 37961 18291 37964
rect 18233 37955 18291 37961
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 19334 37952 19340 38004
rect 19392 37992 19398 38004
rect 23474 37992 23480 38004
rect 19392 37964 23480 37992
rect 19392 37952 19398 37964
rect 23474 37952 23480 37964
rect 23532 37952 23538 38004
rect 23569 37995 23627 38001
rect 23569 37961 23581 37995
rect 23615 37992 23627 37995
rect 24854 37992 24860 38004
rect 23615 37964 24860 37992
rect 23615 37961 23627 37964
rect 23569 37955 23627 37961
rect 24854 37952 24860 37964
rect 24912 37952 24918 38004
rect 25041 37995 25099 38001
rect 25041 37961 25053 37995
rect 25087 37961 25099 37995
rect 25041 37955 25099 37961
rect 9858 37924 9864 37936
rect 8220 37896 9864 37924
rect 7929 37859 7987 37865
rect 7929 37825 7941 37859
rect 7975 37825 7987 37859
rect 7929 37819 7987 37825
rect 8110 37816 8116 37868
rect 8168 37816 8174 37868
rect 8220 37865 8248 37896
rect 9858 37884 9864 37896
rect 9916 37884 9922 37936
rect 10226 37884 10232 37936
rect 10284 37924 10290 37936
rect 14553 37927 14611 37933
rect 10284 37896 14412 37924
rect 10284 37884 10290 37896
rect 8205 37859 8263 37865
rect 8205 37825 8217 37859
rect 8251 37825 8263 37859
rect 8205 37819 8263 37825
rect 9030 37816 9036 37868
rect 9088 37816 9094 37868
rect 10045 37859 10103 37865
rect 10045 37825 10057 37859
rect 10091 37856 10103 37859
rect 10410 37856 10416 37868
rect 10091 37828 10416 37856
rect 10091 37825 10103 37828
rect 10045 37819 10103 37825
rect 10410 37816 10416 37828
rect 10468 37816 10474 37868
rect 10502 37816 10508 37868
rect 10560 37856 10566 37868
rect 10965 37859 11023 37865
rect 10560 37828 10824 37856
rect 10560 37816 10566 37828
rect 7469 37791 7527 37797
rect 7469 37757 7481 37791
rect 7515 37788 7527 37791
rect 9490 37788 9496 37800
rect 7515 37760 9496 37788
rect 7515 37757 7527 37760
rect 7469 37751 7527 37757
rect 9490 37748 9496 37760
rect 9548 37788 9554 37800
rect 9548 37760 10640 37788
rect 9548 37748 9554 37760
rect 8389 37723 8447 37729
rect 8389 37689 8401 37723
rect 8435 37720 8447 37723
rect 9674 37720 9680 37732
rect 8435 37692 9680 37720
rect 8435 37689 8447 37692
rect 8389 37683 8447 37689
rect 9674 37680 9680 37692
rect 9732 37680 9738 37732
rect 10502 37720 10508 37732
rect 9784 37692 10508 37720
rect 5534 37612 5540 37664
rect 5592 37652 5598 37664
rect 5629 37655 5687 37661
rect 5629 37652 5641 37655
rect 5592 37624 5641 37652
rect 5592 37612 5598 37624
rect 5629 37621 5641 37624
rect 5675 37621 5687 37655
rect 5629 37615 5687 37621
rect 7374 37612 7380 37664
rect 7432 37652 7438 37664
rect 8205 37655 8263 37661
rect 8205 37652 8217 37655
rect 7432 37624 8217 37652
rect 7432 37612 7438 37624
rect 8205 37621 8217 37624
rect 8251 37652 8263 37655
rect 9784 37652 9812 37692
rect 10502 37680 10508 37692
rect 10560 37680 10566 37732
rect 10612 37720 10640 37760
rect 10686 37748 10692 37800
rect 10744 37748 10750 37800
rect 10796 37797 10824 37828
rect 10965 37825 10977 37859
rect 11011 37856 11023 37859
rect 11054 37856 11060 37868
rect 11011 37828 11060 37856
rect 11011 37825 11023 37828
rect 10965 37819 11023 37825
rect 11054 37816 11060 37828
rect 11112 37816 11118 37868
rect 11885 37859 11943 37865
rect 11885 37856 11897 37859
rect 11532 37828 11897 37856
rect 10781 37791 10839 37797
rect 10781 37757 10793 37791
rect 10827 37788 10839 37791
rect 11422 37788 11428 37800
rect 10827 37760 11428 37788
rect 10827 37757 10839 37760
rect 10781 37751 10839 37757
rect 11422 37748 11428 37760
rect 11480 37748 11486 37800
rect 11532 37720 11560 37828
rect 11885 37825 11897 37828
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 11977 37859 12035 37865
rect 11977 37825 11989 37859
rect 12023 37825 12035 37859
rect 11977 37819 12035 37825
rect 12161 37859 12219 37865
rect 12161 37825 12173 37859
rect 12207 37825 12219 37859
rect 12161 37819 12219 37825
rect 12253 37859 12311 37865
rect 12253 37825 12265 37859
rect 12299 37856 12311 37859
rect 12342 37856 12348 37868
rect 12299 37828 12348 37856
rect 12299 37825 12311 37828
rect 12253 37819 12311 37825
rect 10612 37692 11560 37720
rect 8251 37624 9812 37652
rect 8251 37621 8263 37624
rect 8205 37615 8263 37621
rect 9858 37612 9864 37664
rect 9916 37652 9922 37664
rect 9953 37655 10011 37661
rect 9953 37652 9965 37655
rect 9916 37624 9965 37652
rect 9916 37612 9922 37624
rect 9953 37621 9965 37624
rect 9999 37652 10011 37655
rect 10686 37652 10692 37664
rect 9999 37624 10692 37652
rect 9999 37621 10011 37624
rect 9953 37615 10011 37621
rect 10686 37612 10692 37624
rect 10744 37612 10750 37664
rect 11149 37655 11207 37661
rect 11149 37621 11161 37655
rect 11195 37652 11207 37655
rect 11514 37652 11520 37664
rect 11195 37624 11520 37652
rect 11195 37621 11207 37624
rect 11149 37615 11207 37621
rect 11514 37612 11520 37624
rect 11572 37612 11578 37664
rect 11606 37612 11612 37664
rect 11664 37652 11670 37664
rect 11701 37655 11759 37661
rect 11701 37652 11713 37655
rect 11664 37624 11713 37652
rect 11664 37612 11670 37624
rect 11701 37621 11713 37624
rect 11747 37621 11759 37655
rect 11992 37652 12020 37819
rect 12176 37720 12204 37819
rect 12342 37816 12348 37828
rect 12400 37816 12406 37868
rect 12713 37859 12771 37865
rect 12713 37825 12725 37859
rect 12759 37856 12771 37859
rect 12802 37856 12808 37868
rect 12759 37828 12808 37856
rect 12759 37825 12771 37828
rect 12713 37819 12771 37825
rect 12802 37816 12808 37828
rect 12860 37816 12866 37868
rect 12897 37859 12955 37865
rect 12897 37825 12909 37859
rect 12943 37856 12955 37859
rect 13078 37856 13084 37868
rect 12943 37828 13084 37856
rect 12943 37825 12955 37828
rect 12897 37819 12955 37825
rect 13078 37816 13084 37828
rect 13136 37816 13142 37868
rect 13814 37816 13820 37868
rect 13872 37816 13878 37868
rect 13998 37816 14004 37868
rect 14056 37816 14062 37868
rect 14090 37816 14096 37868
rect 14148 37816 14154 37868
rect 14384 37865 14412 37896
rect 14553 37893 14565 37927
rect 14599 37924 14611 37927
rect 16117 37927 16175 37933
rect 16117 37924 16129 37927
rect 14599 37896 16129 37924
rect 14599 37893 14611 37896
rect 14553 37887 14611 37893
rect 16117 37893 16129 37896
rect 16163 37893 16175 37927
rect 16117 37887 16175 37893
rect 16666 37884 16672 37936
rect 16724 37924 16730 37936
rect 16724 37896 19196 37924
rect 16724 37884 16730 37896
rect 14369 37859 14427 37865
rect 14369 37825 14381 37859
rect 14415 37856 14427 37859
rect 14826 37856 14832 37868
rect 14415 37828 14832 37856
rect 14415 37825 14427 37828
rect 14369 37819 14427 37825
rect 14826 37816 14832 37828
rect 14884 37816 14890 37868
rect 15930 37816 15936 37868
rect 15988 37816 15994 37868
rect 16025 37859 16083 37865
rect 16025 37825 16037 37859
rect 16071 37856 16083 37859
rect 16574 37856 16580 37868
rect 16071 37828 16580 37856
rect 16071 37825 16083 37828
rect 16025 37819 16083 37825
rect 16574 37816 16580 37828
rect 16632 37816 16638 37868
rect 16853 37859 16911 37865
rect 16853 37825 16865 37859
rect 16899 37825 16911 37859
rect 16853 37819 16911 37825
rect 14182 37748 14188 37800
rect 14240 37788 14246 37800
rect 14240 37760 15884 37788
rect 14240 37748 14246 37760
rect 12710 37720 12716 37732
rect 12176 37692 12716 37720
rect 12710 37680 12716 37692
rect 12768 37720 12774 37732
rect 13081 37723 13139 37729
rect 13081 37720 13093 37723
rect 12768 37692 13093 37720
rect 12768 37680 12774 37692
rect 13081 37689 13093 37692
rect 13127 37720 13139 37723
rect 15102 37720 15108 37732
rect 13127 37692 15108 37720
rect 13127 37689 13139 37692
rect 13081 37683 13139 37689
rect 15102 37680 15108 37692
rect 15160 37680 15166 37732
rect 15746 37680 15752 37732
rect 15804 37680 15810 37732
rect 15856 37720 15884 37760
rect 16482 37748 16488 37800
rect 16540 37788 16546 37800
rect 16868 37788 16896 37819
rect 16942 37816 16948 37868
rect 17000 37856 17006 37868
rect 17037 37859 17095 37865
rect 17037 37856 17049 37859
rect 17000 37828 17049 37856
rect 17000 37816 17006 37828
rect 17037 37825 17049 37828
rect 17083 37825 17095 37859
rect 17037 37819 17095 37825
rect 17773 37859 17831 37865
rect 17773 37825 17785 37859
rect 17819 37825 17831 37859
rect 17773 37819 17831 37825
rect 16540 37760 16896 37788
rect 17788 37788 17816 37819
rect 17954 37816 17960 37868
rect 18012 37816 18018 37868
rect 18046 37816 18052 37868
rect 18104 37816 18110 37868
rect 19168 37856 19196 37896
rect 19426 37884 19432 37936
rect 19484 37924 19490 37936
rect 19705 37927 19763 37933
rect 19705 37924 19717 37927
rect 19484 37896 19717 37924
rect 19484 37884 19490 37896
rect 19705 37893 19717 37896
rect 19751 37893 19763 37927
rect 19705 37887 19763 37893
rect 20254 37884 20260 37936
rect 20312 37924 20318 37936
rect 25056 37924 25084 37955
rect 25406 37952 25412 38004
rect 25464 37992 25470 38004
rect 29733 37995 29791 38001
rect 25464 37964 29500 37992
rect 25464 37952 25470 37964
rect 20312 37896 25084 37924
rect 20312 37884 20318 37896
rect 25222 37884 25228 37936
rect 25280 37924 25286 37936
rect 29472 37924 29500 37964
rect 29733 37961 29745 37995
rect 29779 37992 29791 37995
rect 30374 37992 30380 38004
rect 29779 37964 30380 37992
rect 29779 37961 29791 37964
rect 29733 37955 29791 37961
rect 30374 37952 30380 37964
rect 30432 37952 30438 38004
rect 33594 37952 33600 38004
rect 33652 37992 33658 38004
rect 34330 37992 34336 38004
rect 33652 37964 34336 37992
rect 33652 37952 33658 37964
rect 34330 37952 34336 37964
rect 34388 37992 34394 38004
rect 34609 37995 34667 38001
rect 34609 37992 34621 37995
rect 34388 37964 34621 37992
rect 34388 37952 34394 37964
rect 34609 37961 34621 37964
rect 34655 37961 34667 37995
rect 34609 37955 34667 37961
rect 36078 37952 36084 38004
rect 36136 37952 36142 38004
rect 36170 37952 36176 38004
rect 36228 37952 36234 38004
rect 36262 37952 36268 38004
rect 36320 37992 36326 38004
rect 36449 37995 36507 38001
rect 36449 37992 36461 37995
rect 36320 37964 36461 37992
rect 36320 37952 36326 37964
rect 36449 37961 36461 37964
rect 36495 37961 36507 37995
rect 41233 37995 41291 38001
rect 36449 37955 36507 37961
rect 40696 37964 41092 37992
rect 25280 37896 29408 37924
rect 29472 37896 31616 37924
rect 25280 37884 25286 37896
rect 19168 37828 19840 37856
rect 19812 37788 19840 37828
rect 19886 37816 19892 37868
rect 19944 37816 19950 37868
rect 19988 37859 20046 37865
rect 19988 37825 20000 37859
rect 20034 37856 20046 37859
rect 20162 37856 20168 37868
rect 20034 37828 20168 37856
rect 20034 37825 20046 37828
rect 19988 37819 20046 37825
rect 20162 37816 20168 37828
rect 20220 37856 20226 37868
rect 20714 37856 20720 37868
rect 20220 37828 20720 37856
rect 20220 37816 20226 37828
rect 20714 37816 20720 37828
rect 20772 37816 20778 37868
rect 22189 37859 22247 37865
rect 22189 37825 22201 37859
rect 22235 37825 22247 37859
rect 22189 37819 22247 37825
rect 20073 37791 20131 37797
rect 20073 37788 20085 37791
rect 17788 37760 19748 37788
rect 19812 37760 20085 37788
rect 16540 37748 16546 37760
rect 17865 37723 17923 37729
rect 17865 37720 17877 37723
rect 15856 37692 17877 37720
rect 17865 37689 17877 37692
rect 17911 37689 17923 37723
rect 19720 37720 19748 37760
rect 20073 37757 20085 37760
rect 20119 37788 20131 37791
rect 21082 37788 21088 37800
rect 20119 37760 21088 37788
rect 20119 37757 20131 37760
rect 20073 37751 20131 37757
rect 21082 37748 21088 37760
rect 21140 37748 21146 37800
rect 22204 37732 22232 37819
rect 22554 37816 22560 37868
rect 22612 37816 22618 37868
rect 22738 37816 22744 37868
rect 22796 37816 22802 37868
rect 23382 37816 23388 37868
rect 23440 37816 23446 37868
rect 23474 37816 23480 37868
rect 23532 37856 23538 37868
rect 24397 37859 24455 37865
rect 24397 37856 24409 37859
rect 23532 37828 24409 37856
rect 23532 37816 23538 37828
rect 24397 37825 24409 37828
rect 24443 37856 24455 37859
rect 24486 37856 24492 37868
rect 24443 37828 24492 37856
rect 24443 37825 24455 37828
rect 24397 37819 24455 37825
rect 24486 37816 24492 37828
rect 24544 37816 24550 37868
rect 24857 37859 24915 37865
rect 24857 37825 24869 37859
rect 24903 37825 24915 37859
rect 24857 37819 24915 37825
rect 22370 37748 22376 37800
rect 22428 37748 22434 37800
rect 22462 37748 22468 37800
rect 22520 37748 22526 37800
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37757 23259 37791
rect 23201 37751 23259 37757
rect 19720 37692 22140 37720
rect 17865 37683 17923 37689
rect 12250 37652 12256 37664
rect 11992 37624 12256 37652
rect 11701 37615 11759 37621
rect 12250 37612 12256 37624
rect 12308 37652 12314 37664
rect 12986 37652 12992 37664
rect 12308 37624 12992 37652
rect 12308 37612 12314 37624
rect 12986 37612 12992 37624
rect 13044 37652 13050 37664
rect 14366 37652 14372 37664
rect 13044 37624 14372 37652
rect 13044 37612 13050 37624
rect 14366 37612 14372 37624
rect 14424 37612 14430 37664
rect 16298 37612 16304 37664
rect 16356 37612 16362 37664
rect 16758 37612 16764 37664
rect 16816 37652 16822 37664
rect 17221 37655 17279 37661
rect 17221 37652 17233 37655
rect 16816 37624 17233 37652
rect 16816 37612 16822 37624
rect 17221 37621 17233 37624
rect 17267 37621 17279 37655
rect 17221 37615 17279 37621
rect 21266 37612 21272 37664
rect 21324 37652 21330 37664
rect 22005 37655 22063 37661
rect 22005 37652 22017 37655
rect 21324 37624 22017 37652
rect 21324 37612 21330 37624
rect 22005 37621 22017 37624
rect 22051 37621 22063 37655
rect 22112 37652 22140 37692
rect 22186 37680 22192 37732
rect 22244 37720 22250 37732
rect 23216 37720 23244 37751
rect 24762 37748 24768 37800
rect 24820 37748 24826 37800
rect 22244 37692 23244 37720
rect 24872 37720 24900 37819
rect 25130 37816 25136 37868
rect 25188 37856 25194 37868
rect 25188 37828 25728 37856
rect 25188 37816 25194 37828
rect 25700 37788 25728 37828
rect 25866 37816 25872 37868
rect 25924 37816 25930 37868
rect 26145 37859 26203 37865
rect 26145 37825 26157 37859
rect 26191 37856 26203 37859
rect 26694 37856 26700 37868
rect 26191 37828 26700 37856
rect 26191 37825 26203 37828
rect 26145 37819 26203 37825
rect 26694 37816 26700 37828
rect 26752 37816 26758 37868
rect 27062 37816 27068 37868
rect 27120 37856 27126 37868
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 27120 37828 27169 37856
rect 27120 37816 27126 37828
rect 27157 37825 27169 37828
rect 27203 37825 27215 37859
rect 27157 37819 27215 37825
rect 27341 37859 27399 37865
rect 27341 37825 27353 37859
rect 27387 37856 27399 37859
rect 27522 37856 27528 37868
rect 27387 37828 27528 37856
rect 27387 37825 27399 37828
rect 27341 37819 27399 37825
rect 27522 37816 27528 37828
rect 27580 37856 27586 37868
rect 28074 37856 28080 37868
rect 27580 37828 28080 37856
rect 27580 37816 27586 37828
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 28626 37816 28632 37868
rect 28684 37856 28690 37868
rect 29380 37865 29408 37896
rect 28721 37859 28779 37865
rect 28721 37856 28733 37859
rect 28684 37828 28733 37856
rect 28684 37816 28690 37828
rect 28721 37825 28733 37828
rect 28767 37825 28779 37859
rect 28721 37819 28779 37825
rect 28905 37859 28963 37865
rect 28905 37825 28917 37859
rect 28951 37825 28963 37859
rect 28905 37819 28963 37825
rect 29365 37859 29423 37865
rect 29365 37825 29377 37859
rect 29411 37825 29423 37859
rect 29365 37819 29423 37825
rect 25774 37788 25780 37800
rect 25700 37760 25780 37788
rect 25774 37748 25780 37760
rect 25832 37788 25838 37800
rect 25961 37791 26019 37797
rect 25961 37788 25973 37791
rect 25832 37760 25973 37788
rect 25832 37748 25838 37760
rect 25961 37757 25973 37760
rect 26007 37757 26019 37791
rect 25961 37751 26019 37757
rect 26234 37748 26240 37800
rect 26292 37788 26298 37800
rect 27080 37788 27108 37816
rect 26292 37760 27108 37788
rect 26292 37748 26298 37760
rect 25866 37720 25872 37732
rect 24872 37692 25872 37720
rect 22244 37680 22250 37692
rect 25866 37680 25872 37692
rect 25924 37680 25930 37732
rect 28920 37720 28948 37819
rect 30190 37816 30196 37868
rect 30248 37816 30254 37868
rect 30374 37816 30380 37868
rect 30432 37816 30438 37868
rect 31588 37865 31616 37896
rect 31662 37884 31668 37936
rect 31720 37924 31726 37936
rect 34057 37927 34115 37933
rect 34057 37924 34069 37927
rect 31720 37896 32536 37924
rect 31720 37884 31726 37896
rect 31573 37859 31631 37865
rect 31573 37825 31585 37859
rect 31619 37825 31631 37859
rect 31573 37819 31631 37825
rect 32306 37816 32312 37868
rect 32364 37816 32370 37868
rect 32508 37865 32536 37896
rect 33612 37896 34069 37924
rect 32493 37859 32551 37865
rect 32493 37825 32505 37859
rect 32539 37825 32551 37859
rect 32493 37819 32551 37825
rect 33612 37800 33640 37896
rect 34057 37893 34069 37896
rect 34103 37924 34115 37927
rect 34422 37924 34428 37936
rect 34103 37896 34428 37924
rect 34103 37893 34115 37896
rect 34057 37887 34115 37893
rect 34422 37884 34428 37896
rect 34480 37924 34486 37936
rect 34977 37927 35035 37933
rect 34977 37924 34989 37927
rect 34480 37896 34989 37924
rect 34480 37884 34486 37896
rect 34977 37893 34989 37896
rect 35023 37893 35035 37927
rect 36096 37924 36124 37952
rect 34977 37887 35035 37893
rect 35820 37896 36124 37924
rect 36188 37924 36216 37952
rect 40696 37924 40724 37964
rect 36188 37896 38884 37924
rect 33778 37816 33784 37868
rect 33836 37816 33842 37868
rect 33873 37859 33931 37865
rect 33873 37825 33885 37859
rect 33919 37856 33931 37859
rect 33962 37856 33968 37868
rect 33919 37828 33968 37856
rect 33919 37825 33931 37828
rect 33873 37819 33931 37825
rect 33962 37816 33968 37828
rect 34020 37816 34026 37868
rect 34793 37859 34851 37865
rect 34793 37825 34805 37859
rect 34839 37856 34851 37859
rect 35066 37856 35072 37868
rect 34839 37828 35072 37856
rect 34839 37825 34851 37828
rect 34793 37819 34851 37825
rect 29454 37748 29460 37800
rect 29512 37748 29518 37800
rect 30006 37748 30012 37800
rect 30064 37788 30070 37800
rect 31297 37791 31355 37797
rect 31297 37788 31309 37791
rect 30064 37760 31309 37788
rect 30064 37748 30070 37760
rect 31297 37757 31309 37760
rect 31343 37757 31355 37791
rect 33594 37788 33600 37800
rect 31297 37751 31355 37757
rect 31404 37760 33600 37788
rect 31404 37720 31432 37760
rect 33594 37748 33600 37760
rect 33652 37748 33658 37800
rect 28920 37692 31432 37720
rect 31757 37723 31815 37729
rect 31757 37689 31769 37723
rect 31803 37720 31815 37723
rect 34422 37720 34428 37732
rect 31803 37692 34428 37720
rect 31803 37689 31815 37692
rect 31757 37683 31815 37689
rect 34422 37680 34428 37692
rect 34480 37680 34486 37732
rect 24486 37652 24492 37664
rect 22112 37624 24492 37652
rect 22005 37615 22063 37621
rect 24486 37612 24492 37624
rect 24544 37612 24550 37664
rect 24765 37655 24823 37661
rect 24765 37621 24777 37655
rect 24811 37652 24823 37655
rect 25222 37652 25228 37664
rect 24811 37624 25228 37652
rect 24811 37621 24823 37624
rect 24765 37615 24823 37621
rect 25222 37612 25228 37624
rect 25280 37612 25286 37664
rect 25682 37612 25688 37664
rect 25740 37612 25746 37664
rect 26142 37612 26148 37664
rect 26200 37612 26206 37664
rect 27157 37655 27215 37661
rect 27157 37621 27169 37655
rect 27203 37652 27215 37655
rect 27706 37652 27712 37664
rect 27203 37624 27712 37652
rect 27203 37621 27215 37624
rect 27157 37615 27215 37621
rect 27706 37612 27712 37624
rect 27764 37652 27770 37664
rect 28626 37652 28632 37664
rect 27764 37624 28632 37652
rect 27764 37612 27770 37624
rect 28626 37612 28632 37624
rect 28684 37612 28690 37664
rect 28718 37612 28724 37664
rect 28776 37612 28782 37664
rect 29546 37612 29552 37664
rect 29604 37612 29610 37664
rect 30193 37655 30251 37661
rect 30193 37621 30205 37655
rect 30239 37652 30251 37655
rect 30282 37652 30288 37664
rect 30239 37624 30288 37652
rect 30239 37621 30251 37624
rect 30193 37615 30251 37621
rect 30282 37612 30288 37624
rect 30340 37612 30346 37664
rect 31389 37655 31447 37661
rect 31389 37621 31401 37655
rect 31435 37652 31447 37655
rect 32030 37652 32036 37664
rect 31435 37624 32036 37652
rect 31435 37621 31447 37624
rect 31389 37615 31447 37621
rect 32030 37612 32036 37624
rect 32088 37612 32094 37664
rect 32398 37612 32404 37664
rect 32456 37652 32462 37664
rect 32585 37655 32643 37661
rect 32585 37652 32597 37655
rect 32456 37624 32597 37652
rect 32456 37612 32462 37624
rect 32585 37621 32597 37624
rect 32631 37652 32643 37655
rect 34808 37652 34836 37819
rect 35066 37816 35072 37828
rect 35124 37816 35130 37868
rect 35820 37865 35848 37896
rect 35805 37859 35863 37865
rect 35805 37825 35817 37859
rect 35851 37825 35863 37859
rect 35805 37819 35863 37825
rect 35894 37816 35900 37868
rect 35952 37856 35958 37868
rect 36081 37859 36139 37865
rect 35952 37828 35997 37856
rect 35952 37816 35958 37828
rect 36081 37825 36093 37859
rect 36127 37825 36139 37859
rect 36081 37819 36139 37825
rect 36173 37859 36231 37865
rect 36173 37825 36185 37859
rect 36219 37825 36231 37859
rect 36173 37819 36231 37825
rect 36311 37859 36369 37865
rect 36311 37825 36323 37859
rect 36357 37856 36369 37859
rect 36446 37856 36452 37868
rect 36357 37828 36452 37856
rect 36357 37825 36369 37828
rect 36311 37819 36369 37825
rect 35986 37748 35992 37800
rect 36044 37788 36050 37800
rect 36096 37788 36124 37819
rect 36044 37760 36124 37788
rect 36188 37788 36216 37819
rect 36446 37816 36452 37828
rect 36504 37856 36510 37868
rect 36722 37856 36728 37868
rect 36504 37828 36728 37856
rect 36504 37816 36510 37828
rect 36722 37816 36728 37828
rect 36780 37816 36786 37868
rect 37274 37816 37280 37868
rect 37332 37856 37338 37868
rect 38856 37865 38884 37896
rect 38948 37896 40724 37924
rect 37553 37859 37611 37865
rect 37553 37856 37565 37859
rect 37332 37828 37565 37856
rect 37332 37816 37338 37828
rect 37553 37825 37565 37828
rect 37599 37825 37611 37859
rect 37553 37819 37611 37825
rect 38841 37859 38899 37865
rect 38841 37825 38853 37859
rect 38887 37825 38899 37859
rect 38841 37819 38899 37825
rect 38105 37791 38163 37797
rect 36188 37760 36308 37788
rect 36044 37748 36050 37760
rect 32631 37624 34836 37652
rect 36280 37652 36308 37760
rect 38105 37757 38117 37791
rect 38151 37788 38163 37791
rect 38286 37788 38292 37800
rect 38151 37760 38292 37788
rect 38151 37757 38163 37760
rect 38105 37751 38163 37757
rect 38286 37748 38292 37760
rect 38344 37748 38350 37800
rect 36354 37680 36360 37732
rect 36412 37720 36418 37732
rect 38948 37720 38976 37896
rect 39025 37859 39083 37865
rect 39025 37825 39037 37859
rect 39071 37825 39083 37859
rect 39025 37819 39083 37825
rect 39117 37859 39175 37865
rect 39117 37825 39129 37859
rect 39163 37825 39175 37859
rect 39117 37819 39175 37825
rect 39209 37859 39267 37865
rect 39209 37825 39221 37859
rect 39255 37856 39267 37859
rect 39298 37856 39304 37868
rect 39255 37828 39304 37856
rect 39255 37825 39267 37828
rect 39209 37819 39267 37825
rect 36412 37692 38976 37720
rect 39040 37720 39068 37819
rect 39132 37788 39160 37819
rect 39298 37816 39304 37828
rect 39356 37816 39362 37868
rect 40696 37865 40724 37896
rect 40954 37884 40960 37936
rect 41012 37884 41018 37936
rect 41064 37924 41092 37964
rect 41233 37961 41245 37995
rect 41279 37992 41291 37995
rect 42702 37992 42708 38004
rect 41279 37964 42708 37992
rect 41279 37961 41291 37964
rect 41233 37955 41291 37961
rect 42702 37952 42708 37964
rect 42760 37952 42766 38004
rect 43070 37924 43076 37936
rect 41064 37896 43076 37924
rect 43070 37884 43076 37896
rect 43128 37884 43134 37936
rect 41138 37865 41144 37868
rect 40589 37859 40647 37865
rect 40589 37856 40601 37859
rect 39408 37828 40601 37856
rect 39132 37760 39344 37788
rect 39114 37720 39120 37732
rect 39040 37692 39120 37720
rect 36412 37680 36418 37692
rect 39114 37680 39120 37692
rect 39172 37680 39178 37732
rect 39206 37652 39212 37664
rect 36280 37624 39212 37652
rect 32631 37621 32643 37624
rect 32585 37615 32643 37621
rect 39206 37612 39212 37624
rect 39264 37612 39270 37664
rect 39316 37652 39344 37760
rect 39408 37729 39436 37828
rect 40589 37825 40601 37828
rect 40635 37825 40647 37859
rect 40589 37819 40647 37825
rect 40682 37859 40740 37865
rect 40682 37825 40694 37859
rect 40728 37825 40740 37859
rect 40682 37819 40740 37825
rect 40865 37859 40923 37865
rect 40865 37825 40877 37859
rect 40911 37825 40923 37859
rect 40865 37819 40923 37825
rect 41095 37859 41144 37865
rect 41095 37825 41107 37859
rect 41141 37825 41144 37859
rect 41095 37819 41144 37825
rect 40402 37748 40408 37800
rect 40460 37788 40466 37800
rect 40880 37788 40908 37819
rect 41138 37816 41144 37819
rect 41196 37816 41202 37868
rect 42889 37859 42947 37865
rect 42889 37825 42901 37859
rect 42935 37856 42947 37859
rect 42978 37856 42984 37868
rect 42935 37828 42984 37856
rect 42935 37825 42947 37828
rect 42889 37819 42947 37825
rect 42978 37816 42984 37828
rect 43036 37816 43042 37868
rect 40460 37760 40908 37788
rect 43165 37791 43223 37797
rect 40460 37748 40466 37760
rect 43165 37757 43177 37791
rect 43211 37788 43223 37791
rect 43990 37788 43996 37800
rect 43211 37760 43996 37788
rect 43211 37757 43223 37760
rect 43165 37751 43223 37757
rect 43990 37748 43996 37760
rect 44048 37748 44054 37800
rect 39393 37723 39451 37729
rect 39393 37689 39405 37723
rect 39439 37689 39451 37723
rect 39393 37683 39451 37689
rect 39666 37652 39672 37664
rect 39316 37624 39672 37652
rect 39666 37612 39672 37624
rect 39724 37612 39730 37664
rect 1104 37562 43884 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 43884 37562
rect 1104 37488 43884 37510
rect 4890 37408 4896 37460
rect 4948 37408 4954 37460
rect 11698 37448 11704 37460
rect 11164 37420 11704 37448
rect 11164 37392 11192 37420
rect 11698 37408 11704 37420
rect 11756 37408 11762 37460
rect 11974 37408 11980 37460
rect 12032 37448 12038 37460
rect 12437 37451 12495 37457
rect 12437 37448 12449 37451
rect 12032 37420 12449 37448
rect 12032 37408 12038 37420
rect 12437 37417 12449 37420
rect 12483 37417 12495 37451
rect 12437 37411 12495 37417
rect 12529 37451 12587 37457
rect 12529 37417 12541 37451
rect 12575 37448 12587 37451
rect 13262 37448 13268 37460
rect 12575 37420 13268 37448
rect 12575 37417 12587 37420
rect 12529 37411 12587 37417
rect 13262 37408 13268 37420
rect 13320 37408 13326 37460
rect 14090 37408 14096 37460
rect 14148 37448 14154 37460
rect 14553 37451 14611 37457
rect 14553 37448 14565 37451
rect 14148 37420 14565 37448
rect 14148 37408 14154 37420
rect 14553 37417 14565 37420
rect 14599 37448 14611 37451
rect 14734 37448 14740 37460
rect 14599 37420 14740 37448
rect 14599 37417 14611 37420
rect 14553 37411 14611 37417
rect 14734 37408 14740 37420
rect 14792 37408 14798 37460
rect 20438 37408 20444 37460
rect 20496 37408 20502 37460
rect 22370 37408 22376 37460
rect 22428 37448 22434 37460
rect 22557 37451 22615 37457
rect 22557 37448 22569 37451
rect 22428 37420 22569 37448
rect 22428 37408 22434 37420
rect 22557 37417 22569 37420
rect 22603 37417 22615 37451
rect 22557 37411 22615 37417
rect 25133 37451 25191 37457
rect 25133 37417 25145 37451
rect 25179 37448 25191 37451
rect 26050 37448 26056 37460
rect 25179 37420 26056 37448
rect 25179 37417 25191 37420
rect 25133 37411 25191 37417
rect 26050 37408 26056 37420
rect 26108 37408 26114 37460
rect 26881 37451 26939 37457
rect 26881 37417 26893 37451
rect 26927 37448 26939 37451
rect 27614 37448 27620 37460
rect 26927 37420 27620 37448
rect 26927 37417 26939 37420
rect 26881 37411 26939 37417
rect 27614 37408 27620 37420
rect 27672 37408 27678 37460
rect 36446 37448 36452 37460
rect 32784 37420 36452 37448
rect 9861 37383 9919 37389
rect 9861 37349 9873 37383
rect 9907 37380 9919 37383
rect 11146 37380 11152 37392
rect 9907 37352 11152 37380
rect 9907 37349 9919 37352
rect 9861 37343 9919 37349
rect 11146 37340 11152 37352
rect 11204 37340 11210 37392
rect 11514 37340 11520 37392
rect 11572 37340 11578 37392
rect 11609 37383 11667 37389
rect 11609 37349 11621 37383
rect 11655 37380 11667 37383
rect 12710 37380 12716 37392
rect 11655 37352 12716 37380
rect 11655 37349 11667 37352
rect 11609 37343 11667 37349
rect 12710 37340 12716 37352
rect 12768 37340 12774 37392
rect 13354 37340 13360 37392
rect 13412 37380 13418 37392
rect 22462 37380 22468 37392
rect 13412 37352 22468 37380
rect 13412 37340 13418 37352
rect 22462 37340 22468 37352
rect 22520 37340 22526 37392
rect 24762 37340 24768 37392
rect 24820 37380 24826 37392
rect 25590 37380 25596 37392
rect 24820 37352 25596 37380
rect 24820 37340 24826 37352
rect 25590 37340 25596 37352
rect 25648 37340 25654 37392
rect 5350 37272 5356 37324
rect 5408 37312 5414 37324
rect 5445 37315 5503 37321
rect 5445 37312 5457 37315
rect 5408 37284 5457 37312
rect 5408 37272 5414 37284
rect 5445 37281 5457 37284
rect 5491 37281 5503 37315
rect 5445 37275 5503 37281
rect 6178 37272 6184 37324
rect 6236 37312 6242 37324
rect 6825 37315 6883 37321
rect 6825 37312 6837 37315
rect 6236 37284 6837 37312
rect 6236 37272 6242 37284
rect 6825 37281 6837 37284
rect 6871 37281 6883 37315
rect 6825 37275 6883 37281
rect 7926 37272 7932 37324
rect 7984 37312 7990 37324
rect 9949 37315 10007 37321
rect 9949 37312 9961 37315
rect 7984 37284 9961 37312
rect 7984 37272 7990 37284
rect 9949 37281 9961 37284
rect 9995 37312 10007 37315
rect 12250 37312 12256 37324
rect 9995 37284 12256 37312
rect 9995 37281 10007 37284
rect 9949 37275 10007 37281
rect 12250 37272 12256 37284
rect 12308 37272 12314 37324
rect 12621 37315 12679 37321
rect 12621 37281 12633 37315
rect 12667 37312 12679 37315
rect 13078 37312 13084 37324
rect 12667 37284 13084 37312
rect 12667 37281 12679 37284
rect 12621 37275 12679 37281
rect 13078 37272 13084 37284
rect 13136 37312 13142 37324
rect 13722 37312 13728 37324
rect 13136 37284 13728 37312
rect 13136 37272 13142 37284
rect 13722 37272 13728 37284
rect 13780 37272 13786 37324
rect 15930 37272 15936 37324
rect 15988 37312 15994 37324
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 15988 37284 16589 37312
rect 15988 37272 15994 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 17126 37272 17132 37324
rect 17184 37272 17190 37324
rect 20533 37315 20591 37321
rect 20533 37312 20545 37315
rect 20364 37284 20545 37312
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 6733 37247 6791 37253
rect 6733 37213 6745 37247
rect 6779 37213 6791 37247
rect 6733 37207 6791 37213
rect 5261 37179 5319 37185
rect 5261 37145 5273 37179
rect 5307 37176 5319 37179
rect 5534 37176 5540 37188
rect 5307 37148 5540 37176
rect 5307 37145 5319 37148
rect 5261 37139 5319 37145
rect 5534 37136 5540 37148
rect 5592 37136 5598 37188
rect 5353 37111 5411 37117
rect 5353 37077 5365 37111
rect 5399 37108 5411 37111
rect 6365 37111 6423 37117
rect 6365 37108 6377 37111
rect 5399 37080 6377 37108
rect 5399 37077 5411 37080
rect 5353 37071 5411 37077
rect 6365 37077 6377 37080
rect 6411 37077 6423 37111
rect 6564 37108 6592 37207
rect 6748 37176 6776 37207
rect 7006 37204 7012 37256
rect 7064 37244 7070 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 7064 37216 7389 37244
rect 7064 37204 7070 37216
rect 7377 37213 7389 37216
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 7653 37247 7711 37253
rect 7653 37213 7665 37247
rect 7699 37213 7711 37247
rect 7653 37207 7711 37213
rect 6914 37176 6920 37188
rect 6748 37148 6920 37176
rect 6914 37136 6920 37148
rect 6972 37136 6978 37188
rect 7668 37176 7696 37207
rect 8202 37204 8208 37256
rect 8260 37204 8266 37256
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9769 37247 9827 37253
rect 9769 37244 9781 37247
rect 9732 37216 9781 37244
rect 9732 37204 9738 37216
rect 9769 37213 9781 37216
rect 9815 37213 9827 37247
rect 9769 37207 9827 37213
rect 10042 37204 10048 37256
rect 10100 37204 10106 37256
rect 10318 37204 10324 37256
rect 10376 37204 10382 37256
rect 11425 37247 11483 37253
rect 11425 37213 11437 37247
rect 11471 37244 11483 37247
rect 11606 37244 11612 37256
rect 11471 37216 11612 37244
rect 11471 37213 11483 37216
rect 11425 37207 11483 37213
rect 11606 37204 11612 37216
rect 11664 37204 11670 37256
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37244 11759 37247
rect 11882 37244 11888 37256
rect 11747 37216 11888 37244
rect 11747 37213 11759 37216
rect 11701 37207 11759 37213
rect 7834 37176 7840 37188
rect 7668 37148 7840 37176
rect 7834 37136 7840 37148
rect 7892 37176 7898 37188
rect 8110 37176 8116 37188
rect 7892 37148 8116 37176
rect 7892 37136 7898 37148
rect 8110 37136 8116 37148
rect 8168 37176 8174 37188
rect 8389 37179 8447 37185
rect 8389 37176 8401 37179
rect 8168 37148 8401 37176
rect 8168 37136 8174 37148
rect 8389 37145 8401 37148
rect 8435 37145 8447 37179
rect 8389 37139 8447 37145
rect 8573 37179 8631 37185
rect 8573 37145 8585 37179
rect 8619 37176 8631 37179
rect 11330 37176 11336 37188
rect 8619 37148 11336 37176
rect 8619 37145 8631 37148
rect 8573 37139 8631 37145
rect 11330 37136 11336 37148
rect 11388 37136 11394 37188
rect 11716 37176 11744 37207
rect 11882 37204 11888 37216
rect 11940 37204 11946 37256
rect 12158 37204 12164 37256
rect 12216 37244 12222 37256
rect 12345 37247 12403 37253
rect 12345 37244 12357 37247
rect 12216 37216 12357 37244
rect 12216 37204 12222 37216
rect 12345 37213 12357 37216
rect 12391 37213 12403 37247
rect 12345 37207 12403 37213
rect 14458 37204 14464 37256
rect 14516 37204 14522 37256
rect 16758 37204 16764 37256
rect 16816 37204 16822 37256
rect 17678 37204 17684 37256
rect 17736 37244 17742 37256
rect 20364 37244 20392 37284
rect 20533 37281 20545 37284
rect 20579 37281 20591 37315
rect 25682 37312 25688 37324
rect 20533 37275 20591 37281
rect 20640 37284 25688 37312
rect 17736 37216 20392 37244
rect 17736 37204 17742 37216
rect 12526 37176 12532 37188
rect 11716 37148 12532 37176
rect 12526 37136 12532 37148
rect 12584 37176 12590 37188
rect 14182 37176 14188 37188
rect 12584 37148 14188 37176
rect 12584 37136 12590 37148
rect 14182 37136 14188 37148
rect 14240 37176 14246 37188
rect 14277 37179 14335 37185
rect 14277 37176 14289 37179
rect 14240 37148 14289 37176
rect 14240 37136 14246 37148
rect 14277 37145 14289 37148
rect 14323 37176 14335 37179
rect 15562 37176 15568 37188
rect 14323 37148 15568 37176
rect 14323 37145 14335 37148
rect 14277 37139 14335 37145
rect 15562 37136 15568 37148
rect 15620 37136 15626 37188
rect 17034 37136 17040 37188
rect 17092 37136 17098 37188
rect 6822 37108 6828 37120
rect 6564 37080 6828 37108
rect 6365 37071 6423 37077
rect 6822 37068 6828 37080
rect 6880 37068 6886 37120
rect 7374 37068 7380 37120
rect 7432 37068 7438 37120
rect 10686 37068 10692 37120
rect 10744 37108 10750 37120
rect 11790 37108 11796 37120
rect 10744 37080 11796 37108
rect 10744 37068 10750 37080
rect 11790 37068 11796 37080
rect 11848 37068 11854 37120
rect 11885 37111 11943 37117
rect 11885 37077 11897 37111
rect 11931 37108 11943 37111
rect 15746 37108 15752 37120
rect 11931 37080 15752 37108
rect 11931 37077 11943 37080
rect 11885 37071 11943 37077
rect 15746 37068 15752 37080
rect 15804 37068 15810 37120
rect 20364 37108 20392 37216
rect 20441 37247 20499 37253
rect 20441 37213 20453 37247
rect 20487 37244 20499 37247
rect 20640 37244 20668 37284
rect 25682 37272 25688 37284
rect 25740 37272 25746 37324
rect 26510 37272 26516 37324
rect 26568 37312 26574 37324
rect 26697 37315 26755 37321
rect 26697 37312 26709 37315
rect 26568 37284 26709 37312
rect 26568 37272 26574 37284
rect 26697 37281 26709 37284
rect 26743 37281 26755 37315
rect 26697 37275 26755 37281
rect 27614 37272 27620 37324
rect 27672 37312 27678 37324
rect 28442 37312 28448 37324
rect 27672 37284 28448 37312
rect 27672 37272 27678 37284
rect 28442 37272 28448 37284
rect 28500 37272 28506 37324
rect 31846 37312 31852 37324
rect 30300 37284 31852 37312
rect 20487 37216 20668 37244
rect 20717 37247 20775 37253
rect 20487 37213 20499 37216
rect 20441 37207 20499 37213
rect 20717 37213 20729 37247
rect 20763 37213 20775 37247
rect 20717 37207 20775 37213
rect 22649 37247 22707 37253
rect 22649 37213 22661 37247
rect 22695 37244 22707 37247
rect 23382 37244 23388 37256
rect 22695 37216 23388 37244
rect 22695 37213 22707 37216
rect 22649 37207 22707 37213
rect 20530 37136 20536 37188
rect 20588 37176 20594 37188
rect 20732 37176 20760 37207
rect 23382 37204 23388 37216
rect 23440 37204 23446 37256
rect 24857 37247 24915 37253
rect 24857 37213 24869 37247
rect 24903 37213 24915 37247
rect 24857 37207 24915 37213
rect 21358 37176 21364 37188
rect 20588 37148 20760 37176
rect 20824 37148 21364 37176
rect 20588 37136 20594 37148
rect 20824 37108 20852 37148
rect 21358 37136 21364 37148
rect 21416 37136 21422 37188
rect 24872 37176 24900 37207
rect 24946 37204 24952 37256
rect 25004 37204 25010 37256
rect 25498 37244 25504 37256
rect 25056 37216 25504 37244
rect 25056 37176 25084 37216
rect 25498 37204 25504 37216
rect 25556 37204 25562 37256
rect 25774 37204 25780 37256
rect 25832 37204 25838 37256
rect 26970 37204 26976 37256
rect 27028 37204 27034 37256
rect 27154 37204 27160 37256
rect 27212 37244 27218 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27212 37216 27813 37244
rect 27212 37204 27218 37216
rect 27801 37213 27813 37216
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 24872 37148 25084 37176
rect 25133 37179 25191 37185
rect 25133 37145 25145 37179
rect 25179 37176 25191 37179
rect 25222 37176 25228 37188
rect 25179 37148 25228 37176
rect 25179 37145 25191 37148
rect 25133 37139 25191 37145
rect 25222 37136 25228 37148
rect 25280 37136 25286 37188
rect 25961 37179 26019 37185
rect 25961 37145 25973 37179
rect 26007 37176 26019 37179
rect 26007 37148 27384 37176
rect 26007 37145 26019 37148
rect 25961 37139 26019 37145
rect 20364 37080 20852 37108
rect 20898 37068 20904 37120
rect 20956 37068 20962 37120
rect 24673 37111 24731 37117
rect 24673 37077 24685 37111
rect 24719 37108 24731 37111
rect 25038 37108 25044 37120
rect 24719 37080 25044 37108
rect 24719 37077 24731 37080
rect 24673 37071 24731 37077
rect 25038 37068 25044 37080
rect 25096 37068 25102 37120
rect 26694 37068 26700 37120
rect 26752 37068 26758 37120
rect 27356 37108 27384 37148
rect 27430 37136 27436 37188
rect 27488 37136 27494 37188
rect 27614 37136 27620 37188
rect 27672 37136 27678 37188
rect 27816 37176 27844 37207
rect 27890 37204 27896 37256
rect 27948 37244 27954 37256
rect 28813 37247 28871 37253
rect 28813 37244 28825 37247
rect 27948 37216 28825 37244
rect 27948 37204 27954 37216
rect 28813 37213 28825 37216
rect 28859 37213 28871 37247
rect 28813 37207 28871 37213
rect 29086 37204 29092 37256
rect 29144 37204 29150 37256
rect 29181 37247 29239 37253
rect 29181 37213 29193 37247
rect 29227 37244 29239 37247
rect 30009 37247 30067 37253
rect 30009 37244 30021 37247
rect 29227 37216 30021 37244
rect 29227 37213 29239 37216
rect 29181 37207 29239 37213
rect 30009 37213 30021 37216
rect 30055 37244 30067 37247
rect 30190 37244 30196 37256
rect 30055 37216 30196 37244
rect 30055 37213 30067 37216
rect 30009 37207 30067 37213
rect 30190 37204 30196 37216
rect 30248 37204 30254 37256
rect 30300 37253 30328 37284
rect 31846 37272 31852 37284
rect 31904 37272 31910 37324
rect 32784 37321 32812 37420
rect 36446 37408 36452 37420
rect 36504 37448 36510 37460
rect 37182 37448 37188 37460
rect 36504 37420 37188 37448
rect 36504 37408 36510 37420
rect 37182 37408 37188 37420
rect 37240 37408 37246 37460
rect 37277 37451 37335 37457
rect 37277 37417 37289 37451
rect 37323 37448 37335 37451
rect 37458 37448 37464 37460
rect 37323 37420 37464 37448
rect 37323 37417 37335 37420
rect 37277 37411 37335 37417
rect 37458 37408 37464 37420
rect 37516 37408 37522 37460
rect 39298 37448 39304 37460
rect 37568 37420 39304 37448
rect 33318 37340 33324 37392
rect 33376 37380 33382 37392
rect 33376 37352 35112 37380
rect 33376 37340 33382 37352
rect 35084 37321 35112 37352
rect 35802 37340 35808 37392
rect 35860 37380 35866 37392
rect 37568 37380 37596 37420
rect 39298 37408 39304 37420
rect 39356 37408 39362 37460
rect 39482 37408 39488 37460
rect 39540 37408 39546 37460
rect 35860 37352 37596 37380
rect 35860 37340 35866 37352
rect 37642 37340 37648 37392
rect 37700 37380 37706 37392
rect 40494 37380 40500 37392
rect 37700 37352 40500 37380
rect 37700 37340 37706 37352
rect 40494 37340 40500 37352
rect 40552 37380 40558 37392
rect 41414 37380 41420 37392
rect 40552 37352 41420 37380
rect 40552 37340 40558 37352
rect 41414 37340 41420 37352
rect 41472 37340 41478 37392
rect 32769 37315 32827 37321
rect 32769 37281 32781 37315
rect 32815 37281 32827 37315
rect 32769 37275 32827 37281
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 35434 37312 35440 37324
rect 35115 37284 35440 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 35434 37272 35440 37284
rect 35492 37272 35498 37324
rect 38286 37312 38292 37324
rect 36648 37284 38292 37312
rect 30285 37247 30343 37253
rect 30285 37213 30297 37247
rect 30331 37213 30343 37247
rect 30285 37207 30343 37213
rect 32030 37204 32036 37256
rect 32088 37244 32094 37256
rect 32125 37247 32183 37253
rect 32125 37244 32137 37247
rect 32088 37216 32137 37244
rect 32088 37204 32094 37216
rect 32125 37213 32137 37216
rect 32171 37213 32183 37247
rect 32125 37207 32183 37213
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37244 32367 37247
rect 32490 37244 32496 37256
rect 32355 37216 32496 37244
rect 32355 37213 32367 37216
rect 32309 37207 32367 37213
rect 32490 37204 32496 37216
rect 32548 37204 32554 37256
rect 32674 37204 32680 37256
rect 32732 37204 32738 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33060 37216 33793 37244
rect 31297 37179 31355 37185
rect 31297 37176 31309 37179
rect 27816 37148 31309 37176
rect 31297 37145 31309 37148
rect 31343 37145 31355 37179
rect 31297 37139 31355 37145
rect 28718 37108 28724 37120
rect 27356 37080 28724 37108
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 28810 37068 28816 37120
rect 28868 37108 28874 37120
rect 29825 37111 29883 37117
rect 29825 37108 29837 37111
rect 28868 37080 29837 37108
rect 28868 37068 28874 37080
rect 29825 37077 29837 37080
rect 29871 37077 29883 37111
rect 31312 37108 31340 37139
rect 31478 37136 31484 37188
rect 31536 37136 31542 37188
rect 31570 37136 31576 37188
rect 31628 37176 31634 37188
rect 31665 37179 31723 37185
rect 31665 37176 31677 37179
rect 31628 37148 31677 37176
rect 31628 37136 31634 37148
rect 31665 37145 31677 37148
rect 31711 37145 31723 37179
rect 31665 37139 31723 37145
rect 32766 37108 32772 37120
rect 31312 37080 32772 37108
rect 29825 37071 29883 37077
rect 32766 37068 32772 37080
rect 32824 37108 32830 37120
rect 33060 37108 33088 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 33870 37204 33876 37256
rect 33928 37204 33934 37256
rect 33962 37204 33968 37256
rect 34020 37204 34026 37256
rect 34238 37204 34244 37256
rect 34296 37244 34302 37256
rect 35253 37247 35311 37253
rect 35253 37244 35265 37247
rect 34296 37216 35265 37244
rect 34296 37204 34302 37216
rect 35253 37213 35265 37216
rect 35299 37213 35311 37247
rect 35253 37207 35311 37213
rect 35710 37204 35716 37256
rect 35768 37204 35774 37256
rect 36648 37253 36676 37284
rect 38286 37272 38292 37284
rect 38344 37272 38350 37324
rect 38654 37272 38660 37324
rect 38712 37312 38718 37324
rect 38712 37284 39252 37312
rect 38712 37272 38718 37284
rect 37182 37253 37188 37256
rect 36633 37247 36691 37253
rect 36633 37213 36645 37247
rect 36679 37213 36691 37247
rect 36633 37207 36691 37213
rect 36726 37247 36784 37253
rect 36726 37213 36738 37247
rect 36772 37213 36784 37247
rect 36726 37207 36784 37213
rect 37139 37247 37188 37253
rect 37139 37213 37151 37247
rect 37185 37213 37188 37247
rect 37139 37207 37188 37213
rect 33321 37179 33379 37185
rect 33321 37145 33333 37179
rect 33367 37176 33379 37179
rect 33367 37148 35480 37176
rect 33367 37145 33379 37148
rect 33321 37139 33379 37145
rect 32824 37080 33088 37108
rect 35452 37108 35480 37148
rect 35526 37136 35532 37188
rect 35584 37176 35590 37188
rect 36740 37176 36768 37207
rect 37182 37204 37188 37207
rect 37240 37204 37246 37256
rect 39224 37253 39252 37284
rect 38933 37247 38991 37253
rect 38933 37213 38945 37247
rect 38979 37213 38991 37247
rect 38933 37207 38991 37213
rect 39209 37247 39267 37253
rect 39209 37213 39221 37247
rect 39255 37213 39267 37247
rect 39209 37207 39267 37213
rect 39301 37247 39359 37253
rect 39301 37213 39313 37247
rect 39347 37244 39359 37247
rect 39390 37244 39396 37256
rect 39347 37216 39396 37244
rect 39347 37213 39359 37216
rect 39301 37207 39359 37213
rect 35584 37148 36768 37176
rect 35584 37136 35590 37148
rect 36630 37108 36636 37120
rect 35452 37080 36636 37108
rect 32824 37068 32830 37080
rect 36630 37068 36636 37080
rect 36688 37068 36694 37120
rect 36740 37108 36768 37148
rect 36906 37136 36912 37188
rect 36964 37136 36970 37188
rect 37001 37179 37059 37185
rect 37001 37145 37013 37179
rect 37047 37176 37059 37179
rect 37274 37176 37280 37188
rect 37047 37148 37280 37176
rect 37047 37145 37059 37148
rect 37001 37139 37059 37145
rect 37274 37136 37280 37148
rect 37332 37176 37338 37188
rect 38948 37176 38976 37207
rect 37332 37148 38976 37176
rect 37332 37136 37338 37148
rect 39114 37136 39120 37188
rect 39172 37136 39178 37188
rect 39224 37176 39252 37207
rect 39390 37204 39396 37216
rect 39448 37204 39454 37256
rect 39482 37204 39488 37256
rect 39540 37244 39546 37256
rect 40129 37247 40187 37253
rect 40129 37244 40141 37247
rect 39540 37216 40141 37244
rect 39540 37204 39546 37216
rect 40129 37213 40141 37216
rect 40175 37213 40187 37247
rect 40129 37207 40187 37213
rect 40222 37247 40280 37253
rect 40222 37213 40234 37247
rect 40268 37213 40280 37247
rect 40222 37207 40280 37213
rect 39850 37176 39856 37188
rect 39224 37148 39856 37176
rect 39850 37136 39856 37148
rect 39908 37136 39914 37188
rect 40236 37108 40264 37207
rect 40494 37204 40500 37256
rect 40552 37204 40558 37256
rect 40635 37247 40693 37253
rect 40635 37213 40647 37247
rect 40681 37244 40693 37247
rect 41138 37244 41144 37256
rect 40681 37216 41144 37244
rect 40681 37213 40693 37216
rect 40635 37207 40693 37213
rect 41138 37204 41144 37216
rect 41196 37204 41202 37256
rect 41693 37247 41751 37253
rect 41693 37213 41705 37247
rect 41739 37244 41751 37247
rect 41782 37244 41788 37256
rect 41739 37216 41788 37244
rect 41739 37213 41751 37216
rect 41693 37207 41751 37213
rect 41782 37204 41788 37216
rect 41840 37204 41846 37256
rect 41892 37216 42748 37244
rect 40402 37136 40408 37188
rect 40460 37136 40466 37188
rect 41892 37176 41920 37216
rect 40512 37148 41920 37176
rect 41960 37179 42018 37185
rect 40512 37108 40540 37148
rect 41960 37145 41972 37179
rect 42006 37176 42018 37179
rect 42610 37176 42616 37188
rect 42006 37148 42616 37176
rect 42006 37145 42018 37148
rect 41960 37139 42018 37145
rect 42610 37136 42616 37148
rect 42668 37136 42674 37188
rect 42720 37176 42748 37216
rect 42720 37148 43116 37176
rect 43088 37120 43116 37148
rect 36740 37080 40540 37108
rect 40773 37111 40831 37117
rect 40773 37077 40785 37111
rect 40819 37108 40831 37111
rect 42978 37108 42984 37120
rect 40819 37080 42984 37108
rect 40819 37077 40831 37080
rect 40773 37071 40831 37077
rect 42978 37068 42984 37080
rect 43036 37068 43042 37120
rect 43070 37068 43076 37120
rect 43128 37068 43134 37120
rect 1104 37018 43884 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 43884 37018
rect 1104 36944 43884 36966
rect 8110 36904 8116 36916
rect 6656 36876 8116 36904
rect 6656 36845 6684 36876
rect 8110 36864 8116 36876
rect 8168 36864 8174 36916
rect 9950 36864 9956 36916
rect 10008 36904 10014 36916
rect 12342 36904 12348 36916
rect 10008 36876 12348 36904
rect 10008 36864 10014 36876
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 13725 36907 13783 36913
rect 13725 36873 13737 36907
rect 13771 36904 13783 36907
rect 13998 36904 14004 36916
rect 13771 36876 14004 36904
rect 13771 36873 13783 36876
rect 13725 36867 13783 36873
rect 13998 36864 14004 36876
rect 14056 36864 14062 36916
rect 15010 36904 15016 36916
rect 14108 36876 15016 36904
rect 6641 36839 6699 36845
rect 6641 36805 6653 36839
rect 6687 36805 6699 36839
rect 10686 36836 10692 36848
rect 6641 36799 6699 36805
rect 6840 36808 7880 36836
rect 6840 36777 6868 36808
rect 7852 36780 7880 36808
rect 9140 36808 10692 36836
rect 6825 36771 6883 36777
rect 6825 36737 6837 36771
rect 6871 36737 6883 36771
rect 6825 36731 6883 36737
rect 6917 36771 6975 36777
rect 6917 36737 6929 36771
rect 6963 36737 6975 36771
rect 6917 36731 6975 36737
rect 6932 36632 6960 36731
rect 7834 36728 7840 36780
rect 7892 36728 7898 36780
rect 8018 36728 8024 36780
rect 8076 36728 8082 36780
rect 8938 36728 8944 36780
rect 8996 36728 9002 36780
rect 9140 36777 9168 36808
rect 10686 36796 10692 36808
rect 10744 36796 10750 36848
rect 14108 36836 14136 36876
rect 15010 36864 15016 36876
rect 15068 36864 15074 36916
rect 15841 36907 15899 36913
rect 15841 36873 15853 36907
rect 15887 36904 15899 36907
rect 17126 36904 17132 36916
rect 15887 36876 17132 36904
rect 15887 36873 15899 36876
rect 15841 36867 15899 36873
rect 17126 36864 17132 36876
rect 17184 36864 17190 36916
rect 20257 36907 20315 36913
rect 20257 36873 20269 36907
rect 20303 36904 20315 36907
rect 20622 36904 20628 36916
rect 20303 36876 20628 36904
rect 20303 36873 20315 36876
rect 20257 36867 20315 36873
rect 20622 36864 20628 36876
rect 20680 36864 20686 36916
rect 24578 36864 24584 36916
rect 24636 36904 24642 36916
rect 24673 36907 24731 36913
rect 24673 36904 24685 36907
rect 24636 36876 24685 36904
rect 24636 36864 24642 36876
rect 24673 36873 24685 36876
rect 24719 36873 24731 36907
rect 33134 36904 33140 36916
rect 24673 36867 24731 36873
rect 27724 36876 33140 36904
rect 16482 36836 16488 36848
rect 11900 36808 14136 36836
rect 15488 36808 16488 36836
rect 9125 36771 9183 36777
rect 9125 36737 9137 36771
rect 9171 36737 9183 36771
rect 9125 36731 9183 36737
rect 9217 36771 9275 36777
rect 9217 36737 9229 36771
rect 9263 36768 9275 36771
rect 9674 36768 9680 36780
rect 9263 36740 9680 36768
rect 9263 36737 9275 36740
rect 9217 36731 9275 36737
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 10226 36728 10232 36780
rect 10284 36768 10290 36780
rect 10321 36771 10379 36777
rect 10321 36768 10333 36771
rect 10284 36740 10333 36768
rect 10284 36728 10290 36740
rect 10321 36737 10333 36740
rect 10367 36737 10379 36771
rect 10321 36731 10379 36737
rect 10410 36728 10416 36780
rect 10468 36768 10474 36780
rect 11072 36777 11284 36790
rect 10965 36771 11023 36777
rect 10965 36768 10977 36771
rect 10468 36740 10977 36768
rect 10468 36728 10474 36740
rect 10965 36737 10977 36740
rect 11011 36737 11023 36771
rect 10965 36731 11023 36737
rect 11057 36774 11284 36777
rect 11057 36771 11376 36774
rect 11057 36737 11069 36771
rect 11103 36768 11376 36771
rect 11422 36768 11428 36780
rect 11103 36762 11428 36768
rect 11103 36737 11115 36762
rect 11256 36746 11428 36762
rect 11348 36740 11428 36746
rect 11057 36731 11115 36737
rect 8202 36660 8208 36712
rect 8260 36700 8266 36712
rect 9033 36703 9091 36709
rect 9033 36700 9045 36703
rect 8260 36672 9045 36700
rect 8260 36660 8266 36672
rect 9033 36669 9045 36672
rect 9079 36669 9091 36703
rect 9033 36663 9091 36669
rect 10042 36660 10048 36712
rect 10100 36660 10106 36712
rect 10502 36660 10508 36712
rect 10560 36700 10566 36712
rect 10781 36703 10839 36709
rect 10781 36700 10793 36703
rect 10560 36672 10793 36700
rect 10560 36660 10566 36672
rect 10781 36669 10793 36672
rect 10827 36669 10839 36703
rect 10980 36700 11008 36731
rect 11422 36728 11428 36740
rect 11480 36768 11486 36780
rect 11900 36768 11928 36808
rect 15488 36780 15516 36808
rect 16482 36796 16488 36808
rect 16540 36796 16546 36848
rect 16574 36796 16580 36848
rect 16632 36836 16638 36848
rect 17589 36839 17647 36845
rect 17589 36836 17601 36839
rect 16632 36808 17601 36836
rect 16632 36796 16638 36808
rect 17589 36805 17601 36808
rect 17635 36805 17647 36839
rect 17589 36799 17647 36805
rect 17862 36796 17868 36848
rect 17920 36836 17926 36848
rect 22002 36836 22008 36848
rect 17920 36808 22008 36836
rect 17920 36796 17926 36808
rect 22002 36796 22008 36808
rect 22060 36796 22066 36848
rect 25866 36836 25872 36848
rect 24044 36808 25872 36836
rect 11480 36740 11928 36768
rect 11480 36728 11486 36740
rect 12618 36728 12624 36780
rect 12676 36768 12682 36780
rect 12713 36771 12771 36777
rect 12713 36768 12725 36771
rect 12676 36740 12725 36768
rect 12676 36728 12682 36740
rect 12713 36737 12725 36740
rect 12759 36768 12771 36771
rect 13078 36768 13084 36780
rect 12759 36740 13084 36768
rect 12759 36737 12771 36740
rect 12713 36731 12771 36737
rect 13078 36728 13084 36740
rect 13136 36728 13142 36780
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36768 13599 36771
rect 13630 36768 13636 36780
rect 13587 36740 13636 36768
rect 13587 36737 13599 36740
rect 13541 36731 13599 36737
rect 13630 36728 13636 36740
rect 13688 36728 13694 36780
rect 14642 36728 14648 36780
rect 14700 36777 14706 36780
rect 14700 36731 14708 36777
rect 14700 36728 14706 36731
rect 15470 36728 15476 36780
rect 15528 36728 15534 36780
rect 15562 36728 15568 36780
rect 15620 36728 15626 36780
rect 16850 36728 16856 36780
rect 16908 36728 16914 36780
rect 17034 36728 17040 36780
rect 17092 36768 17098 36780
rect 17221 36771 17279 36777
rect 17221 36768 17233 36771
rect 17092 36740 17233 36768
rect 17092 36728 17098 36740
rect 17221 36737 17233 36740
rect 17267 36737 17279 36771
rect 17221 36731 17279 36737
rect 17313 36771 17371 36777
rect 17313 36737 17325 36771
rect 17359 36737 17371 36771
rect 17313 36731 17371 36737
rect 11977 36703 12035 36709
rect 11977 36700 11989 36703
rect 10980 36672 11989 36700
rect 10781 36663 10839 36669
rect 11977 36669 11989 36672
rect 12023 36669 12035 36703
rect 11977 36663 12035 36669
rect 13265 36703 13323 36709
rect 13265 36669 13277 36703
rect 13311 36700 13323 36703
rect 13311 36672 14596 36700
rect 13311 36669 13323 36672
rect 13265 36663 13323 36669
rect 8846 36632 8852 36644
rect 6932 36604 8852 36632
rect 8846 36592 8852 36604
rect 8904 36592 8910 36644
rect 9766 36592 9772 36644
rect 9824 36632 9830 36644
rect 11422 36632 11428 36644
rect 9824 36604 11428 36632
rect 9824 36592 9830 36604
rect 11422 36592 11428 36604
rect 11480 36592 11486 36644
rect 13280 36632 13308 36663
rect 12406 36604 13308 36632
rect 6730 36524 6736 36576
rect 6788 36524 6794 36576
rect 7101 36567 7159 36573
rect 7101 36533 7113 36567
rect 7147 36564 7159 36567
rect 7282 36564 7288 36576
rect 7147 36536 7288 36564
rect 7147 36533 7159 36536
rect 7101 36527 7159 36533
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 7558 36524 7564 36576
rect 7616 36564 7622 36576
rect 7653 36567 7711 36573
rect 7653 36564 7665 36567
rect 7616 36536 7665 36564
rect 7616 36524 7622 36536
rect 7653 36533 7665 36536
rect 7699 36533 7711 36567
rect 7653 36527 7711 36533
rect 9401 36567 9459 36573
rect 9401 36533 9413 36567
rect 9447 36564 9459 36567
rect 10870 36564 10876 36576
rect 9447 36536 10876 36564
rect 9447 36533 9459 36536
rect 9401 36527 9459 36533
rect 10870 36524 10876 36536
rect 10928 36524 10934 36576
rect 10962 36524 10968 36576
rect 11020 36564 11026 36576
rect 12406 36564 12434 36604
rect 14568 36576 14596 36672
rect 14734 36660 14740 36712
rect 14792 36660 14798 36712
rect 15746 36632 15752 36644
rect 14844 36604 15752 36632
rect 11020 36536 12434 36564
rect 11020 36524 11026 36536
rect 12986 36524 12992 36576
rect 13044 36564 13050 36576
rect 13357 36567 13415 36573
rect 13357 36564 13369 36567
rect 13044 36536 13369 36564
rect 13044 36524 13050 36536
rect 13357 36533 13369 36536
rect 13403 36533 13415 36567
rect 13357 36527 13415 36533
rect 14550 36524 14556 36576
rect 14608 36564 14614 36576
rect 14844 36573 14872 36604
rect 15746 36592 15752 36604
rect 15804 36592 15810 36644
rect 15838 36592 15844 36644
rect 15896 36632 15902 36644
rect 17328 36632 17356 36731
rect 19150 36728 19156 36780
rect 19208 36728 19214 36780
rect 20625 36771 20683 36777
rect 20625 36768 20637 36771
rect 19260 36740 20637 36768
rect 17770 36660 17776 36712
rect 17828 36700 17834 36712
rect 19260 36700 19288 36740
rect 20625 36737 20637 36740
rect 20671 36737 20683 36771
rect 20625 36731 20683 36737
rect 22094 36728 22100 36780
rect 22152 36728 22158 36780
rect 22278 36728 22284 36780
rect 22336 36728 22342 36780
rect 24044 36777 24072 36808
rect 25866 36796 25872 36808
rect 25924 36836 25930 36848
rect 27522 36836 27528 36848
rect 25924 36808 27528 36836
rect 25924 36796 25930 36808
rect 27522 36796 27528 36808
rect 27580 36796 27586 36848
rect 24029 36771 24087 36777
rect 24029 36737 24041 36771
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 24213 36771 24271 36777
rect 24213 36737 24225 36771
rect 24259 36737 24271 36771
rect 24213 36731 24271 36737
rect 17828 36672 19288 36700
rect 17828 36660 17834 36672
rect 19426 36660 19432 36712
rect 19484 36660 19490 36712
rect 20530 36660 20536 36712
rect 20588 36660 20594 36712
rect 20806 36660 20812 36712
rect 20864 36700 20870 36712
rect 22005 36703 22063 36709
rect 22005 36700 22017 36703
rect 20864 36672 22017 36700
rect 20864 36660 20870 36672
rect 22005 36669 22017 36672
rect 22051 36669 22063 36703
rect 24228 36700 24256 36731
rect 24854 36728 24860 36780
rect 24912 36728 24918 36780
rect 25038 36728 25044 36780
rect 25096 36728 25102 36780
rect 27338 36728 27344 36780
rect 27396 36728 27402 36780
rect 27724 36777 27752 36876
rect 33134 36864 33140 36876
rect 33192 36864 33198 36916
rect 34422 36864 34428 36916
rect 34480 36904 34486 36916
rect 34480 36876 36308 36904
rect 34480 36864 34486 36876
rect 30374 36836 30380 36848
rect 30024 36808 30380 36836
rect 30024 36777 30052 36808
rect 30374 36796 30380 36808
rect 30432 36836 30438 36848
rect 30432 36808 32904 36836
rect 30432 36796 30438 36808
rect 27709 36771 27767 36777
rect 27709 36737 27721 36771
rect 27755 36737 27767 36771
rect 27709 36731 27767 36737
rect 29733 36771 29791 36777
rect 29733 36737 29745 36771
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 30009 36771 30067 36777
rect 30009 36737 30021 36771
rect 30055 36737 30067 36771
rect 30009 36731 30067 36737
rect 27154 36700 27160 36712
rect 24228 36672 27160 36700
rect 22005 36663 22063 36669
rect 27154 36660 27160 36672
rect 27212 36660 27218 36712
rect 27249 36703 27307 36709
rect 27249 36669 27261 36703
rect 27295 36700 27307 36703
rect 27522 36700 27528 36712
rect 27295 36672 27528 36700
rect 27295 36669 27307 36672
rect 27249 36663 27307 36669
rect 27522 36660 27528 36672
rect 27580 36660 27586 36712
rect 28810 36700 28816 36712
rect 27632 36672 28816 36700
rect 18874 36632 18880 36644
rect 15896 36604 18880 36632
rect 15896 36592 15902 36604
rect 18874 36592 18880 36604
rect 18932 36592 18938 36644
rect 20640 36604 22508 36632
rect 14829 36567 14887 36573
rect 14829 36564 14841 36567
rect 14608 36536 14841 36564
rect 14608 36524 14614 36536
rect 14829 36533 14841 36536
rect 14875 36533 14887 36567
rect 14829 36527 14887 36533
rect 15010 36524 15016 36576
rect 15068 36524 15074 36576
rect 15102 36524 15108 36576
rect 15160 36564 15166 36576
rect 15473 36567 15531 36573
rect 15473 36564 15485 36567
rect 15160 36536 15485 36564
rect 15160 36524 15166 36536
rect 15473 36533 15485 36536
rect 15519 36533 15531 36567
rect 15473 36527 15531 36533
rect 15562 36524 15568 36576
rect 15620 36564 15626 36576
rect 16390 36564 16396 36576
rect 15620 36536 16396 36564
rect 15620 36524 15626 36536
rect 16390 36524 16396 36536
rect 16448 36564 16454 36576
rect 20640 36573 20668 36604
rect 22480 36576 22508 36604
rect 24854 36592 24860 36644
rect 24912 36632 24918 36644
rect 24912 36604 26004 36632
rect 24912 36592 24918 36604
rect 25976 36576 26004 36604
rect 16945 36567 17003 36573
rect 16945 36564 16957 36567
rect 16448 36536 16957 36564
rect 16448 36524 16454 36536
rect 16945 36533 16957 36536
rect 16991 36533 17003 36567
rect 16945 36527 17003 36533
rect 20625 36567 20683 36573
rect 20625 36533 20637 36567
rect 20671 36533 20683 36567
rect 20625 36527 20683 36533
rect 22462 36524 22468 36576
rect 22520 36524 22526 36576
rect 23658 36524 23664 36576
rect 23716 36564 23722 36576
rect 24213 36567 24271 36573
rect 24213 36564 24225 36567
rect 23716 36536 24225 36564
rect 23716 36524 23722 36536
rect 24213 36533 24225 36536
rect 24259 36533 24271 36567
rect 24213 36527 24271 36533
rect 25041 36567 25099 36573
rect 25041 36533 25053 36567
rect 25087 36564 25099 36567
rect 25590 36564 25596 36576
rect 25087 36536 25596 36564
rect 25087 36533 25099 36536
rect 25041 36527 25099 36533
rect 25590 36524 25596 36536
rect 25648 36524 25654 36576
rect 25958 36524 25964 36576
rect 26016 36564 26022 36576
rect 27632 36564 27660 36672
rect 28810 36660 28816 36672
rect 28868 36660 28874 36712
rect 29748 36632 29776 36731
rect 31018 36728 31024 36780
rect 31076 36728 31082 36780
rect 31205 36771 31263 36777
rect 31205 36737 31217 36771
rect 31251 36737 31263 36771
rect 31205 36731 31263 36737
rect 29914 36660 29920 36712
rect 29972 36660 29978 36712
rect 30742 36660 30748 36712
rect 30800 36660 30806 36712
rect 31036 36632 31064 36728
rect 29748 36604 31064 36632
rect 31220 36700 31248 36731
rect 31662 36728 31668 36780
rect 31720 36768 31726 36780
rect 32309 36771 32367 36777
rect 32309 36768 32321 36771
rect 31720 36740 32321 36768
rect 31720 36728 31726 36740
rect 32309 36737 32321 36740
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 32582 36728 32588 36780
rect 32640 36728 32646 36780
rect 32876 36700 32904 36808
rect 33042 36796 33048 36848
rect 33100 36836 33106 36848
rect 33100 36808 34560 36836
rect 33100 36796 33106 36808
rect 33410 36728 33416 36780
rect 33468 36768 33474 36780
rect 33505 36771 33563 36777
rect 33505 36768 33517 36771
rect 33468 36740 33517 36768
rect 33468 36728 33474 36740
rect 33505 36737 33517 36740
rect 33551 36737 33563 36771
rect 33505 36731 33563 36737
rect 33594 36728 33600 36780
rect 33652 36768 33658 36780
rect 33689 36771 33747 36777
rect 33689 36768 33701 36771
rect 33652 36740 33701 36768
rect 33652 36728 33658 36740
rect 33689 36737 33701 36740
rect 33735 36737 33747 36771
rect 33689 36731 33747 36737
rect 34054 36728 34060 36780
rect 34112 36768 34118 36780
rect 34532 36777 34560 36808
rect 34790 36796 34796 36848
rect 34848 36836 34854 36848
rect 34848 36808 34928 36836
rect 34848 36796 34854 36808
rect 34900 36777 34928 36808
rect 34333 36771 34391 36777
rect 34333 36768 34345 36771
rect 34112 36740 34345 36768
rect 34112 36728 34118 36740
rect 34333 36737 34345 36740
rect 34379 36737 34391 36771
rect 34333 36731 34391 36737
rect 34517 36771 34575 36777
rect 34517 36737 34529 36771
rect 34563 36737 34575 36771
rect 34517 36731 34575 36737
rect 34885 36771 34943 36777
rect 34885 36737 34897 36771
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 36173 36771 36231 36777
rect 36173 36737 36185 36771
rect 36219 36737 36231 36771
rect 36280 36768 36308 36876
rect 36630 36864 36636 36916
rect 36688 36904 36694 36916
rect 39114 36904 39120 36916
rect 36688 36876 39120 36904
rect 36688 36864 36694 36876
rect 39114 36864 39120 36876
rect 39172 36904 39178 36916
rect 39942 36904 39948 36916
rect 39172 36876 39948 36904
rect 39172 36864 39178 36876
rect 39942 36864 39948 36876
rect 40000 36864 40006 36916
rect 42610 36864 42616 36916
rect 42668 36864 42674 36916
rect 42978 36864 42984 36916
rect 43036 36904 43042 36916
rect 43073 36907 43131 36913
rect 43073 36904 43085 36907
rect 43036 36876 43085 36904
rect 43036 36864 43042 36876
rect 43073 36873 43085 36876
rect 43119 36873 43131 36907
rect 43073 36867 43131 36873
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 36280 36740 36369 36768
rect 36173 36731 36231 36737
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 36541 36771 36599 36777
rect 36541 36737 36553 36771
rect 36587 36768 36599 36771
rect 41598 36768 41604 36780
rect 36587 36740 41604 36768
rect 36587 36737 36599 36740
rect 36541 36731 36599 36737
rect 33045 36703 33103 36709
rect 33045 36700 33057 36703
rect 31220 36672 32536 36700
rect 32876 36672 33057 36700
rect 26016 36536 27660 36564
rect 26016 36524 26022 36536
rect 27706 36524 27712 36576
rect 27764 36524 27770 36576
rect 27893 36567 27951 36573
rect 27893 36533 27905 36567
rect 27939 36564 27951 36567
rect 27982 36564 27988 36576
rect 27939 36536 27988 36564
rect 27939 36533 27951 36536
rect 27893 36527 27951 36533
rect 27982 36524 27988 36536
rect 28040 36524 28046 36576
rect 28074 36524 28080 36576
rect 28132 36564 28138 36576
rect 31220 36564 31248 36672
rect 32401 36635 32459 36641
rect 32401 36601 32413 36635
rect 32447 36601 32459 36635
rect 32508 36632 32536 36672
rect 33045 36669 33057 36672
rect 33091 36700 33103 36703
rect 34238 36700 34244 36712
rect 33091 36672 34244 36700
rect 33091 36669 33103 36672
rect 33045 36663 33103 36669
rect 34238 36660 34244 36672
rect 34296 36660 34302 36712
rect 34790 36660 34796 36712
rect 34848 36660 34854 36712
rect 36188 36700 36216 36731
rect 41598 36728 41604 36740
rect 41656 36728 41662 36780
rect 42981 36771 43039 36777
rect 42981 36737 42993 36771
rect 43027 36768 43039 36771
rect 43070 36768 43076 36780
rect 43027 36740 43076 36768
rect 43027 36737 43039 36740
rect 42981 36731 43039 36737
rect 43070 36728 43076 36740
rect 43128 36728 43134 36780
rect 36814 36700 36820 36712
rect 36188 36672 36820 36700
rect 36814 36660 36820 36672
rect 36872 36660 36878 36712
rect 43162 36660 43168 36712
rect 43220 36660 43226 36712
rect 33410 36632 33416 36644
rect 32508 36604 33416 36632
rect 32401 36595 32459 36601
rect 28132 36536 31248 36564
rect 28132 36524 28138 36536
rect 31478 36524 31484 36576
rect 31536 36564 31542 36576
rect 32416 36564 32444 36595
rect 33410 36592 33416 36604
rect 33468 36592 33474 36644
rect 33781 36635 33839 36641
rect 33781 36601 33793 36635
rect 33827 36632 33839 36635
rect 34808 36632 34836 36660
rect 33827 36604 34836 36632
rect 33827 36601 33839 36604
rect 33781 36595 33839 36601
rect 31536 36536 32444 36564
rect 35437 36567 35495 36573
rect 31536 36524 31542 36536
rect 35437 36533 35449 36567
rect 35483 36564 35495 36567
rect 37826 36564 37832 36576
rect 35483 36536 37832 36564
rect 35483 36533 35495 36536
rect 35437 36527 35495 36533
rect 37826 36524 37832 36536
rect 37884 36524 37890 36576
rect 1104 36474 43884 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 43884 36474
rect 1104 36400 43884 36422
rect 6730 36320 6736 36372
rect 6788 36360 6794 36372
rect 9950 36360 9956 36372
rect 6788 36332 9956 36360
rect 6788 36320 6794 36332
rect 9950 36320 9956 36332
rect 10008 36320 10014 36372
rect 11514 36360 11520 36372
rect 10244 36332 11520 36360
rect 10244 36304 10272 36332
rect 11514 36320 11520 36332
rect 11572 36320 11578 36372
rect 11698 36320 11704 36372
rect 11756 36360 11762 36372
rect 12437 36363 12495 36369
rect 12437 36360 12449 36363
rect 11756 36332 12449 36360
rect 11756 36320 11762 36332
rect 12437 36329 12449 36332
rect 12483 36329 12495 36363
rect 12437 36323 12495 36329
rect 13630 36320 13636 36372
rect 13688 36320 13694 36372
rect 14550 36320 14556 36372
rect 14608 36320 14614 36372
rect 14737 36363 14795 36369
rect 14737 36329 14749 36363
rect 14783 36360 14795 36363
rect 15838 36360 15844 36372
rect 14783 36332 15844 36360
rect 14783 36329 14795 36332
rect 14737 36323 14795 36329
rect 15838 36320 15844 36332
rect 15896 36320 15902 36372
rect 16022 36320 16028 36372
rect 16080 36320 16086 36372
rect 17126 36320 17132 36372
rect 17184 36320 17190 36372
rect 17221 36363 17279 36369
rect 17221 36329 17233 36363
rect 17267 36360 17279 36363
rect 17678 36360 17684 36372
rect 17267 36332 17684 36360
rect 17267 36329 17279 36332
rect 17221 36323 17279 36329
rect 17678 36320 17684 36332
rect 17736 36320 17742 36372
rect 17770 36320 17776 36372
rect 17828 36320 17834 36372
rect 17862 36320 17868 36372
rect 17920 36360 17926 36372
rect 18509 36363 18567 36369
rect 18509 36360 18521 36363
rect 17920 36332 18521 36360
rect 17920 36320 17926 36332
rect 18509 36329 18521 36332
rect 18555 36329 18567 36363
rect 18509 36323 18567 36329
rect 19058 36320 19064 36372
rect 19116 36360 19122 36372
rect 19886 36360 19892 36372
rect 19116 36332 19892 36360
rect 19116 36320 19122 36332
rect 19886 36320 19892 36332
rect 19944 36320 19950 36372
rect 19981 36363 20039 36369
rect 19981 36329 19993 36363
rect 20027 36360 20039 36363
rect 20346 36360 20352 36372
rect 20027 36332 20352 36360
rect 20027 36329 20039 36332
rect 19981 36323 20039 36329
rect 20346 36320 20352 36332
rect 20404 36320 20410 36372
rect 20530 36320 20536 36372
rect 20588 36360 20594 36372
rect 21177 36363 21235 36369
rect 21177 36360 21189 36363
rect 20588 36332 21189 36360
rect 20588 36320 20594 36332
rect 21177 36329 21189 36332
rect 21223 36329 21235 36363
rect 21177 36323 21235 36329
rect 22462 36320 22468 36372
rect 22520 36360 22526 36372
rect 23477 36363 23535 36369
rect 23477 36360 23489 36363
rect 22520 36332 23489 36360
rect 22520 36320 22526 36332
rect 23477 36329 23489 36332
rect 23523 36329 23535 36363
rect 23477 36323 23535 36329
rect 23750 36320 23756 36372
rect 23808 36360 23814 36372
rect 23937 36363 23995 36369
rect 23937 36360 23949 36363
rect 23808 36332 23949 36360
rect 23808 36320 23814 36332
rect 23937 36329 23949 36332
rect 23983 36329 23995 36363
rect 23937 36323 23995 36329
rect 24596 36332 25084 36360
rect 8018 36252 8024 36304
rect 8076 36292 8082 36304
rect 10226 36292 10232 36304
rect 8076 36264 10232 36292
rect 8076 36252 8082 36264
rect 10226 36252 10232 36264
rect 10284 36252 10290 36304
rect 10502 36252 10508 36304
rect 10560 36252 10566 36304
rect 11054 36252 11060 36304
rect 11112 36292 11118 36304
rect 12802 36292 12808 36304
rect 11112 36264 12808 36292
rect 11112 36252 11118 36264
rect 12802 36252 12808 36264
rect 12860 36292 12866 36304
rect 15562 36292 15568 36304
rect 12860 36264 15568 36292
rect 12860 36252 12866 36264
rect 15562 36252 15568 36264
rect 15620 36252 15626 36304
rect 15654 36252 15660 36304
rect 15712 36252 15718 36304
rect 15930 36252 15936 36304
rect 15988 36292 15994 36304
rect 16209 36295 16267 36301
rect 16209 36292 16221 36295
rect 15988 36264 16221 36292
rect 15988 36252 15994 36264
rect 16209 36261 16221 36264
rect 16255 36261 16267 36295
rect 20947 36295 21005 36301
rect 20947 36292 20959 36295
rect 16209 36255 16267 36261
rect 17236 36264 17908 36292
rect 6089 36227 6147 36233
rect 6089 36193 6101 36227
rect 6135 36224 6147 36227
rect 10413 36227 10471 36233
rect 10413 36224 10425 36227
rect 6135 36196 6960 36224
rect 6135 36193 6147 36196
rect 6089 36187 6147 36193
rect 6932 36168 6960 36196
rect 7024 36196 10425 36224
rect 4065 36159 4123 36165
rect 4065 36125 4077 36159
rect 4111 36156 4123 36159
rect 4614 36156 4620 36168
rect 4111 36128 4620 36156
rect 4111 36125 4123 36128
rect 4065 36119 4123 36125
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 6181 36159 6239 36165
rect 6181 36125 6193 36159
rect 6227 36125 6239 36159
rect 6181 36119 6239 36125
rect 4332 36091 4390 36097
rect 4332 36057 4344 36091
rect 4378 36088 4390 36091
rect 4982 36088 4988 36100
rect 4378 36060 4988 36088
rect 4378 36057 4390 36060
rect 4332 36051 4390 36057
rect 4982 36048 4988 36060
rect 5040 36048 5046 36100
rect 6196 36088 6224 36119
rect 6822 36116 6828 36168
rect 6880 36116 6886 36168
rect 6914 36116 6920 36168
rect 6972 36116 6978 36168
rect 7024 36165 7052 36196
rect 10413 36193 10425 36196
rect 10459 36193 10471 36227
rect 10520 36224 10548 36252
rect 14461 36227 14519 36233
rect 14461 36224 14473 36227
rect 10520 36196 11744 36224
rect 10413 36187 10471 36193
rect 7009 36159 7067 36165
rect 7009 36125 7021 36159
rect 7055 36125 7067 36159
rect 7009 36119 7067 36125
rect 7190 36116 7196 36168
rect 7248 36116 7254 36168
rect 8110 36116 8116 36168
rect 8168 36156 8174 36168
rect 8297 36159 8355 36165
rect 8297 36156 8309 36159
rect 8168 36128 8309 36156
rect 8168 36116 8174 36128
rect 8297 36125 8309 36128
rect 8343 36125 8355 36159
rect 8297 36119 8355 36125
rect 8573 36159 8631 36165
rect 8573 36125 8585 36159
rect 8619 36156 8631 36159
rect 9766 36156 9772 36168
rect 8619 36128 9772 36156
rect 8619 36125 8631 36128
rect 8573 36119 8631 36125
rect 9766 36116 9772 36128
rect 9824 36116 9830 36168
rect 9861 36159 9919 36165
rect 9861 36125 9873 36159
rect 9907 36125 9919 36159
rect 9861 36119 9919 36125
rect 7558 36088 7564 36100
rect 6196 36060 7564 36088
rect 7558 36048 7564 36060
rect 7616 36048 7622 36100
rect 8846 36048 8852 36100
rect 8904 36088 8910 36100
rect 9585 36091 9643 36097
rect 9585 36088 9597 36091
rect 8904 36060 9597 36088
rect 8904 36048 8910 36060
rect 9585 36057 9597 36060
rect 9631 36057 9643 36091
rect 9585 36051 9643 36057
rect 5445 36023 5503 36029
rect 5445 35989 5457 36023
rect 5491 36020 5503 36023
rect 5534 36020 5540 36032
rect 5491 35992 5540 36020
rect 5491 35989 5503 35992
rect 5445 35983 5503 35989
rect 5534 35980 5540 35992
rect 5592 35980 5598 36032
rect 6638 35980 6644 36032
rect 6696 35980 6702 36032
rect 8294 35980 8300 36032
rect 8352 36020 8358 36032
rect 8481 36023 8539 36029
rect 8481 36020 8493 36023
rect 8352 35992 8493 36020
rect 8352 35980 8358 35992
rect 8481 35989 8493 35992
rect 8527 36020 8539 36023
rect 8570 36020 8576 36032
rect 8527 35992 8576 36020
rect 8527 35989 8539 35992
rect 8481 35983 8539 35989
rect 8570 35980 8576 35992
rect 8628 35980 8634 36032
rect 9876 36020 9904 36119
rect 10318 36116 10324 36168
rect 10376 36116 10382 36168
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36125 10563 36159
rect 10505 36119 10563 36125
rect 10520 36088 10548 36119
rect 11054 36116 11060 36168
rect 11112 36116 11118 36168
rect 11330 36116 11336 36168
rect 11388 36116 11394 36168
rect 11514 36116 11520 36168
rect 11572 36116 11578 36168
rect 11716 36165 11744 36196
rect 13556 36196 14473 36224
rect 11701 36159 11759 36165
rect 11701 36125 11713 36159
rect 11747 36156 11759 36159
rect 11882 36156 11888 36168
rect 11747 36128 11888 36156
rect 11747 36125 11759 36128
rect 11701 36119 11759 36125
rect 11882 36116 11888 36128
rect 11940 36116 11946 36168
rect 12526 36116 12532 36168
rect 12584 36116 12590 36168
rect 12621 36159 12679 36165
rect 12621 36125 12633 36159
rect 12667 36156 12679 36159
rect 12894 36156 12900 36168
rect 12667 36128 12900 36156
rect 12667 36125 12679 36128
rect 12621 36119 12679 36125
rect 12894 36116 12900 36128
rect 12952 36116 12958 36168
rect 13078 36116 13084 36168
rect 13136 36156 13142 36168
rect 13556 36165 13584 36196
rect 14461 36193 14473 36196
rect 14507 36224 14519 36227
rect 14642 36224 14648 36236
rect 14507 36196 14648 36224
rect 14507 36193 14519 36196
rect 14461 36187 14519 36193
rect 14642 36184 14648 36196
rect 14700 36184 14706 36236
rect 15672 36224 15700 36252
rect 17236 36224 17264 36264
rect 15672 36196 17264 36224
rect 17310 36184 17316 36236
rect 17368 36184 17374 36236
rect 13541 36159 13599 36165
rect 13541 36156 13553 36159
rect 13136 36128 13553 36156
rect 13136 36116 13142 36128
rect 13541 36125 13553 36128
rect 13587 36125 13599 36159
rect 13541 36119 13599 36125
rect 14182 36116 14188 36168
rect 14240 36156 14246 36168
rect 14553 36159 14611 36165
rect 14553 36156 14565 36159
rect 14240 36128 14565 36156
rect 14240 36116 14246 36128
rect 14553 36125 14565 36128
rect 14599 36125 14611 36159
rect 15102 36156 15108 36168
rect 14553 36119 14611 36125
rect 14660 36128 15108 36156
rect 11974 36088 11980 36100
rect 10520 36060 11980 36088
rect 11974 36048 11980 36060
rect 12032 36088 12038 36100
rect 12345 36091 12403 36097
rect 12345 36088 12357 36091
rect 12032 36060 12357 36088
rect 12032 36048 12038 36060
rect 12345 36057 12357 36060
rect 12391 36088 12403 36091
rect 13357 36091 13415 36097
rect 13357 36088 13369 36091
rect 12391 36060 13369 36088
rect 12391 36057 12403 36060
rect 12345 36051 12403 36057
rect 13357 36057 13369 36060
rect 13403 36057 13415 36091
rect 13357 36051 13415 36057
rect 14277 36091 14335 36097
rect 14277 36057 14289 36091
rect 14323 36088 14335 36091
rect 14660 36088 14688 36128
rect 15102 36116 15108 36128
rect 15160 36116 15166 36168
rect 16942 36116 16948 36168
rect 17000 36156 17006 36168
rect 17037 36159 17095 36165
rect 17037 36156 17049 36159
rect 17000 36128 17049 36156
rect 17000 36116 17006 36128
rect 17037 36125 17049 36128
rect 17083 36156 17095 36159
rect 17678 36156 17684 36168
rect 17083 36128 17684 36156
rect 17083 36125 17095 36128
rect 17037 36119 17095 36125
rect 17678 36116 17684 36128
rect 17736 36116 17742 36168
rect 17773 36159 17831 36165
rect 17773 36125 17785 36159
rect 17819 36125 17831 36159
rect 17773 36119 17831 36125
rect 14323 36060 14688 36088
rect 14323 36057 14335 36060
rect 14277 36051 14335 36057
rect 15010 36048 15016 36100
rect 15068 36088 15074 36100
rect 16025 36091 16083 36097
rect 16025 36088 16037 36091
rect 15068 36060 16037 36088
rect 15068 36048 15074 36060
rect 16025 36057 16037 36060
rect 16071 36088 16083 36091
rect 17788 36088 17816 36119
rect 16071 36060 17816 36088
rect 17880 36088 17908 36264
rect 18524 36264 20959 36292
rect 18524 36168 18552 36264
rect 20947 36261 20959 36264
rect 20993 36292 21005 36295
rect 22094 36292 22100 36304
rect 20993 36264 22100 36292
rect 20993 36261 21005 36264
rect 20947 36255 21005 36261
rect 22094 36252 22100 36264
rect 22152 36252 22158 36304
rect 23382 36252 23388 36304
rect 23440 36292 23446 36304
rect 24596 36292 24624 36332
rect 24946 36292 24952 36304
rect 23440 36264 24624 36292
rect 24688 36264 24952 36292
rect 23440 36252 23446 36264
rect 21821 36227 21879 36233
rect 21821 36224 21833 36227
rect 19720 36196 21833 36224
rect 17954 36116 17960 36168
rect 18012 36116 18018 36168
rect 18506 36116 18512 36168
rect 18564 36116 18570 36168
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36156 18751 36159
rect 19058 36156 19064 36168
rect 18739 36128 19064 36156
rect 18739 36125 18751 36128
rect 18693 36119 18751 36125
rect 19058 36116 19064 36128
rect 19116 36116 19122 36168
rect 19426 36116 19432 36168
rect 19484 36116 19490 36168
rect 19720 36165 19748 36196
rect 21821 36193 21833 36196
rect 21867 36224 21879 36227
rect 21867 36196 22600 36224
rect 21867 36193 21879 36196
rect 21821 36187 21879 36193
rect 19705 36159 19763 36165
rect 19705 36125 19717 36159
rect 19751 36125 19763 36159
rect 19705 36119 19763 36125
rect 19797 36159 19855 36165
rect 19797 36125 19809 36159
rect 19843 36125 19855 36159
rect 19797 36119 19855 36125
rect 19613 36091 19671 36097
rect 19613 36088 19625 36091
rect 17880 36060 19625 36088
rect 16071 36057 16083 36060
rect 16025 36051 16083 36057
rect 19613 36057 19625 36060
rect 19659 36057 19671 36091
rect 19613 36051 19671 36057
rect 10502 36020 10508 36032
rect 9876 35992 10508 36020
rect 10502 35980 10508 35992
rect 10560 35980 10566 36032
rect 11238 35980 11244 36032
rect 11296 35980 11302 36032
rect 11514 35980 11520 36032
rect 11572 36020 11578 36032
rect 12710 36020 12716 36032
rect 11572 35992 12716 36020
rect 11572 35980 11578 35992
rect 12710 35980 12716 35992
rect 12768 35980 12774 36032
rect 12805 36023 12863 36029
rect 12805 35989 12817 36023
rect 12851 36020 12863 36023
rect 17126 36020 17132 36032
rect 12851 35992 17132 36020
rect 12851 35989 12863 35992
rect 12805 35983 12863 35989
rect 17126 35980 17132 35992
rect 17184 35980 17190 36032
rect 18877 36023 18935 36029
rect 18877 35989 18889 36023
rect 18923 36020 18935 36023
rect 19812 36020 19840 36119
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20806 36156 20812 36168
rect 19944 36128 20812 36156
rect 19944 36116 19950 36128
rect 20806 36116 20812 36128
rect 20864 36116 20870 36168
rect 21082 36116 21088 36168
rect 21140 36116 21146 36168
rect 21266 36116 21272 36168
rect 21324 36116 21330 36168
rect 21729 36159 21787 36165
rect 21729 36125 21741 36159
rect 21775 36125 21787 36159
rect 21729 36119 21787 36125
rect 21913 36159 21971 36165
rect 21913 36125 21925 36159
rect 21959 36156 21971 36159
rect 22094 36156 22100 36168
rect 21959 36128 22100 36156
rect 21959 36125 21971 36128
rect 21913 36119 21971 36125
rect 21744 36088 21772 36119
rect 22094 36116 22100 36128
rect 22152 36116 22158 36168
rect 22462 36156 22468 36168
rect 22204 36128 22468 36156
rect 22204 36088 22232 36128
rect 22462 36116 22468 36128
rect 22520 36116 22526 36168
rect 22572 36165 22600 36196
rect 24486 36184 24492 36236
rect 24544 36224 24550 36236
rect 24581 36227 24639 36233
rect 24581 36224 24593 36227
rect 24544 36196 24593 36224
rect 24544 36184 24550 36196
rect 24581 36193 24593 36196
rect 24627 36193 24639 36227
rect 24581 36187 24639 36193
rect 22557 36159 22615 36165
rect 22557 36125 22569 36159
rect 22603 36125 22615 36159
rect 23658 36156 23664 36168
rect 22557 36119 22615 36125
rect 23308 36128 23664 36156
rect 21744 36060 22232 36088
rect 22278 36048 22284 36100
rect 22336 36088 22342 36100
rect 22373 36091 22431 36097
rect 22373 36088 22385 36091
rect 22336 36060 22385 36088
rect 22336 36048 22342 36060
rect 22373 36057 22385 36060
rect 22419 36057 22431 36091
rect 23308 36088 23336 36128
rect 23658 36116 23664 36128
rect 23716 36116 23722 36168
rect 23753 36159 23811 36165
rect 23753 36125 23765 36159
rect 23799 36156 23811 36159
rect 24688 36156 24716 36264
rect 24946 36252 24952 36264
rect 25004 36252 25010 36304
rect 25056 36292 25084 36332
rect 27522 36320 27528 36372
rect 27580 36320 27586 36372
rect 28626 36320 28632 36372
rect 28684 36320 28690 36372
rect 30006 36360 30012 36372
rect 28736 36332 30012 36360
rect 28736 36292 28764 36332
rect 30006 36320 30012 36332
rect 30064 36320 30070 36372
rect 30282 36320 30288 36372
rect 30340 36369 30346 36372
rect 30340 36363 30362 36369
rect 30350 36329 30362 36363
rect 30340 36323 30362 36329
rect 30340 36320 30346 36323
rect 37366 36320 37372 36372
rect 37424 36320 37430 36372
rect 37476 36332 38884 36360
rect 25056 36264 28764 36292
rect 29362 36252 29368 36304
rect 29420 36292 29426 36304
rect 29914 36292 29920 36304
rect 29420 36264 29920 36292
rect 29420 36252 29426 36264
rect 29914 36252 29920 36264
rect 29972 36292 29978 36304
rect 30193 36295 30251 36301
rect 30193 36292 30205 36295
rect 29972 36264 30205 36292
rect 29972 36252 29978 36264
rect 30193 36261 30205 36264
rect 30239 36261 30251 36295
rect 32674 36292 32680 36304
rect 30193 36255 30251 36261
rect 30300 36264 32680 36292
rect 26878 36224 26884 36236
rect 23799 36128 24716 36156
rect 24780 36196 26884 36224
rect 23799 36125 23811 36128
rect 23753 36119 23811 36125
rect 22373 36051 22431 36057
rect 22572 36060 23336 36088
rect 18923 35992 19840 36020
rect 18923 35989 18935 35992
rect 18877 35983 18935 35989
rect 21910 35980 21916 36032
rect 21968 36020 21974 36032
rect 22572 36020 22600 36060
rect 23474 36048 23480 36100
rect 23532 36048 23538 36100
rect 21968 35992 22600 36020
rect 22649 36023 22707 36029
rect 21968 35980 21974 35992
rect 22649 35989 22661 36023
rect 22695 36020 22707 36023
rect 24780 36020 24808 36196
rect 26878 36184 26884 36196
rect 26936 36184 26942 36236
rect 27154 36184 27160 36236
rect 27212 36224 27218 36236
rect 27890 36224 27896 36236
rect 27212 36196 27896 36224
rect 27212 36184 27218 36196
rect 27890 36184 27896 36196
rect 27948 36184 27954 36236
rect 28074 36184 28080 36236
rect 28132 36224 28138 36236
rect 30101 36227 30159 36233
rect 30101 36224 30113 36227
rect 28132 36196 30113 36224
rect 28132 36184 28138 36196
rect 30101 36193 30113 36196
rect 30147 36224 30159 36227
rect 30300 36224 30328 36264
rect 32674 36252 32680 36264
rect 32732 36252 32738 36304
rect 33226 36252 33232 36304
rect 33284 36252 33290 36304
rect 34885 36295 34943 36301
rect 34885 36261 34897 36295
rect 34931 36292 34943 36295
rect 35710 36292 35716 36304
rect 34931 36264 35716 36292
rect 34931 36261 34943 36264
rect 34885 36255 34943 36261
rect 35710 36252 35716 36264
rect 35768 36252 35774 36304
rect 37476 36292 37504 36332
rect 37108 36264 37504 36292
rect 38105 36295 38163 36301
rect 30147 36196 30328 36224
rect 30147 36193 30159 36196
rect 30101 36187 30159 36193
rect 31018 36184 31024 36236
rect 31076 36224 31082 36236
rect 31849 36227 31907 36233
rect 31849 36224 31861 36227
rect 31076 36196 31861 36224
rect 31076 36184 31082 36196
rect 31849 36193 31861 36196
rect 31895 36193 31907 36227
rect 31849 36187 31907 36193
rect 31938 36184 31944 36236
rect 31996 36224 32002 36236
rect 34790 36224 34796 36236
rect 31996 36196 32996 36224
rect 31996 36184 32002 36196
rect 32968 36168 32996 36196
rect 34256 36196 34796 36224
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36125 24915 36159
rect 24857 36119 24915 36125
rect 24949 36159 25007 36165
rect 24949 36125 24961 36159
rect 24995 36125 25007 36159
rect 24949 36119 25007 36125
rect 22695 35992 24808 36020
rect 24872 36020 24900 36119
rect 24964 36088 24992 36119
rect 25038 36116 25044 36168
rect 25096 36116 25102 36168
rect 25225 36159 25283 36165
rect 25225 36125 25237 36159
rect 25271 36156 25283 36159
rect 26510 36156 26516 36168
rect 25271 36128 26516 36156
rect 25271 36125 25283 36128
rect 25225 36119 25283 36125
rect 26510 36116 26516 36128
rect 26568 36116 26574 36168
rect 27706 36116 27712 36168
rect 27764 36116 27770 36168
rect 27801 36159 27859 36165
rect 27801 36125 27813 36159
rect 27847 36125 27859 36159
rect 27801 36119 27859 36125
rect 27985 36159 28043 36165
rect 27985 36125 27997 36159
rect 28031 36156 28043 36159
rect 28442 36156 28448 36168
rect 28031 36128 28448 36156
rect 28031 36125 28043 36128
rect 27985 36119 28043 36125
rect 26528 36088 26556 36116
rect 24964 36060 25452 36088
rect 26528 36060 27568 36088
rect 25424 36032 25452 36060
rect 25130 36020 25136 36032
rect 24872 35992 25136 36020
rect 22695 35989 22707 35992
rect 22649 35983 22707 35989
rect 25130 35980 25136 35992
rect 25188 35980 25194 36032
rect 25406 35980 25412 36032
rect 25464 36020 25470 36032
rect 27430 36020 27436 36032
rect 25464 35992 27436 36020
rect 25464 35980 25470 35992
rect 27430 35980 27436 35992
rect 27488 35980 27494 36032
rect 27540 36020 27568 36060
rect 27614 36048 27620 36100
rect 27672 36088 27678 36100
rect 27816 36088 27844 36119
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 28537 36159 28595 36165
rect 28537 36125 28549 36159
rect 28583 36156 28595 36159
rect 28810 36156 28816 36168
rect 28583 36128 28816 36156
rect 28583 36125 28595 36128
rect 28537 36119 28595 36125
rect 27672 36060 27844 36088
rect 27672 36048 27678 36060
rect 27890 36048 27896 36100
rect 27948 36088 27954 36100
rect 28552 36088 28580 36119
rect 28810 36116 28816 36128
rect 28868 36116 28874 36168
rect 28902 36116 28908 36168
rect 28960 36116 28966 36168
rect 28997 36159 29055 36165
rect 28997 36125 29009 36159
rect 29043 36156 29055 36159
rect 30282 36156 30288 36168
rect 29043 36128 30288 36156
rect 29043 36125 29055 36128
rect 28997 36119 29055 36125
rect 30282 36116 30288 36128
rect 30340 36116 30346 36168
rect 30374 36116 30380 36168
rect 30432 36156 30438 36168
rect 30469 36159 30527 36165
rect 30469 36156 30481 36159
rect 30432 36128 30481 36156
rect 30432 36116 30438 36128
rect 30469 36125 30481 36128
rect 30515 36156 30527 36159
rect 30558 36156 30564 36168
rect 30515 36128 30564 36156
rect 30515 36125 30527 36128
rect 30469 36119 30527 36125
rect 30558 36116 30564 36128
rect 30616 36116 30622 36168
rect 31662 36116 31668 36168
rect 31720 36156 31726 36168
rect 31757 36159 31815 36165
rect 31757 36156 31769 36159
rect 31720 36128 31769 36156
rect 31720 36116 31726 36128
rect 31757 36125 31769 36128
rect 31803 36125 31815 36159
rect 31757 36119 31815 36125
rect 32033 36159 32091 36165
rect 32033 36125 32045 36159
rect 32079 36156 32091 36159
rect 32122 36156 32128 36168
rect 32079 36128 32128 36156
rect 32079 36125 32091 36128
rect 32033 36119 32091 36125
rect 32122 36116 32128 36128
rect 32180 36156 32186 36168
rect 32582 36156 32588 36168
rect 32180 36128 32588 36156
rect 32180 36116 32186 36128
rect 32582 36116 32588 36128
rect 32640 36116 32646 36168
rect 32950 36116 32956 36168
rect 33008 36116 33014 36168
rect 33134 36116 33140 36168
rect 33192 36156 33198 36168
rect 34054 36156 34060 36168
rect 33192 36128 34060 36156
rect 33192 36116 33198 36128
rect 34054 36116 34060 36128
rect 34112 36116 34118 36168
rect 34256 36165 34284 36196
rect 34790 36184 34796 36196
rect 34848 36224 34854 36236
rect 34848 36196 35006 36224
rect 34848 36184 34854 36196
rect 36170 36184 36176 36236
rect 36228 36224 36234 36236
rect 37108 36224 37136 36264
rect 38105 36261 38117 36295
rect 38151 36261 38163 36295
rect 38105 36255 38163 36261
rect 36228 36196 37136 36224
rect 36228 36184 36234 36196
rect 34241 36159 34299 36165
rect 34241 36125 34253 36159
rect 34287 36125 34299 36159
rect 34241 36119 34299 36125
rect 35066 36116 35072 36168
rect 35124 36116 35130 36168
rect 35621 36159 35679 36165
rect 35621 36125 35633 36159
rect 35667 36125 35679 36159
rect 35621 36119 35679 36125
rect 35713 36159 35771 36165
rect 35713 36125 35725 36159
rect 35759 36125 35771 36159
rect 35713 36119 35771 36125
rect 30742 36088 30748 36100
rect 27948 36060 28580 36088
rect 29104 36060 30748 36088
rect 27948 36048 27954 36060
rect 29104 36020 29132 36060
rect 30742 36048 30748 36060
rect 30800 36048 30806 36100
rect 32493 36091 32551 36097
rect 32493 36057 32505 36091
rect 32539 36088 32551 36091
rect 33229 36091 33287 36097
rect 32539 36060 33180 36088
rect 32539 36057 32551 36060
rect 32493 36051 32551 36057
rect 27540 35992 29132 36020
rect 29178 35980 29184 36032
rect 29236 35980 29242 36032
rect 32766 35980 32772 36032
rect 32824 36020 32830 36032
rect 33045 36023 33103 36029
rect 33045 36020 33057 36023
rect 32824 35992 33057 36020
rect 32824 35980 32830 35992
rect 33045 35989 33057 35992
rect 33091 35989 33103 36023
rect 33152 36020 33180 36060
rect 33229 36057 33241 36091
rect 33275 36088 33287 36091
rect 33318 36088 33324 36100
rect 33275 36060 33324 36088
rect 33275 36057 33287 36060
rect 33229 36051 33287 36057
rect 33318 36048 33324 36060
rect 33376 36048 33382 36100
rect 33410 36048 33416 36100
rect 33468 36048 33474 36100
rect 34072 36088 34100 36116
rect 35636 36088 35664 36119
rect 34072 36060 35664 36088
rect 33428 36020 33456 36048
rect 33152 35992 33456 36020
rect 33045 35983 33103 35989
rect 33686 35980 33692 36032
rect 33744 36020 33750 36032
rect 34149 36023 34207 36029
rect 34149 36020 34161 36023
rect 33744 35992 34161 36020
rect 33744 35980 33750 35992
rect 34149 35989 34161 35992
rect 34195 35989 34207 36023
rect 34149 35983 34207 35989
rect 34514 35980 34520 36032
rect 34572 36020 34578 36032
rect 35728 36020 35756 36119
rect 36078 36116 36084 36168
rect 36136 36156 36142 36168
rect 36630 36156 36636 36168
rect 36136 36128 36636 36156
rect 36136 36116 36142 36128
rect 36630 36116 36636 36128
rect 36688 36156 36694 36168
rect 36906 36165 36912 36168
rect 36725 36159 36783 36165
rect 36725 36156 36737 36159
rect 36688 36128 36737 36156
rect 36688 36116 36694 36128
rect 36725 36125 36737 36128
rect 36771 36125 36783 36159
rect 36725 36119 36783 36125
rect 36873 36159 36912 36165
rect 36873 36125 36885 36159
rect 36873 36119 36912 36125
rect 36906 36116 36912 36119
rect 36964 36116 36970 36168
rect 37108 36165 37136 36196
rect 37093 36159 37151 36165
rect 37093 36125 37105 36159
rect 37139 36125 37151 36159
rect 37093 36119 37151 36125
rect 37190 36159 37248 36165
rect 37190 36125 37202 36159
rect 37236 36125 37248 36159
rect 37190 36119 37248 36125
rect 37829 36159 37887 36165
rect 37829 36125 37841 36159
rect 37875 36156 37887 36159
rect 38010 36156 38016 36168
rect 37875 36128 38016 36156
rect 37875 36125 37887 36128
rect 37829 36119 37887 36125
rect 36354 36048 36360 36100
rect 36412 36088 36418 36100
rect 36998 36088 37004 36100
rect 36412 36060 37004 36088
rect 36412 36048 36418 36060
rect 36998 36048 37004 36060
rect 37056 36048 37062 36100
rect 34572 35992 35756 36020
rect 34572 35980 34578 35992
rect 35986 35980 35992 36032
rect 36044 36020 36050 36032
rect 36446 36020 36452 36032
rect 36044 35992 36452 36020
rect 36044 35980 36050 35992
rect 36446 35980 36452 35992
rect 36504 36020 36510 36032
rect 37200 36020 37228 36119
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 38120 36156 38148 36255
rect 38565 36159 38623 36165
rect 38565 36156 38577 36159
rect 38120 36128 38577 36156
rect 38565 36125 38577 36128
rect 38611 36125 38623 36159
rect 38565 36119 38623 36125
rect 38746 36116 38752 36168
rect 38804 36116 38810 36168
rect 38856 36156 38884 36332
rect 39758 36184 39764 36236
rect 39816 36224 39822 36236
rect 39816 36196 40540 36224
rect 39816 36184 39822 36196
rect 40037 36159 40095 36165
rect 40037 36156 40049 36159
rect 38856 36128 40049 36156
rect 40037 36125 40049 36128
rect 40083 36125 40095 36159
rect 40405 36159 40463 36165
rect 40405 36156 40417 36159
rect 40037 36119 40095 36125
rect 40144 36128 40417 36156
rect 38105 36091 38163 36097
rect 38105 36057 38117 36091
rect 38151 36057 38163 36091
rect 38105 36051 38163 36057
rect 36504 35992 37228 36020
rect 36504 35980 36510 35992
rect 37918 35980 37924 36032
rect 37976 35980 37982 36032
rect 38010 35980 38016 36032
rect 38068 36020 38074 36032
rect 38120 36020 38148 36051
rect 39390 36048 39396 36100
rect 39448 36088 39454 36100
rect 40144 36088 40172 36128
rect 40405 36125 40417 36128
rect 40451 36125 40463 36159
rect 40405 36119 40463 36125
rect 39448 36060 40172 36088
rect 40221 36091 40279 36097
rect 39448 36048 39454 36060
rect 40221 36057 40233 36091
rect 40267 36057 40279 36091
rect 40221 36051 40279 36057
rect 40313 36091 40371 36097
rect 40313 36057 40325 36091
rect 40359 36088 40371 36091
rect 40512 36088 40540 36196
rect 41874 36116 41880 36168
rect 41932 36116 41938 36168
rect 40359 36060 40540 36088
rect 42144 36091 42202 36097
rect 40359 36057 40371 36060
rect 40313 36051 40371 36057
rect 42144 36057 42156 36091
rect 42190 36088 42202 36091
rect 42610 36088 42616 36100
rect 42190 36060 42616 36088
rect 42190 36057 42202 36060
rect 42144 36051 42202 36057
rect 38068 35992 38148 36020
rect 38657 36023 38715 36029
rect 38068 35980 38074 35992
rect 38657 35989 38669 36023
rect 38703 36020 38715 36023
rect 39114 36020 39120 36032
rect 38703 35992 39120 36020
rect 38703 35989 38715 35992
rect 38657 35983 38715 35989
rect 39114 35980 39120 35992
rect 39172 35980 39178 36032
rect 39298 35980 39304 36032
rect 39356 36020 39362 36032
rect 39942 36020 39948 36032
rect 39356 35992 39948 36020
rect 39356 35980 39362 35992
rect 39942 35980 39948 35992
rect 40000 36020 40006 36032
rect 40236 36020 40264 36051
rect 42610 36048 42616 36060
rect 42668 36048 42674 36100
rect 40000 35992 40264 36020
rect 40589 36023 40647 36029
rect 40000 35980 40006 35992
rect 40589 35989 40601 36023
rect 40635 36020 40647 36023
rect 40954 36020 40960 36032
rect 40635 35992 40960 36020
rect 40635 35989 40647 35992
rect 40589 35983 40647 35989
rect 40954 35980 40960 35992
rect 41012 35980 41018 36032
rect 43254 35980 43260 36032
rect 43312 35980 43318 36032
rect 1104 35930 43884 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 43884 35930
rect 1104 35856 43884 35878
rect 4982 35776 4988 35828
rect 5040 35776 5046 35828
rect 6822 35776 6828 35828
rect 6880 35816 6886 35828
rect 8202 35816 8208 35828
rect 6880 35788 8208 35816
rect 6880 35776 6886 35788
rect 7190 35708 7196 35760
rect 7248 35748 7254 35760
rect 7484 35757 7512 35788
rect 8202 35776 8208 35788
rect 8260 35776 8266 35828
rect 8297 35819 8355 35825
rect 8297 35785 8309 35819
rect 8343 35816 8355 35819
rect 8938 35816 8944 35828
rect 8343 35788 8944 35816
rect 8343 35785 8355 35788
rect 8297 35779 8355 35785
rect 7377 35751 7435 35757
rect 7377 35748 7389 35751
rect 7248 35720 7389 35748
rect 7248 35708 7254 35720
rect 7377 35717 7389 35720
rect 7423 35717 7435 35751
rect 7377 35711 7435 35717
rect 7469 35751 7527 35757
rect 7469 35717 7481 35751
rect 7515 35717 7527 35751
rect 8312 35748 8340 35779
rect 8938 35776 8944 35788
rect 8996 35776 9002 35828
rect 9766 35776 9772 35828
rect 9824 35816 9830 35828
rect 10318 35816 10324 35828
rect 9824 35788 10324 35816
rect 9824 35776 9830 35788
rect 10318 35776 10324 35788
rect 10376 35776 10382 35828
rect 11974 35776 11980 35828
rect 12032 35816 12038 35828
rect 12069 35819 12127 35825
rect 12069 35816 12081 35819
rect 12032 35788 12081 35816
rect 12032 35776 12038 35788
rect 12069 35785 12081 35788
rect 12115 35816 12127 35819
rect 12115 35788 12434 35816
rect 12115 35785 12127 35788
rect 12069 35779 12127 35785
rect 10042 35748 10048 35760
rect 7469 35711 7527 35717
rect 7668 35720 8340 35748
rect 9232 35720 10048 35748
rect 7668 35689 7696 35720
rect 9232 35692 9260 35720
rect 10042 35708 10048 35720
rect 10100 35708 10106 35760
rect 11882 35708 11888 35760
rect 11940 35708 11946 35760
rect 7285 35683 7343 35689
rect 7285 35649 7297 35683
rect 7331 35649 7343 35683
rect 7285 35643 7343 35649
rect 7653 35683 7711 35689
rect 7653 35649 7665 35683
rect 7699 35649 7711 35683
rect 7653 35643 7711 35649
rect 5166 35572 5172 35624
rect 5224 35572 5230 35624
rect 5261 35615 5319 35621
rect 5261 35581 5273 35615
rect 5307 35581 5319 35615
rect 5261 35575 5319 35581
rect 5276 35544 5304 35575
rect 5350 35572 5356 35624
rect 5408 35572 5414 35624
rect 5442 35572 5448 35624
rect 5500 35572 5506 35624
rect 7300 35612 7328 35643
rect 7834 35640 7840 35692
rect 7892 35680 7898 35692
rect 8205 35683 8263 35689
rect 8205 35680 8217 35683
rect 7892 35652 8217 35680
rect 7892 35640 7898 35652
rect 8205 35649 8217 35652
rect 8251 35649 8263 35683
rect 8205 35643 8263 35649
rect 8389 35683 8447 35689
rect 8389 35649 8401 35683
rect 8435 35680 8447 35683
rect 8754 35680 8760 35692
rect 8435 35652 8760 35680
rect 8435 35649 8447 35652
rect 8389 35643 8447 35649
rect 8754 35640 8760 35652
rect 8812 35640 8818 35692
rect 8846 35640 8852 35692
rect 8904 35680 8910 35692
rect 8941 35683 8999 35689
rect 8941 35680 8953 35683
rect 8904 35652 8953 35680
rect 8904 35640 8910 35652
rect 8941 35649 8953 35652
rect 8987 35649 8999 35683
rect 8941 35643 8999 35649
rect 9214 35640 9220 35692
rect 9272 35640 9278 35692
rect 9674 35640 9680 35692
rect 9732 35680 9738 35692
rect 9950 35680 9956 35692
rect 9732 35652 9956 35680
rect 9732 35640 9738 35652
rect 9950 35640 9956 35652
rect 10008 35640 10014 35692
rect 10134 35640 10140 35692
rect 10192 35680 10198 35692
rect 10594 35680 10600 35692
rect 10192 35652 10600 35680
rect 10192 35640 10198 35652
rect 10594 35640 10600 35652
rect 10652 35640 10658 35692
rect 11606 35640 11612 35692
rect 11664 35680 11670 35692
rect 11701 35683 11759 35689
rect 11701 35680 11713 35683
rect 11664 35652 11713 35680
rect 11664 35640 11670 35652
rect 11701 35649 11713 35652
rect 11747 35649 11759 35683
rect 12406 35680 12434 35788
rect 12802 35776 12808 35828
rect 12860 35776 12866 35828
rect 13354 35776 13360 35828
rect 13412 35816 13418 35828
rect 15194 35816 15200 35828
rect 13412 35788 15200 35816
rect 13412 35776 13418 35788
rect 15194 35776 15200 35788
rect 15252 35776 15258 35828
rect 15565 35819 15623 35825
rect 15565 35785 15577 35819
rect 15611 35816 15623 35819
rect 16022 35816 16028 35828
rect 15611 35788 16028 35816
rect 15611 35785 15623 35788
rect 15565 35779 15623 35785
rect 16022 35776 16028 35788
rect 16080 35776 16086 35828
rect 19334 35816 19340 35828
rect 16132 35788 19340 35816
rect 12710 35708 12716 35760
rect 12768 35748 12774 35760
rect 13538 35748 13544 35760
rect 12768 35720 13544 35748
rect 12768 35708 12774 35720
rect 13538 35708 13544 35720
rect 13596 35708 13602 35760
rect 14277 35751 14335 35757
rect 14277 35717 14289 35751
rect 14323 35748 14335 35751
rect 14458 35748 14464 35760
rect 14323 35720 14464 35748
rect 14323 35717 14335 35720
rect 14277 35711 14335 35717
rect 14458 35708 14464 35720
rect 14516 35708 14522 35760
rect 16132 35748 16160 35788
rect 17034 35748 17040 35760
rect 14936 35720 16160 35748
rect 16224 35720 17040 35748
rect 12897 35683 12955 35689
rect 12897 35680 12909 35683
rect 12406 35652 12909 35680
rect 11701 35643 11759 35649
rect 12897 35649 12909 35652
rect 12943 35649 12955 35683
rect 12897 35643 12955 35649
rect 12986 35640 12992 35692
rect 13044 35680 13050 35692
rect 13081 35683 13139 35689
rect 13081 35680 13093 35683
rect 13044 35652 13093 35680
rect 13044 35640 13050 35652
rect 13081 35649 13093 35652
rect 13127 35649 13139 35683
rect 13081 35643 13139 35649
rect 14550 35640 14556 35692
rect 14608 35680 14614 35692
rect 14826 35680 14832 35692
rect 14608 35652 14832 35680
rect 14608 35640 14614 35652
rect 14826 35640 14832 35652
rect 14884 35640 14890 35692
rect 7300 35584 8432 35612
rect 8404 35556 8432 35584
rect 14366 35572 14372 35624
rect 14424 35572 14430 35624
rect 14936 35612 14964 35720
rect 15378 35640 15384 35692
rect 15436 35640 15442 35692
rect 15565 35683 15623 35689
rect 15565 35649 15577 35683
rect 15611 35649 15623 35683
rect 15565 35643 15623 35649
rect 14476 35584 14964 35612
rect 15580 35612 15608 35643
rect 15746 35640 15752 35692
rect 15804 35680 15810 35692
rect 16224 35689 16252 35720
rect 17034 35708 17040 35720
rect 17092 35708 17098 35760
rect 16025 35683 16083 35689
rect 16025 35680 16037 35683
rect 15804 35652 16037 35680
rect 15804 35640 15810 35652
rect 16025 35649 16037 35652
rect 16071 35649 16083 35683
rect 16025 35643 16083 35649
rect 16209 35683 16267 35689
rect 16209 35649 16221 35683
rect 16255 35649 16267 35683
rect 16209 35643 16267 35649
rect 16942 35640 16948 35692
rect 17000 35640 17006 35692
rect 17126 35640 17132 35692
rect 17184 35640 17190 35692
rect 17696 35689 17724 35788
rect 19334 35776 19340 35788
rect 19392 35776 19398 35828
rect 19886 35776 19892 35828
rect 19944 35816 19950 35828
rect 20070 35816 20076 35828
rect 19944 35788 20076 35816
rect 19944 35776 19950 35788
rect 20070 35776 20076 35788
rect 20128 35776 20134 35828
rect 20625 35819 20683 35825
rect 20625 35785 20637 35819
rect 20671 35816 20683 35819
rect 20714 35816 20720 35828
rect 20671 35788 20720 35816
rect 20671 35785 20683 35788
rect 20625 35779 20683 35785
rect 20714 35776 20720 35788
rect 20772 35776 20778 35828
rect 21082 35776 21088 35828
rect 21140 35816 21146 35828
rect 22005 35819 22063 35825
rect 22005 35816 22017 35819
rect 21140 35788 22017 35816
rect 21140 35776 21146 35788
rect 22005 35785 22017 35788
rect 22051 35785 22063 35819
rect 22005 35779 22063 35785
rect 23474 35776 23480 35828
rect 23532 35776 23538 35828
rect 23842 35776 23848 35828
rect 23900 35816 23906 35828
rect 24578 35816 24584 35828
rect 23900 35788 24584 35816
rect 23900 35776 23906 35788
rect 24578 35776 24584 35788
rect 24636 35816 24642 35828
rect 24949 35819 25007 35825
rect 24949 35816 24961 35819
rect 24636 35788 24961 35816
rect 24636 35776 24642 35788
rect 24949 35785 24961 35788
rect 24995 35785 25007 35819
rect 27614 35816 27620 35828
rect 24949 35779 25007 35785
rect 27264 35788 27620 35816
rect 17957 35751 18015 35757
rect 17957 35717 17969 35751
rect 18003 35748 18015 35751
rect 18138 35748 18144 35760
rect 18003 35720 18144 35748
rect 18003 35717 18015 35720
rect 17957 35711 18015 35717
rect 18138 35708 18144 35720
rect 18196 35708 18202 35760
rect 18785 35751 18843 35757
rect 18785 35717 18797 35751
rect 18831 35748 18843 35751
rect 20165 35751 20223 35757
rect 20165 35748 20177 35751
rect 18831 35720 20177 35748
rect 18831 35717 18843 35720
rect 18785 35711 18843 35717
rect 20165 35717 20177 35720
rect 20211 35717 20223 35751
rect 25038 35748 25044 35760
rect 20165 35711 20223 35717
rect 22066 35720 25044 35748
rect 17681 35683 17739 35689
rect 17681 35649 17693 35683
rect 17727 35649 17739 35683
rect 17681 35643 17739 35649
rect 17862 35640 17868 35692
rect 17920 35640 17926 35692
rect 18046 35640 18052 35692
rect 18104 35680 18110 35692
rect 18693 35683 18751 35689
rect 18693 35680 18705 35683
rect 18104 35652 18705 35680
rect 18104 35640 18110 35652
rect 18693 35649 18705 35652
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 18874 35640 18880 35692
rect 18932 35640 18938 35692
rect 20441 35683 20499 35689
rect 20441 35649 20453 35683
rect 20487 35680 20499 35683
rect 21266 35680 21272 35692
rect 20487 35652 21272 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 21266 35640 21272 35652
rect 21324 35640 21330 35692
rect 15654 35612 15660 35624
rect 15580 35584 15660 35612
rect 7006 35544 7012 35556
rect 5276 35516 7012 35544
rect 7006 35504 7012 35516
rect 7064 35544 7070 35556
rect 7064 35516 8156 35544
rect 7064 35504 7070 35516
rect 8128 35488 8156 35516
rect 8386 35504 8392 35556
rect 8444 35504 8450 35556
rect 9125 35547 9183 35553
rect 9125 35513 9137 35547
rect 9171 35544 9183 35547
rect 9674 35544 9680 35556
rect 9171 35516 9680 35544
rect 9171 35513 9183 35516
rect 9125 35507 9183 35513
rect 9674 35504 9680 35516
rect 9732 35544 9738 35556
rect 10962 35544 10968 35556
rect 9732 35516 10968 35544
rect 9732 35504 9738 35516
rect 10962 35504 10968 35516
rect 11020 35504 11026 35556
rect 12710 35504 12716 35556
rect 12768 35544 12774 35556
rect 14476 35544 14504 35584
rect 15654 35572 15660 35584
rect 15712 35612 15718 35624
rect 16117 35615 16175 35621
rect 16117 35612 16129 35615
rect 15712 35584 16129 35612
rect 15712 35572 15718 35584
rect 16117 35581 16129 35584
rect 16163 35581 16175 35615
rect 16117 35575 16175 35581
rect 17037 35615 17095 35621
rect 17037 35581 17049 35615
rect 17083 35612 17095 35615
rect 17880 35612 17908 35640
rect 17083 35584 17908 35612
rect 20349 35615 20407 35621
rect 17083 35581 17095 35584
rect 17037 35575 17095 35581
rect 20349 35581 20361 35615
rect 20395 35612 20407 35615
rect 21910 35612 21916 35624
rect 20395 35584 21916 35612
rect 20395 35581 20407 35584
rect 20349 35575 20407 35581
rect 21910 35572 21916 35584
rect 21968 35572 21974 35624
rect 12768 35516 14504 35544
rect 14737 35547 14795 35553
rect 12768 35504 12774 35516
rect 14737 35513 14749 35547
rect 14783 35544 14795 35547
rect 22066 35544 22094 35720
rect 22186 35640 22192 35692
rect 22244 35640 22250 35692
rect 22281 35683 22339 35689
rect 22281 35649 22293 35683
rect 22327 35680 22339 35683
rect 22554 35680 22560 35692
rect 22327 35652 22560 35680
rect 22327 35649 22339 35652
rect 22281 35643 22339 35649
rect 22554 35640 22560 35652
rect 22612 35640 22618 35692
rect 22649 35683 22707 35689
rect 22649 35649 22661 35683
rect 22695 35680 22707 35683
rect 23290 35680 23296 35692
rect 22695 35652 23296 35680
rect 22695 35649 22707 35652
rect 22649 35643 22707 35649
rect 23290 35640 23296 35652
rect 23348 35640 23354 35692
rect 23492 35689 23520 35720
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 25130 35708 25136 35760
rect 25188 35748 25194 35760
rect 25188 35720 25452 35748
rect 25188 35708 25194 35720
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35649 23535 35683
rect 23477 35643 23535 35649
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35680 23719 35683
rect 24026 35680 24032 35692
rect 23707 35652 24032 35680
rect 23707 35649 23719 35652
rect 23661 35643 23719 35649
rect 24026 35640 24032 35652
rect 24084 35640 24090 35692
rect 24210 35640 24216 35692
rect 24268 35640 24274 35692
rect 25424 35689 25452 35720
rect 25409 35683 25467 35689
rect 25409 35649 25421 35683
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 25682 35640 25688 35692
rect 25740 35680 25746 35692
rect 26053 35683 26111 35689
rect 26053 35680 26065 35683
rect 25740 35652 26065 35680
rect 25740 35640 25746 35652
rect 26053 35649 26065 35652
rect 26099 35649 26111 35683
rect 26053 35643 26111 35649
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 27062 35680 27068 35692
rect 26467 35652 27068 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 27062 35640 27068 35652
rect 27120 35640 27126 35692
rect 22373 35615 22431 35621
rect 22373 35581 22385 35615
rect 22419 35581 22431 35615
rect 22373 35575 22431 35581
rect 14783 35516 22094 35544
rect 14783 35513 14795 35516
rect 14737 35507 14795 35513
rect 22186 35504 22192 35556
rect 22244 35544 22250 35556
rect 22388 35544 22416 35575
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 23382 35544 23388 35556
rect 22244 35516 23388 35544
rect 22244 35504 22250 35516
rect 23382 35504 23388 35516
rect 23440 35504 23446 35556
rect 24228 35544 24256 35640
rect 25130 35572 25136 35624
rect 25188 35612 25194 35624
rect 25961 35615 26019 35621
rect 25961 35612 25973 35615
rect 25188 35584 25973 35612
rect 25188 35572 25194 35584
rect 25961 35581 25973 35584
rect 26007 35581 26019 35615
rect 25961 35575 26019 35581
rect 26326 35572 26332 35624
rect 26384 35612 26390 35624
rect 27264 35621 27292 35788
rect 27614 35776 27620 35788
rect 27672 35776 27678 35828
rect 27706 35776 27712 35828
rect 27764 35816 27770 35828
rect 31481 35819 31539 35825
rect 31481 35816 31493 35819
rect 27764 35788 31493 35816
rect 27764 35776 27770 35788
rect 31481 35785 31493 35788
rect 31527 35816 31539 35819
rect 31938 35816 31944 35828
rect 31527 35788 31944 35816
rect 31527 35785 31539 35788
rect 31481 35779 31539 35785
rect 31938 35776 31944 35788
rect 31996 35776 32002 35828
rect 33042 35776 33048 35828
rect 33100 35816 33106 35828
rect 36906 35816 36912 35828
rect 33100 35788 36912 35816
rect 33100 35776 33106 35788
rect 36906 35776 36912 35788
rect 36964 35776 36970 35828
rect 38289 35819 38347 35825
rect 38289 35785 38301 35819
rect 38335 35816 38347 35819
rect 38746 35816 38752 35828
rect 38335 35788 38752 35816
rect 38335 35785 38347 35788
rect 38289 35779 38347 35785
rect 38746 35776 38752 35788
rect 38804 35776 38810 35828
rect 42610 35776 42616 35828
rect 42668 35776 42674 35828
rect 28350 35708 28356 35760
rect 28408 35748 28414 35760
rect 28902 35748 28908 35760
rect 28408 35720 28908 35748
rect 28408 35708 28414 35720
rect 28902 35708 28908 35720
rect 28960 35708 28966 35760
rect 30374 35708 30380 35760
rect 30432 35748 30438 35760
rect 30432 35720 31754 35748
rect 30432 35708 30438 35720
rect 27706 35689 27712 35692
rect 27663 35683 27712 35689
rect 27663 35649 27675 35683
rect 27709 35649 27712 35683
rect 27663 35643 27712 35649
rect 27706 35640 27712 35643
rect 27764 35640 27770 35692
rect 27890 35640 27896 35692
rect 27948 35680 27954 35692
rect 29089 35683 29147 35689
rect 29089 35680 29101 35683
rect 27948 35652 29101 35680
rect 27948 35640 27954 35652
rect 29089 35649 29101 35652
rect 29135 35649 29147 35683
rect 29089 35643 29147 35649
rect 30098 35640 30104 35692
rect 30156 35680 30162 35692
rect 30558 35680 30564 35692
rect 30156 35652 30564 35680
rect 30156 35640 30162 35652
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 31113 35683 31171 35689
rect 31113 35649 31125 35683
rect 31159 35680 31171 35683
rect 31478 35680 31484 35692
rect 31159 35652 31484 35680
rect 31159 35649 31171 35652
rect 31113 35643 31171 35649
rect 27249 35615 27307 35621
rect 27249 35612 27261 35615
rect 26384 35584 27261 35612
rect 26384 35572 26390 35584
rect 27249 35581 27261 35584
rect 27295 35581 27307 35615
rect 27249 35575 27307 35581
rect 27525 35615 27583 35621
rect 27525 35581 27537 35615
rect 27571 35612 27583 35615
rect 28350 35612 28356 35624
rect 27571 35584 28356 35612
rect 27571 35581 27583 35584
rect 27525 35575 27583 35581
rect 28350 35572 28356 35584
rect 28408 35572 28414 35624
rect 30193 35615 30251 35621
rect 30193 35581 30205 35615
rect 30239 35581 30251 35615
rect 30193 35575 30251 35581
rect 25317 35547 25375 35553
rect 24228 35516 25268 35544
rect 7098 35436 7104 35488
rect 7156 35436 7162 35488
rect 8110 35436 8116 35488
rect 8168 35476 8174 35488
rect 10321 35479 10379 35485
rect 10321 35476 10333 35479
rect 8168 35448 10333 35476
rect 8168 35436 8174 35448
rect 10321 35445 10333 35448
rect 10367 35445 10379 35479
rect 10321 35439 10379 35445
rect 14274 35436 14280 35488
rect 14332 35436 14338 35488
rect 18230 35436 18236 35488
rect 18288 35436 18294 35488
rect 20438 35436 20444 35488
rect 20496 35436 20502 35488
rect 22554 35436 22560 35488
rect 22612 35476 22618 35488
rect 24210 35476 24216 35488
rect 22612 35448 24216 35476
rect 22612 35436 22618 35448
rect 24210 35436 24216 35448
rect 24268 35436 24274 35488
rect 24305 35479 24363 35485
rect 24305 35445 24317 35479
rect 24351 35476 24363 35479
rect 24762 35476 24768 35488
rect 24351 35448 24768 35476
rect 24351 35445 24363 35448
rect 24305 35439 24363 35445
rect 24762 35436 24768 35448
rect 24820 35436 24826 35488
rect 25240 35476 25268 35516
rect 25317 35513 25329 35547
rect 25363 35544 25375 35547
rect 25406 35544 25412 35556
rect 25363 35516 25412 35544
rect 25363 35513 25375 35516
rect 25317 35507 25375 35513
rect 25406 35504 25412 35516
rect 25464 35504 25470 35556
rect 26068 35516 27752 35544
rect 26068 35476 26096 35516
rect 25240 35448 26096 35476
rect 26142 35436 26148 35488
rect 26200 35476 26206 35488
rect 26329 35479 26387 35485
rect 26329 35476 26341 35479
rect 26200 35448 26341 35476
rect 26200 35436 26206 35448
rect 26329 35445 26341 35448
rect 26375 35445 26387 35479
rect 26329 35439 26387 35445
rect 26602 35436 26608 35488
rect 26660 35436 26666 35488
rect 27724 35485 27752 35516
rect 27982 35504 27988 35556
rect 28040 35544 28046 35556
rect 28077 35547 28135 35553
rect 28077 35544 28089 35547
rect 28040 35516 28089 35544
rect 28040 35504 28046 35516
rect 28077 35513 28089 35516
rect 28123 35513 28135 35547
rect 30208 35544 30236 35575
rect 30374 35572 30380 35624
rect 30432 35572 30438 35624
rect 30653 35615 30711 35621
rect 30653 35581 30665 35615
rect 30699 35612 30711 35615
rect 30834 35612 30840 35624
rect 30699 35584 30840 35612
rect 30699 35581 30711 35584
rect 30653 35575 30711 35581
rect 30834 35572 30840 35584
rect 30892 35572 30898 35624
rect 30926 35544 30932 35556
rect 30208 35516 30932 35544
rect 28077 35507 28135 35513
rect 30926 35504 30932 35516
rect 30984 35544 30990 35556
rect 31128 35544 31156 35643
rect 31478 35640 31484 35652
rect 31536 35640 31542 35692
rect 31726 35680 31754 35720
rect 32674 35708 32680 35760
rect 32732 35748 32738 35760
rect 36170 35748 36176 35760
rect 32732 35720 36176 35748
rect 32732 35708 32738 35720
rect 36170 35708 36176 35720
rect 36228 35708 36234 35760
rect 37918 35708 37924 35760
rect 37976 35708 37982 35760
rect 38010 35708 38016 35760
rect 38068 35748 38074 35760
rect 38105 35751 38163 35757
rect 38105 35748 38117 35751
rect 38068 35720 38117 35748
rect 38068 35708 38074 35720
rect 38105 35717 38117 35720
rect 38151 35717 38163 35751
rect 41782 35748 41788 35760
rect 38105 35711 38163 35717
rect 39040 35720 41788 35748
rect 33229 35683 33287 35689
rect 33229 35680 33241 35683
rect 31726 35652 33241 35680
rect 33229 35649 33241 35652
rect 33275 35680 33287 35683
rect 33318 35680 33324 35692
rect 33275 35652 33324 35680
rect 33275 35649 33287 35652
rect 33229 35643 33287 35649
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 33410 35640 33416 35692
rect 33468 35640 33474 35692
rect 34149 35683 34207 35689
rect 34149 35649 34161 35683
rect 34195 35680 34207 35683
rect 34238 35680 34244 35692
rect 34195 35652 34244 35680
rect 34195 35649 34207 35652
rect 34149 35643 34207 35649
rect 34238 35640 34244 35652
rect 34296 35640 34302 35692
rect 34330 35640 34336 35692
rect 34388 35640 34394 35692
rect 37936 35680 37964 35708
rect 38378 35680 38384 35692
rect 37936 35652 38384 35680
rect 38378 35640 38384 35652
rect 38436 35640 38442 35692
rect 31202 35572 31208 35624
rect 31260 35612 31266 35624
rect 31754 35612 31760 35624
rect 31260 35584 31760 35612
rect 31260 35572 31266 35584
rect 31754 35572 31760 35584
rect 31812 35612 31818 35624
rect 32030 35612 32036 35624
rect 31812 35584 32036 35612
rect 31812 35572 31818 35584
rect 32030 35572 32036 35584
rect 32088 35572 32094 35624
rect 33134 35572 33140 35624
rect 33192 35572 33198 35624
rect 35618 35572 35624 35624
rect 35676 35612 35682 35624
rect 39040 35621 39068 35720
rect 41782 35708 41788 35720
rect 41840 35708 41846 35760
rect 43254 35708 43260 35760
rect 43312 35708 43318 35760
rect 39114 35640 39120 35692
rect 39172 35680 39178 35692
rect 39281 35683 39339 35689
rect 39281 35680 39293 35683
rect 39172 35652 39293 35680
rect 39172 35640 39178 35652
rect 39281 35649 39293 35652
rect 39327 35649 39339 35683
rect 39281 35643 39339 35649
rect 40954 35640 40960 35692
rect 41012 35640 41018 35692
rect 41050 35683 41108 35689
rect 41050 35649 41062 35683
rect 41096 35649 41108 35683
rect 41050 35643 41108 35649
rect 39025 35615 39083 35621
rect 39025 35612 39037 35615
rect 35676 35584 39037 35612
rect 35676 35572 35682 35584
rect 39025 35581 39037 35584
rect 39071 35581 39083 35615
rect 39025 35575 39083 35581
rect 30984 35516 31156 35544
rect 31312 35516 31754 35544
rect 30984 35504 30990 35516
rect 27709 35479 27767 35485
rect 27709 35445 27721 35479
rect 27755 35445 27767 35479
rect 27709 35439 27767 35445
rect 28994 35436 29000 35488
rect 29052 35476 29058 35488
rect 29365 35479 29423 35485
rect 29365 35476 29377 35479
rect 29052 35448 29377 35476
rect 29052 35436 29058 35448
rect 29365 35445 29377 35448
rect 29411 35476 29423 35479
rect 29638 35476 29644 35488
rect 29411 35448 29644 35476
rect 29411 35445 29423 35448
rect 29365 35439 29423 35445
rect 29638 35436 29644 35448
rect 29696 35436 29702 35488
rect 31312 35485 31340 35516
rect 31297 35479 31355 35485
rect 31297 35445 31309 35479
rect 31343 35445 31355 35479
rect 31726 35476 31754 35516
rect 36906 35504 36912 35556
rect 36964 35544 36970 35556
rect 41064 35544 41092 35643
rect 41230 35640 41236 35692
rect 41288 35640 41294 35692
rect 41322 35640 41328 35692
rect 41380 35640 41386 35692
rect 41422 35683 41480 35689
rect 41422 35649 41434 35683
rect 41468 35649 41480 35683
rect 42981 35683 43039 35689
rect 42981 35680 42993 35683
rect 41422 35643 41480 35649
rect 41524 35652 42993 35680
rect 41432 35612 41460 35643
rect 41386 35584 41460 35612
rect 36964 35516 39068 35544
rect 36964 35504 36970 35516
rect 32122 35476 32128 35488
rect 31726 35448 32128 35476
rect 31297 35439 31355 35445
rect 32122 35436 32128 35448
rect 32180 35436 32186 35488
rect 33594 35436 33600 35488
rect 33652 35476 33658 35488
rect 34241 35479 34299 35485
rect 34241 35476 34253 35479
rect 33652 35448 34253 35476
rect 33652 35436 33658 35448
rect 34241 35445 34253 35448
rect 34287 35445 34299 35479
rect 34241 35439 34299 35445
rect 38102 35436 38108 35488
rect 38160 35436 38166 35488
rect 39040 35476 39068 35516
rect 40236 35516 41092 35544
rect 40236 35476 40264 35516
rect 39040 35448 40264 35476
rect 40310 35436 40316 35488
rect 40368 35476 40374 35488
rect 40405 35479 40463 35485
rect 40405 35476 40417 35479
rect 40368 35448 40417 35476
rect 40368 35436 40374 35448
rect 40405 35445 40417 35448
rect 40451 35445 40463 35479
rect 41064 35476 41092 35516
rect 41138 35504 41144 35556
rect 41196 35544 41202 35556
rect 41386 35544 41414 35584
rect 41196 35516 41414 35544
rect 41196 35504 41202 35516
rect 41524 35476 41552 35652
rect 42981 35649 42993 35652
rect 43027 35680 43039 35683
rect 43272 35680 43300 35708
rect 43027 35652 43300 35680
rect 43027 35649 43039 35652
rect 42981 35643 43039 35649
rect 41966 35612 41972 35624
rect 41616 35584 41972 35612
rect 41616 35553 41644 35584
rect 41966 35572 41972 35584
rect 42024 35612 42030 35624
rect 43073 35615 43131 35621
rect 43073 35612 43085 35615
rect 42024 35584 43085 35612
rect 42024 35572 42030 35584
rect 43073 35581 43085 35584
rect 43119 35581 43131 35615
rect 43073 35575 43131 35581
rect 43254 35572 43260 35624
rect 43312 35572 43318 35624
rect 41601 35547 41659 35553
rect 41601 35513 41613 35547
rect 41647 35513 41659 35547
rect 41601 35507 41659 35513
rect 41064 35448 41552 35476
rect 40405 35439 40463 35445
rect 1104 35386 43884 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 43884 35386
rect 1104 35312 43884 35334
rect 5353 35275 5411 35281
rect 5353 35241 5365 35275
rect 5399 35272 5411 35275
rect 5442 35272 5448 35284
rect 5399 35244 5448 35272
rect 5399 35241 5411 35244
rect 5353 35235 5411 35241
rect 5442 35232 5448 35244
rect 5500 35232 5506 35284
rect 9582 35232 9588 35284
rect 9640 35272 9646 35284
rect 9640 35244 11836 35272
rect 9640 35232 9646 35244
rect 5166 35164 5172 35216
rect 5224 35204 5230 35216
rect 5224 35176 8432 35204
rect 5224 35164 5230 35176
rect 7558 35096 7564 35148
rect 7616 35096 7622 35148
rect 7926 35136 7932 35148
rect 7852 35108 7932 35136
rect 5534 35028 5540 35080
rect 5592 35028 5598 35080
rect 5626 35028 5632 35080
rect 5684 35028 5690 35080
rect 7282 35028 7288 35080
rect 7340 35028 7346 35080
rect 7469 35071 7527 35077
rect 7469 35037 7481 35071
rect 7515 35037 7527 35071
rect 7469 35031 7527 35037
rect 7484 35000 7512 35031
rect 7650 35028 7656 35080
rect 7708 35028 7714 35080
rect 7852 35077 7880 35108
rect 7926 35096 7932 35108
rect 7984 35096 7990 35148
rect 7837 35071 7895 35077
rect 7837 35037 7849 35071
rect 7883 35037 7895 35071
rect 7837 35031 7895 35037
rect 7926 35000 7932 35012
rect 7484 34972 7932 35000
rect 7926 34960 7932 34972
rect 7984 34960 7990 35012
rect 7558 34892 7564 34944
rect 7616 34932 7622 34944
rect 8021 34935 8079 34941
rect 8021 34932 8033 34935
rect 7616 34904 8033 34932
rect 7616 34892 7622 34904
rect 8021 34901 8033 34904
rect 8067 34901 8079 34935
rect 8404 34932 8432 35176
rect 8754 35164 8760 35216
rect 8812 35204 8818 35216
rect 11698 35204 11704 35216
rect 8812 35176 11704 35204
rect 8812 35164 8818 35176
rect 9309 35071 9367 35077
rect 9309 35037 9321 35071
rect 9355 35068 9367 35071
rect 9416 35068 9444 35176
rect 11698 35164 11704 35176
rect 11756 35164 11762 35216
rect 11808 35204 11836 35244
rect 12250 35232 12256 35284
rect 12308 35272 12314 35284
rect 12618 35272 12624 35284
rect 12308 35244 12624 35272
rect 12308 35232 12314 35244
rect 12618 35232 12624 35244
rect 12676 35272 12682 35284
rect 14277 35275 14335 35281
rect 14277 35272 14289 35275
rect 12676 35244 14289 35272
rect 12676 35232 12682 35244
rect 14277 35241 14289 35244
rect 14323 35241 14335 35275
rect 14277 35235 14335 35241
rect 15654 35232 15660 35284
rect 15712 35232 15718 35284
rect 17862 35232 17868 35284
rect 17920 35272 17926 35284
rect 19705 35275 19763 35281
rect 19705 35272 19717 35275
rect 17920 35244 19717 35272
rect 17920 35232 17926 35244
rect 19705 35241 19717 35244
rect 19751 35241 19763 35275
rect 19705 35235 19763 35241
rect 20165 35275 20223 35281
rect 20165 35241 20177 35275
rect 20211 35272 20223 35275
rect 20438 35272 20444 35284
rect 20211 35244 20444 35272
rect 20211 35241 20223 35244
rect 20165 35235 20223 35241
rect 20438 35232 20444 35244
rect 20496 35232 20502 35284
rect 22278 35232 22284 35284
rect 22336 35232 22342 35284
rect 25130 35232 25136 35284
rect 25188 35232 25194 35284
rect 27062 35232 27068 35284
rect 27120 35232 27126 35284
rect 27798 35232 27804 35284
rect 27856 35232 27862 35284
rect 27890 35232 27896 35284
rect 27948 35232 27954 35284
rect 29546 35232 29552 35284
rect 29604 35272 29610 35284
rect 29825 35275 29883 35281
rect 29825 35272 29837 35275
rect 29604 35244 29837 35272
rect 29604 35232 29610 35244
rect 29825 35241 29837 35244
rect 29871 35241 29883 35275
rect 31202 35272 31208 35284
rect 29825 35235 29883 35241
rect 30760 35244 31208 35272
rect 14737 35207 14795 35213
rect 11808 35176 14320 35204
rect 9508 35108 11008 35136
rect 9508 35080 9536 35108
rect 9355 35040 9444 35068
rect 9355 35037 9367 35040
rect 9309 35031 9367 35037
rect 9490 35028 9496 35080
rect 9548 35028 9554 35080
rect 10226 35028 10232 35080
rect 10284 35068 10290 35080
rect 10778 35068 10784 35080
rect 10284 35040 10784 35068
rect 10284 35028 10290 35040
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 10980 35077 11008 35108
rect 10965 35071 11023 35077
rect 10965 35037 10977 35071
rect 11011 35068 11023 35071
rect 11698 35068 11704 35080
rect 11011 35040 11704 35068
rect 11011 35037 11023 35040
rect 10965 35031 11023 35037
rect 11698 35028 11704 35040
rect 11756 35028 11762 35080
rect 11790 35028 11796 35080
rect 11848 35068 11854 35080
rect 12069 35071 12127 35077
rect 12069 35068 12081 35071
rect 11848 35040 12081 35068
rect 11848 35028 11854 35040
rect 12069 35037 12081 35040
rect 12115 35037 12127 35071
rect 12069 35031 12127 35037
rect 12526 35028 12532 35080
rect 12584 35028 12590 35080
rect 14292 35077 14320 35176
rect 14737 35173 14749 35207
rect 14783 35173 14795 35207
rect 14737 35167 14795 35173
rect 15841 35207 15899 35213
rect 15841 35173 15853 35207
rect 15887 35204 15899 35207
rect 19886 35204 19892 35216
rect 15887 35176 19892 35204
rect 15887 35173 15899 35176
rect 15841 35167 15899 35173
rect 14366 35096 14372 35148
rect 14424 35096 14430 35148
rect 14277 35071 14335 35077
rect 14277 35037 14289 35071
rect 14323 35068 14335 35071
rect 14458 35068 14464 35080
rect 14323 35040 14464 35068
rect 14323 35037 14335 35040
rect 14277 35031 14335 35037
rect 14458 35028 14464 35040
rect 14516 35028 14522 35080
rect 14550 35028 14556 35080
rect 14608 35028 14614 35080
rect 14752 35068 14780 35167
rect 19886 35164 19892 35176
rect 19944 35164 19950 35216
rect 22094 35164 22100 35216
rect 22152 35204 22158 35216
rect 22554 35204 22560 35216
rect 22152 35176 22560 35204
rect 22152 35164 22158 35176
rect 22554 35164 22560 35176
rect 22612 35164 22618 35216
rect 27816 35204 27844 35232
rect 26988 35176 27844 35204
rect 23290 35136 23296 35148
rect 22296 35108 23296 35136
rect 22296 35077 22324 35108
rect 23290 35096 23296 35108
rect 23348 35096 23354 35148
rect 23382 35096 23388 35148
rect 23440 35136 23446 35148
rect 26988 35145 27016 35176
rect 27982 35164 27988 35216
rect 28040 35204 28046 35216
rect 30760 35204 30788 35244
rect 31202 35232 31208 35244
rect 31260 35232 31266 35284
rect 32309 35275 32367 35281
rect 32309 35272 32321 35275
rect 31312 35244 32321 35272
rect 28040 35176 30788 35204
rect 28040 35164 28046 35176
rect 26973 35139 27031 35145
rect 23440 35108 26188 35136
rect 23440 35096 23446 35108
rect 26160 35080 26188 35108
rect 26973 35105 26985 35139
rect 27019 35105 27031 35139
rect 26973 35099 27031 35105
rect 27062 35096 27068 35148
rect 27120 35096 27126 35148
rect 27157 35139 27215 35145
rect 27157 35105 27169 35139
rect 27203 35136 27215 35139
rect 28534 35136 28540 35148
rect 27203 35108 28540 35136
rect 27203 35105 27215 35108
rect 27157 35099 27215 35105
rect 19613 35071 19671 35077
rect 19613 35068 19625 35071
rect 14752 35040 19625 35068
rect 19613 35037 19625 35040
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 19981 35071 20039 35077
rect 19981 35037 19993 35071
rect 20027 35068 20039 35071
rect 22281 35071 22339 35077
rect 20027 35040 22094 35068
rect 20027 35037 20039 35040
rect 19981 35031 20039 35037
rect 8478 34960 8484 35012
rect 8536 35000 8542 35012
rect 9125 35003 9183 35009
rect 9125 35000 9137 35003
rect 8536 34972 9137 35000
rect 8536 34960 8542 34972
rect 9125 34969 9137 34972
rect 9171 34969 9183 35003
rect 9125 34963 9183 34969
rect 9766 34960 9772 35012
rect 9824 35000 9830 35012
rect 12544 35000 12572 35028
rect 9824 34972 12572 35000
rect 9824 34960 9830 34972
rect 15470 34960 15476 35012
rect 15528 34960 15534 35012
rect 17218 34960 17224 35012
rect 17276 34960 17282 35012
rect 17494 34960 17500 35012
rect 17552 35000 17558 35012
rect 17957 35003 18015 35009
rect 17957 35000 17969 35003
rect 17552 34972 17969 35000
rect 17552 34960 17558 34972
rect 17957 34969 17969 34972
rect 18003 34969 18015 35003
rect 17957 34963 18015 34969
rect 11054 34932 11060 34944
rect 8404 34904 11060 34932
rect 8021 34895 8079 34901
rect 11054 34892 11060 34904
rect 11112 34892 11118 34944
rect 11330 34892 11336 34944
rect 11388 34932 11394 34944
rect 12161 34935 12219 34941
rect 12161 34932 12173 34935
rect 11388 34904 12173 34932
rect 11388 34892 11394 34904
rect 12161 34901 12173 34904
rect 12207 34932 12219 34935
rect 15378 34932 15384 34944
rect 12207 34904 15384 34932
rect 12207 34901 12219 34904
rect 12161 34895 12219 34901
rect 15378 34892 15384 34904
rect 15436 34932 15442 34944
rect 15657 34935 15715 34941
rect 15657 34932 15669 34935
rect 15436 34904 15669 34932
rect 15436 34892 15442 34904
rect 15657 34901 15669 34904
rect 15703 34901 15715 34935
rect 22066 34932 22094 35040
rect 22281 35037 22293 35071
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 22462 35028 22468 35080
rect 22520 35028 22526 35080
rect 22925 35071 22983 35077
rect 22925 35037 22937 35071
rect 22971 35068 22983 35071
rect 23014 35068 23020 35080
rect 22971 35040 23020 35068
rect 22971 35037 22983 35040
rect 22925 35031 22983 35037
rect 23014 35028 23020 35040
rect 23072 35068 23078 35080
rect 23072 35040 23888 35068
rect 23072 35028 23078 35040
rect 23106 34960 23112 35012
rect 23164 34960 23170 35012
rect 23198 34960 23204 35012
rect 23256 35000 23262 35012
rect 23293 35003 23351 35009
rect 23293 35000 23305 35003
rect 23256 34972 23305 35000
rect 23256 34960 23262 34972
rect 23293 34969 23305 34972
rect 23339 34969 23351 35003
rect 23860 35000 23888 35040
rect 23934 35028 23940 35080
rect 23992 35068 23998 35080
rect 25501 35071 25559 35077
rect 25501 35068 25513 35071
rect 23992 35040 25513 35068
rect 23992 35028 23998 35040
rect 25501 35037 25513 35040
rect 25547 35068 25559 35071
rect 25774 35068 25780 35080
rect 25547 35040 25780 35068
rect 25547 35037 25559 35040
rect 25501 35031 25559 35037
rect 25774 35028 25780 35040
rect 25832 35028 25838 35080
rect 26142 35028 26148 35080
rect 26200 35028 26206 35080
rect 26234 35028 26240 35080
rect 26292 35028 26298 35080
rect 27080 35068 27108 35096
rect 27249 35071 27307 35077
rect 27249 35068 27261 35071
rect 27080 35040 27261 35068
rect 27249 35037 27261 35040
rect 27295 35068 27307 35071
rect 27522 35068 27528 35080
rect 27295 35040 27528 35068
rect 27295 35037 27307 35040
rect 27249 35031 27307 35037
rect 27522 35028 27528 35040
rect 27580 35028 27586 35080
rect 27614 35028 27620 35080
rect 27672 35068 27678 35080
rect 27908 35077 27936 35108
rect 28534 35096 28540 35108
rect 28592 35136 28598 35148
rect 30760 35145 30788 35176
rect 30834 35164 30840 35216
rect 30892 35164 30898 35216
rect 30926 35164 30932 35216
rect 30984 35204 30990 35216
rect 31312 35204 31340 35244
rect 32309 35241 32321 35244
rect 32355 35241 32367 35275
rect 32309 35235 32367 35241
rect 32582 35232 32588 35284
rect 32640 35272 32646 35284
rect 33413 35275 33471 35281
rect 33413 35272 33425 35275
rect 32640 35244 33425 35272
rect 32640 35232 32646 35244
rect 33413 35241 33425 35244
rect 33459 35241 33471 35275
rect 33413 35235 33471 35241
rect 34882 35232 34888 35284
rect 34940 35272 34946 35284
rect 35802 35272 35808 35284
rect 34940 35244 35808 35272
rect 34940 35232 34946 35244
rect 35802 35232 35808 35244
rect 35860 35232 35866 35284
rect 36449 35275 36507 35281
rect 36449 35241 36461 35275
rect 36495 35272 36507 35275
rect 38010 35272 38016 35284
rect 36495 35244 38016 35272
rect 36495 35241 36507 35244
rect 36449 35235 36507 35241
rect 38010 35232 38016 35244
rect 38068 35232 38074 35284
rect 30984 35176 31340 35204
rect 30984 35164 30990 35176
rect 31386 35164 31392 35216
rect 31444 35204 31450 35216
rect 33597 35207 33655 35213
rect 31444 35176 32444 35204
rect 31444 35164 31450 35176
rect 28905 35139 28963 35145
rect 28905 35136 28917 35139
rect 28592 35108 28917 35136
rect 28592 35096 28598 35108
rect 28905 35105 28917 35108
rect 28951 35105 28963 35139
rect 28905 35099 28963 35105
rect 29181 35139 29239 35145
rect 29181 35105 29193 35139
rect 29227 35136 29239 35139
rect 30745 35139 30803 35145
rect 29227 35108 29960 35136
rect 29227 35105 29239 35108
rect 29181 35099 29239 35105
rect 29932 35080 29960 35108
rect 30745 35105 30757 35139
rect 30791 35105 30803 35139
rect 30852 35136 30880 35164
rect 31849 35139 31907 35145
rect 31849 35136 31861 35139
rect 30852 35108 31861 35136
rect 30745 35099 30803 35105
rect 31849 35105 31861 35108
rect 31895 35136 31907 35139
rect 32122 35136 32128 35148
rect 31895 35108 32128 35136
rect 31895 35105 31907 35108
rect 31849 35099 31907 35105
rect 32122 35096 32128 35108
rect 32180 35096 32186 35148
rect 32416 35145 32444 35176
rect 33597 35173 33609 35207
rect 33643 35204 33655 35207
rect 33643 35176 36032 35204
rect 33643 35173 33655 35176
rect 33597 35167 33655 35173
rect 32401 35139 32459 35145
rect 32401 35105 32413 35139
rect 32447 35105 32459 35139
rect 32401 35099 32459 35105
rect 32766 35096 32772 35148
rect 32824 35096 32830 35148
rect 32950 35096 32956 35148
rect 33008 35136 33014 35148
rect 36004 35136 36032 35176
rect 36078 35164 36084 35216
rect 36136 35204 36142 35216
rect 37553 35207 37611 35213
rect 36136 35176 37320 35204
rect 36136 35164 36142 35176
rect 36722 35136 36728 35148
rect 33008 35108 34376 35136
rect 36004 35108 36728 35136
rect 33008 35096 33014 35108
rect 27709 35071 27767 35077
rect 27709 35068 27721 35071
rect 27672 35040 27721 35068
rect 27672 35028 27678 35040
rect 27709 35037 27721 35040
rect 27755 35037 27767 35071
rect 27709 35031 27767 35037
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35037 27951 35071
rect 27893 35031 27951 35037
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 28721 35071 28779 35077
rect 28721 35068 28733 35071
rect 28500 35040 28733 35068
rect 28500 35028 28506 35040
rect 28721 35037 28733 35040
rect 28767 35037 28779 35071
rect 28721 35031 28779 35037
rect 28810 35028 28816 35080
rect 28868 35028 28874 35080
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35037 29055 35071
rect 28997 35031 29055 35037
rect 24854 35000 24860 35012
rect 23860 34972 24860 35000
rect 23293 34963 23351 34969
rect 24854 34960 24860 34972
rect 24912 34960 24918 35012
rect 25038 34960 25044 35012
rect 25096 35000 25102 35012
rect 25317 35003 25375 35009
rect 25317 35000 25329 35003
rect 25096 34972 25329 35000
rect 25096 34960 25102 34972
rect 25317 34969 25329 34972
rect 25363 35000 25375 35003
rect 25866 35000 25872 35012
rect 25363 34972 25872 35000
rect 25363 34969 25375 34972
rect 25317 34963 25375 34969
rect 25866 34960 25872 34972
rect 25924 34960 25930 35012
rect 27062 34960 27068 35012
rect 27120 35000 27126 35012
rect 29012 35000 29040 35031
rect 29454 35028 29460 35080
rect 29512 35068 29518 35080
rect 29733 35071 29791 35077
rect 29733 35068 29745 35071
rect 29512 35040 29745 35068
rect 29512 35028 29518 35040
rect 29733 35037 29745 35040
rect 29779 35037 29791 35071
rect 29733 35031 29791 35037
rect 29914 35028 29920 35080
rect 29972 35028 29978 35080
rect 31297 35071 31355 35077
rect 31297 35037 31309 35071
rect 31343 35068 31355 35071
rect 31386 35068 31392 35080
rect 31343 35040 31392 35068
rect 31343 35037 31355 35040
rect 31297 35031 31355 35037
rect 31386 35028 31392 35040
rect 31444 35028 31450 35080
rect 31941 35071 31999 35077
rect 31941 35037 31953 35071
rect 31987 35068 31999 35071
rect 32030 35068 32036 35080
rect 31987 35040 32036 35068
rect 31987 35037 31999 35040
rect 31941 35031 31999 35037
rect 32030 35028 32036 35040
rect 32088 35028 32094 35080
rect 32416 35040 33364 35068
rect 27120 34972 29040 35000
rect 27120 34960 27126 34972
rect 25406 34932 25412 34944
rect 22066 34904 25412 34932
rect 15657 34895 15715 34901
rect 25406 34892 25412 34904
rect 25464 34932 25470 34944
rect 26053 34935 26111 34941
rect 26053 34932 26065 34935
rect 25464 34904 26065 34932
rect 25464 34892 25470 34904
rect 26053 34901 26065 34904
rect 26099 34901 26111 34935
rect 26053 34895 26111 34901
rect 27614 34892 27620 34944
rect 27672 34932 27678 34944
rect 28902 34932 28908 34944
rect 27672 34904 28908 34932
rect 27672 34892 27678 34904
rect 28902 34892 28908 34904
rect 28960 34892 28966 34944
rect 29012 34932 29040 34972
rect 29546 34960 29552 35012
rect 29604 35000 29610 35012
rect 32416 35000 32444 35040
rect 33229 35003 33287 35009
rect 33229 35000 33241 35003
rect 29604 34972 32444 35000
rect 32508 34972 33241 35000
rect 29604 34960 29610 34972
rect 30374 34932 30380 34944
rect 29012 34904 30380 34932
rect 30374 34892 30380 34904
rect 30432 34892 30438 34944
rect 30466 34892 30472 34944
rect 30524 34892 30530 34944
rect 30650 34892 30656 34944
rect 30708 34932 30714 34944
rect 32508 34932 32536 34972
rect 33229 34969 33241 34972
rect 33275 34969 33287 35003
rect 33336 35000 33364 35040
rect 33410 35028 33416 35080
rect 33468 35068 33474 35080
rect 33962 35068 33968 35080
rect 33468 35040 33968 35068
rect 33468 35028 33474 35040
rect 33962 35028 33968 35040
rect 34020 35068 34026 35080
rect 34348 35077 34376 35108
rect 36722 35096 36728 35108
rect 36780 35096 36786 35148
rect 37292 35136 37320 35176
rect 37553 35173 37565 35207
rect 37599 35204 37611 35207
rect 38102 35204 38108 35216
rect 37599 35176 38108 35204
rect 37599 35173 37611 35176
rect 37553 35167 37611 35173
rect 38102 35164 38108 35176
rect 38160 35204 38166 35216
rect 38160 35176 38240 35204
rect 38160 35164 38166 35176
rect 37734 35136 37740 35148
rect 37292 35108 37740 35136
rect 34149 35071 34207 35077
rect 34149 35068 34161 35071
rect 34020 35040 34161 35068
rect 34020 35028 34026 35040
rect 34149 35037 34161 35040
rect 34195 35037 34207 35071
rect 34149 35031 34207 35037
rect 34333 35071 34391 35077
rect 34333 35037 34345 35071
rect 34379 35037 34391 35071
rect 34333 35031 34391 35037
rect 35802 35028 35808 35080
rect 35860 35028 35866 35080
rect 35894 35028 35900 35080
rect 35952 35068 35958 35080
rect 36311 35071 36369 35077
rect 35952 35040 35997 35068
rect 35952 35028 35958 35040
rect 36311 35037 36323 35071
rect 36357 35068 36369 35071
rect 36446 35068 36452 35080
rect 36357 35040 36452 35068
rect 36357 35037 36369 35040
rect 36311 35031 36369 35037
rect 35710 35000 35716 35012
rect 33336 34972 35716 35000
rect 33229 34963 33287 34969
rect 35710 34960 35716 34972
rect 35768 34960 35774 35012
rect 36078 34960 36084 35012
rect 36136 34960 36142 35012
rect 36170 34960 36176 35012
rect 36228 34960 36234 35012
rect 30708 34904 32536 34932
rect 30708 34892 30714 34904
rect 33042 34892 33048 34944
rect 33100 34932 33106 34944
rect 33413 34935 33471 34941
rect 33413 34932 33425 34935
rect 33100 34904 33425 34932
rect 33100 34892 33106 34904
rect 33413 34901 33425 34904
rect 33459 34901 33471 34935
rect 33413 34895 33471 34901
rect 34238 34892 34244 34944
rect 34296 34892 34302 34944
rect 35342 34892 35348 34944
rect 35400 34932 35406 34944
rect 36326 34932 36354 35031
rect 36446 35028 36452 35040
rect 36504 35028 36510 35080
rect 36906 35028 36912 35080
rect 36964 35028 36970 35080
rect 37047 35071 37105 35077
rect 37047 35037 37059 35071
rect 37093 35037 37105 35071
rect 37292 35068 37320 35108
rect 37734 35096 37740 35108
rect 37792 35096 37798 35148
rect 38212 35145 38240 35176
rect 38197 35139 38255 35145
rect 38197 35105 38209 35139
rect 38243 35105 38255 35139
rect 38197 35099 38255 35105
rect 38657 35139 38715 35145
rect 38657 35105 38669 35139
rect 38703 35105 38715 35139
rect 38657 35099 38715 35105
rect 37047 35031 37105 35037
rect 37200 35040 37320 35068
rect 35400 34904 36354 34932
rect 37072 34932 37100 35031
rect 37200 35009 37228 35040
rect 37366 35028 37372 35080
rect 37424 35077 37430 35080
rect 37424 35071 37473 35077
rect 37424 35037 37427 35071
rect 37461 35068 37473 35071
rect 37826 35068 37832 35080
rect 37461 35040 37832 35068
rect 37461 35037 37473 35040
rect 37424 35031 37473 35037
rect 37424 35028 37430 35031
rect 37826 35028 37832 35040
rect 37884 35028 37890 35080
rect 38289 35071 38347 35077
rect 38289 35037 38301 35071
rect 38335 35068 38347 35071
rect 38378 35068 38384 35080
rect 38335 35040 38384 35068
rect 38335 35037 38347 35040
rect 38289 35031 38347 35037
rect 38378 35028 38384 35040
rect 38436 35028 38442 35080
rect 37185 35003 37243 35009
rect 37185 34969 37197 35003
rect 37231 34969 37243 35003
rect 37185 34963 37243 34969
rect 37274 34960 37280 35012
rect 37332 34960 37338 35012
rect 38672 35000 38700 35099
rect 40034 35096 40040 35148
rect 40092 35096 40098 35148
rect 42245 35139 42303 35145
rect 42245 35105 42257 35139
rect 42291 35136 42303 35139
rect 43990 35136 43996 35148
rect 42291 35108 43996 35136
rect 42291 35105 42303 35108
rect 42245 35099 42303 35105
rect 43990 35096 43996 35108
rect 44048 35096 44054 35148
rect 40052 35068 40080 35096
rect 41414 35068 41420 35080
rect 40052 35040 41420 35068
rect 41414 35028 41420 35040
rect 41472 35068 41478 35080
rect 41874 35068 41880 35080
rect 41472 35040 41880 35068
rect 41472 35028 41478 35040
rect 41874 35028 41880 35040
rect 41932 35028 41938 35080
rect 41966 35028 41972 35080
rect 42024 35028 42030 35080
rect 42886 35028 42892 35080
rect 42944 35028 42950 35080
rect 40282 35003 40340 35009
rect 40282 35000 40294 35003
rect 38672 34972 40294 35000
rect 40282 34969 40294 34972
rect 40328 34969 40340 35003
rect 40282 34963 40340 34969
rect 40586 34960 40592 35012
rect 40644 35000 40650 35012
rect 41230 35000 41236 35012
rect 40644 34972 41236 35000
rect 40644 34960 40650 34972
rect 41230 34960 41236 34972
rect 41288 34960 41294 35012
rect 43165 35003 43223 35009
rect 43165 34969 43177 35003
rect 43211 35000 43223 35003
rect 43990 35000 43996 35012
rect 43211 34972 43996 35000
rect 43211 34969 43223 34972
rect 43165 34963 43223 34969
rect 43990 34960 43996 34972
rect 44048 34960 44054 35012
rect 40770 34932 40776 34944
rect 37072 34904 40776 34932
rect 35400 34892 35406 34904
rect 40770 34892 40776 34904
rect 40828 34932 40834 34944
rect 41417 34935 41475 34941
rect 41417 34932 41429 34935
rect 40828 34904 41429 34932
rect 40828 34892 40834 34904
rect 41417 34901 41429 34904
rect 41463 34901 41475 34935
rect 41417 34895 41475 34901
rect 1104 34842 43884 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 43884 34842
rect 1104 34768 43884 34790
rect 8938 34688 8944 34740
rect 8996 34728 9002 34740
rect 9398 34728 9404 34740
rect 8996 34700 9404 34728
rect 8996 34688 9002 34700
rect 9398 34688 9404 34700
rect 9456 34688 9462 34740
rect 9858 34688 9864 34740
rect 9916 34728 9922 34740
rect 9916 34700 13952 34728
rect 9916 34688 9922 34700
rect 4614 34660 4620 34672
rect 4172 34632 4620 34660
rect 4172 34601 4200 34632
rect 4614 34620 4620 34632
rect 4672 34620 4678 34672
rect 7558 34620 7564 34672
rect 7616 34620 7622 34672
rect 9217 34663 9275 34669
rect 9217 34660 9229 34663
rect 7760 34632 9229 34660
rect 4157 34595 4215 34601
rect 4157 34561 4169 34595
rect 4203 34561 4215 34595
rect 4157 34555 4215 34561
rect 4424 34595 4482 34601
rect 4424 34561 4436 34595
rect 4470 34592 4482 34595
rect 5810 34592 5816 34604
rect 4470 34564 5816 34592
rect 4470 34561 4482 34564
rect 4424 34555 4482 34561
rect 5810 34552 5816 34564
rect 5868 34552 5874 34604
rect 7098 34552 7104 34604
rect 7156 34552 7162 34604
rect 7282 34552 7288 34604
rect 7340 34592 7346 34604
rect 7760 34592 7788 34632
rect 9217 34629 9229 34632
rect 9263 34629 9275 34663
rect 9674 34660 9680 34672
rect 9217 34623 9275 34629
rect 9324 34632 9680 34660
rect 7340 34564 7788 34592
rect 7340 34552 7346 34564
rect 8478 34552 8484 34604
rect 8536 34552 8542 34604
rect 8665 34595 8723 34601
rect 8665 34561 8677 34595
rect 8711 34592 8723 34595
rect 9324 34592 9352 34632
rect 9674 34620 9680 34632
rect 9732 34620 9738 34672
rect 10060 34604 10088 34700
rect 10594 34620 10600 34672
rect 10652 34660 10658 34672
rect 10652 34632 12020 34660
rect 10652 34620 10658 34632
rect 8711 34564 9352 34592
rect 8711 34561 8723 34564
rect 8665 34555 8723 34561
rect 9398 34552 9404 34604
rect 9456 34552 9462 34604
rect 10042 34552 10048 34604
rect 10100 34552 10106 34604
rect 10229 34595 10287 34601
rect 10229 34561 10241 34595
rect 10275 34561 10287 34595
rect 10229 34555 10287 34561
rect 8386 34484 8392 34536
rect 8444 34484 8450 34536
rect 8846 34524 8852 34536
rect 8496 34496 8852 34524
rect 7558 34416 7564 34468
rect 7616 34456 7622 34468
rect 8496 34456 8524 34496
rect 8846 34484 8852 34496
rect 8904 34484 8910 34536
rect 9214 34484 9220 34536
rect 9272 34524 9278 34536
rect 9585 34527 9643 34533
rect 9585 34524 9597 34527
rect 9272 34496 9597 34524
rect 9272 34484 9278 34496
rect 9585 34493 9597 34496
rect 9631 34524 9643 34527
rect 10244 34524 10272 34555
rect 11698 34552 11704 34604
rect 11756 34552 11762 34604
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34561 11943 34595
rect 11992 34592 12020 34632
rect 12434 34620 12440 34672
rect 12492 34660 12498 34672
rect 12897 34663 12955 34669
rect 12897 34660 12909 34663
rect 12492 34632 12909 34660
rect 12492 34620 12498 34632
rect 12897 34629 12909 34632
rect 12943 34629 12955 34663
rect 12897 34623 12955 34629
rect 13078 34620 13084 34672
rect 13136 34660 13142 34672
rect 13722 34660 13728 34672
rect 13136 34632 13728 34660
rect 13136 34620 13142 34632
rect 13722 34620 13728 34632
rect 13780 34620 13786 34672
rect 12710 34592 12716 34604
rect 11992 34564 12716 34592
rect 11885 34555 11943 34561
rect 9631 34496 10272 34524
rect 9631 34493 9643 34496
rect 9585 34487 9643 34493
rect 10244 34468 10272 34496
rect 10318 34484 10324 34536
rect 10376 34524 10382 34536
rect 11793 34527 11851 34533
rect 11793 34524 11805 34527
rect 10376 34496 11805 34524
rect 10376 34484 10382 34496
rect 11793 34493 11805 34496
rect 11839 34493 11851 34527
rect 11900 34524 11928 34555
rect 12710 34552 12716 34564
rect 12768 34552 12774 34604
rect 13096 34524 13124 34620
rect 13538 34552 13544 34604
rect 13596 34552 13602 34604
rect 13814 34552 13820 34604
rect 13872 34552 13878 34604
rect 13924 34592 13952 34700
rect 17954 34688 17960 34740
rect 18012 34728 18018 34740
rect 19521 34731 19579 34737
rect 19521 34728 19533 34731
rect 18012 34700 19533 34728
rect 18012 34688 18018 34700
rect 19521 34697 19533 34700
rect 19567 34728 19579 34731
rect 22738 34728 22744 34740
rect 19567 34700 22744 34728
rect 19567 34697 19579 34700
rect 19521 34691 19579 34697
rect 22738 34688 22744 34700
rect 22796 34688 22802 34740
rect 24578 34688 24584 34740
rect 24636 34728 24642 34740
rect 28166 34728 28172 34740
rect 24636 34700 28172 34728
rect 24636 34688 24642 34700
rect 28166 34688 28172 34700
rect 28224 34688 28230 34740
rect 28442 34688 28448 34740
rect 28500 34728 28506 34740
rect 31294 34728 31300 34740
rect 28500 34700 31300 34728
rect 28500 34688 28506 34700
rect 31294 34688 31300 34700
rect 31352 34688 31358 34740
rect 31478 34688 31484 34740
rect 31536 34728 31542 34740
rect 32582 34728 32588 34740
rect 31536 34700 32588 34728
rect 31536 34688 31542 34700
rect 32582 34688 32588 34700
rect 32640 34688 32646 34740
rect 33042 34688 33048 34740
rect 33100 34688 33106 34740
rect 33134 34688 33140 34740
rect 33192 34728 33198 34740
rect 34422 34728 34428 34740
rect 33192 34700 34428 34728
rect 33192 34688 33198 34700
rect 34422 34688 34428 34700
rect 34480 34688 34486 34740
rect 35802 34688 35808 34740
rect 35860 34728 35866 34740
rect 35989 34731 36047 34737
rect 35989 34728 36001 34731
rect 35860 34700 36001 34728
rect 35860 34688 35866 34700
rect 35989 34697 36001 34700
rect 36035 34697 36047 34731
rect 35989 34691 36047 34697
rect 36722 34688 36728 34740
rect 36780 34728 36786 34740
rect 38470 34728 38476 34740
rect 36780 34700 38476 34728
rect 36780 34688 36786 34700
rect 38470 34688 38476 34700
rect 38528 34728 38534 34740
rect 38528 34700 41414 34728
rect 38528 34688 38534 34700
rect 14461 34663 14519 34669
rect 14461 34629 14473 34663
rect 14507 34660 14519 34663
rect 17034 34660 17040 34672
rect 14507 34632 17040 34660
rect 14507 34629 14519 34632
rect 14461 34623 14519 34629
rect 14369 34595 14427 34601
rect 14369 34592 14381 34595
rect 13924 34564 14381 34592
rect 14369 34561 14381 34564
rect 14415 34561 14427 34595
rect 14369 34555 14427 34561
rect 11900 34496 13124 34524
rect 13909 34527 13967 34533
rect 11793 34487 11851 34493
rect 13909 34493 13921 34527
rect 13955 34524 13967 34527
rect 14458 34524 14464 34536
rect 13955 34496 14464 34524
rect 13955 34493 13967 34496
rect 13909 34487 13967 34493
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 7616 34428 8524 34456
rect 7616 34416 7622 34428
rect 10226 34416 10232 34468
rect 10284 34456 10290 34468
rect 10284 34428 12434 34456
rect 10284 34416 10290 34428
rect 5537 34391 5595 34397
rect 5537 34357 5549 34391
rect 5583 34388 5595 34391
rect 6362 34388 6368 34400
rect 5583 34360 6368 34388
rect 5583 34357 5595 34360
rect 5537 34351 5595 34357
rect 6362 34348 6368 34360
rect 6420 34348 6426 34400
rect 6914 34348 6920 34400
rect 6972 34348 6978 34400
rect 7466 34348 7472 34400
rect 7524 34348 7530 34400
rect 9674 34348 9680 34400
rect 9732 34388 9738 34400
rect 10137 34391 10195 34397
rect 10137 34388 10149 34391
rect 9732 34360 10149 34388
rect 9732 34348 9738 34360
rect 10137 34357 10149 34360
rect 10183 34357 10195 34391
rect 12406 34388 12434 34428
rect 12894 34416 12900 34468
rect 12952 34456 12958 34468
rect 13538 34456 13544 34468
rect 12952 34428 13544 34456
rect 12952 34416 12958 34428
rect 13538 34416 13544 34428
rect 13596 34456 13602 34468
rect 14568 34456 14596 34632
rect 17034 34620 17040 34632
rect 17092 34620 17098 34672
rect 18230 34620 18236 34672
rect 18288 34660 18294 34672
rect 18386 34663 18444 34669
rect 18386 34660 18398 34663
rect 18288 34632 18398 34660
rect 18288 34620 18294 34632
rect 18386 34629 18398 34632
rect 18432 34629 18444 34663
rect 24854 34660 24860 34672
rect 18386 34623 18444 34629
rect 22066 34632 24860 34660
rect 17218 34552 17224 34604
rect 17276 34592 17282 34604
rect 18141 34595 18199 34601
rect 18141 34592 18153 34595
rect 17276 34564 18153 34592
rect 17276 34552 17282 34564
rect 18141 34561 18153 34564
rect 18187 34561 18199 34595
rect 19518 34592 19524 34604
rect 18141 34555 18199 34561
rect 18248 34564 19524 34592
rect 15470 34484 15476 34536
rect 15528 34524 15534 34536
rect 18248 34524 18276 34564
rect 19518 34552 19524 34564
rect 19576 34552 19582 34604
rect 15528 34496 18276 34524
rect 15528 34484 15534 34496
rect 19150 34484 19156 34536
rect 19208 34524 19214 34536
rect 22066 34524 22094 34632
rect 24854 34620 24860 34632
rect 24912 34620 24918 34672
rect 25774 34620 25780 34672
rect 25832 34620 25838 34672
rect 27154 34660 27160 34672
rect 26160 34632 27160 34660
rect 22462 34552 22468 34604
rect 22520 34592 22526 34604
rect 23109 34595 23167 34601
rect 23109 34592 23121 34595
rect 22520 34564 23121 34592
rect 22520 34552 22526 34564
rect 23109 34561 23121 34564
rect 23155 34561 23167 34595
rect 23109 34555 23167 34561
rect 23201 34595 23259 34601
rect 23201 34561 23213 34595
rect 23247 34592 23259 34595
rect 23382 34592 23388 34604
rect 23247 34564 23388 34592
rect 23247 34561 23259 34564
rect 23201 34555 23259 34561
rect 19208 34496 22094 34524
rect 23124 34524 23152 34555
rect 23382 34552 23388 34564
rect 23440 34552 23446 34604
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 23934 34592 23940 34604
rect 23799 34564 23940 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 23934 34552 23940 34564
rect 23992 34552 23998 34604
rect 24121 34595 24179 34601
rect 24121 34561 24133 34595
rect 24167 34592 24179 34595
rect 24302 34592 24308 34604
rect 24167 34564 24308 34592
rect 24167 34561 24179 34564
rect 24121 34555 24179 34561
rect 24302 34552 24308 34564
rect 24360 34552 24366 34604
rect 25225 34595 25283 34601
rect 25225 34561 25237 34595
rect 25271 34592 25283 34595
rect 25314 34592 25320 34604
rect 25271 34564 25320 34592
rect 25271 34561 25283 34564
rect 25225 34555 25283 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 26160 34601 26188 34632
rect 27154 34620 27160 34632
rect 27212 34620 27218 34672
rect 27801 34663 27859 34669
rect 27356 34632 27660 34660
rect 26145 34595 26203 34601
rect 26145 34561 26157 34595
rect 26191 34561 26203 34595
rect 26145 34555 26203 34561
rect 26326 34552 26332 34604
rect 26384 34592 26390 34604
rect 27356 34592 27384 34632
rect 27632 34601 27660 34632
rect 27801 34629 27813 34663
rect 27847 34660 27859 34663
rect 28074 34660 28080 34672
rect 27847 34632 28080 34660
rect 27847 34629 27859 34632
rect 27801 34623 27859 34629
rect 28074 34620 28080 34632
rect 28132 34660 28138 34672
rect 28626 34660 28632 34672
rect 28132 34632 28632 34660
rect 28132 34620 28138 34632
rect 28626 34620 28632 34632
rect 28684 34620 28690 34672
rect 28902 34660 28908 34672
rect 28736 34632 28908 34660
rect 26384 34564 27384 34592
rect 27525 34595 27583 34601
rect 26384 34552 26390 34564
rect 27525 34561 27537 34595
rect 27571 34561 27583 34595
rect 27525 34555 27583 34561
rect 27617 34595 27675 34601
rect 27617 34561 27629 34595
rect 27663 34561 27675 34595
rect 27617 34555 27675 34561
rect 25038 34524 25044 34536
rect 23124 34496 25044 34524
rect 19208 34484 19214 34496
rect 25038 34484 25044 34496
rect 25096 34484 25102 34536
rect 25866 34484 25872 34536
rect 25924 34524 25930 34536
rect 25961 34527 26019 34533
rect 25961 34524 25973 34527
rect 25924 34496 25973 34524
rect 25924 34484 25930 34496
rect 25961 34493 25973 34496
rect 26007 34493 26019 34527
rect 25961 34487 26019 34493
rect 26053 34527 26111 34533
rect 26053 34493 26065 34527
rect 26099 34524 26111 34527
rect 27540 34524 27568 34555
rect 28350 34552 28356 34604
rect 28408 34592 28414 34604
rect 28736 34601 28764 34632
rect 28902 34620 28908 34632
rect 28960 34620 28966 34672
rect 29178 34620 29184 34672
rect 29236 34660 29242 34672
rect 34517 34663 34575 34669
rect 34517 34660 34529 34663
rect 29236 34632 34529 34660
rect 29236 34620 29242 34632
rect 34517 34629 34529 34632
rect 34563 34629 34575 34663
rect 34517 34623 34575 34629
rect 35894 34620 35900 34672
rect 35952 34660 35958 34672
rect 40310 34660 40316 34672
rect 35952 34632 40316 34660
rect 35952 34620 35958 34632
rect 40310 34620 40316 34632
rect 40368 34620 40374 34672
rect 41386 34660 41414 34700
rect 42797 34663 42855 34669
rect 42797 34660 42809 34663
rect 41386 34632 42809 34660
rect 42797 34629 42809 34632
rect 42843 34629 42855 34663
rect 42797 34623 42855 34629
rect 28721 34595 28779 34601
rect 28408 34564 28672 34592
rect 28408 34552 28414 34564
rect 27706 34524 27712 34536
rect 26099 34496 26280 34524
rect 27540 34496 27712 34524
rect 26099 34493 26111 34496
rect 26053 34487 26111 34493
rect 13596 34428 14596 34456
rect 23017 34459 23075 34465
rect 13596 34416 13602 34428
rect 23017 34425 23029 34459
rect 23063 34456 23075 34459
rect 23106 34456 23112 34468
rect 23063 34428 23112 34456
rect 23063 34425 23075 34428
rect 23017 34419 23075 34425
rect 23106 34416 23112 34428
rect 23164 34416 23170 34468
rect 24762 34416 24768 34468
rect 24820 34456 24826 34468
rect 26252 34456 26280 34496
rect 27706 34484 27712 34496
rect 27764 34484 27770 34536
rect 27798 34484 27804 34536
rect 27856 34524 27862 34536
rect 28445 34527 28503 34533
rect 28445 34524 28457 34527
rect 27856 34496 28457 34524
rect 27856 34484 27862 34496
rect 28445 34493 28457 34496
rect 28491 34493 28503 34527
rect 28644 34524 28672 34564
rect 28721 34561 28733 34595
rect 28767 34561 28779 34595
rect 28721 34555 28779 34561
rect 28828 34564 30328 34592
rect 28828 34524 28856 34564
rect 28644 34496 28856 34524
rect 28997 34527 29055 34533
rect 28445 34487 28503 34493
rect 28997 34493 29009 34527
rect 29043 34524 29055 34527
rect 29454 34524 29460 34536
rect 29043 34496 29460 34524
rect 29043 34493 29055 34496
rect 28997 34487 29055 34493
rect 29454 34484 29460 34496
rect 29512 34484 29518 34536
rect 30300 34524 30328 34564
rect 31294 34552 31300 34604
rect 31352 34552 31358 34604
rect 33226 34552 33232 34604
rect 33284 34552 33290 34604
rect 33686 34552 33692 34604
rect 33744 34552 33750 34604
rect 34422 34552 34428 34604
rect 34480 34592 34486 34604
rect 35986 34592 35992 34604
rect 34480 34564 35992 34592
rect 34480 34552 34486 34564
rect 35986 34552 35992 34564
rect 36044 34592 36050 34604
rect 36127 34595 36185 34601
rect 36127 34592 36139 34595
rect 36044 34564 36139 34592
rect 36044 34552 36050 34564
rect 36127 34561 36139 34564
rect 36173 34561 36185 34595
rect 36127 34555 36185 34561
rect 36265 34595 36323 34601
rect 36265 34561 36277 34595
rect 36311 34561 36323 34595
rect 36265 34555 36323 34561
rect 31386 34524 31392 34536
rect 30300 34496 31392 34524
rect 31386 34484 31392 34496
rect 31444 34484 31450 34536
rect 32490 34484 32496 34536
rect 32548 34524 32554 34536
rect 33321 34527 33379 34533
rect 33321 34524 33333 34527
rect 32548 34496 33333 34524
rect 32548 34484 32554 34496
rect 33321 34493 33333 34496
rect 33367 34493 33379 34527
rect 33321 34487 33379 34493
rect 34882 34484 34888 34536
rect 34940 34484 34946 34536
rect 35253 34527 35311 34533
rect 35253 34493 35265 34527
rect 35299 34524 35311 34527
rect 36280 34524 36308 34555
rect 36354 34552 36360 34604
rect 36412 34552 36418 34604
rect 36446 34552 36452 34604
rect 36504 34601 36510 34604
rect 36504 34595 36543 34601
rect 36531 34561 36543 34595
rect 36504 34555 36543 34561
rect 36504 34552 36510 34555
rect 36630 34552 36636 34604
rect 36688 34552 36694 34604
rect 38194 34524 38200 34536
rect 35299 34496 36124 34524
rect 35299 34493 35311 34496
rect 35253 34487 35311 34493
rect 26970 34456 26976 34468
rect 24820 34428 26096 34456
rect 26252 34428 26976 34456
rect 24820 34416 24826 34428
rect 14274 34388 14280 34400
rect 12406 34360 14280 34388
rect 10137 34351 10195 34357
rect 14274 34348 14280 34360
rect 14332 34348 14338 34400
rect 25406 34348 25412 34400
rect 25464 34388 25470 34400
rect 25961 34391 26019 34397
rect 25961 34388 25973 34391
rect 25464 34360 25973 34388
rect 25464 34348 25470 34360
rect 25961 34357 25973 34360
rect 26007 34357 26019 34391
rect 26068 34388 26096 34428
rect 26970 34416 26976 34428
rect 27028 34456 27034 34468
rect 29086 34456 29092 34468
rect 27028 34428 29092 34456
rect 27028 34416 27034 34428
rect 29086 34416 29092 34428
rect 29144 34416 29150 34468
rect 29638 34416 29644 34468
rect 29696 34456 29702 34468
rect 34146 34456 34152 34468
rect 29696 34428 34152 34456
rect 29696 34416 29702 34428
rect 34146 34416 34152 34428
rect 34204 34416 34210 34468
rect 34238 34416 34244 34468
rect 34296 34456 34302 34468
rect 34655 34459 34713 34465
rect 34655 34456 34667 34459
rect 34296 34428 34667 34456
rect 34296 34416 34302 34428
rect 34655 34425 34667 34428
rect 34701 34425 34713 34459
rect 34655 34419 34713 34425
rect 28442 34388 28448 34400
rect 26068 34360 28448 34388
rect 25961 34351 26019 34357
rect 28442 34348 28448 34360
rect 28500 34388 28506 34400
rect 28537 34391 28595 34397
rect 28537 34388 28549 34391
rect 28500 34360 28549 34388
rect 28500 34348 28506 34360
rect 28537 34357 28549 34360
rect 28583 34357 28595 34391
rect 28537 34351 28595 34357
rect 28629 34391 28687 34397
rect 28629 34357 28641 34391
rect 28675 34388 28687 34391
rect 28994 34388 29000 34400
rect 28675 34360 29000 34388
rect 28675 34357 28687 34360
rect 28629 34351 28687 34357
rect 28994 34348 29000 34360
rect 29052 34388 29058 34400
rect 30006 34388 30012 34400
rect 29052 34360 30012 34388
rect 29052 34348 29058 34360
rect 30006 34348 30012 34360
rect 30064 34348 30070 34400
rect 32858 34348 32864 34400
rect 32916 34388 32922 34400
rect 33042 34388 33048 34400
rect 32916 34360 33048 34388
rect 32916 34348 32922 34360
rect 33042 34348 33048 34360
rect 33100 34348 33106 34400
rect 33594 34348 33600 34400
rect 33652 34348 33658 34400
rect 34793 34391 34851 34397
rect 34793 34357 34805 34391
rect 34839 34388 34851 34391
rect 35802 34388 35808 34400
rect 34839 34360 35808 34388
rect 34839 34357 34851 34360
rect 34793 34351 34851 34357
rect 35802 34348 35808 34360
rect 35860 34348 35866 34400
rect 36096 34388 36124 34496
rect 36188 34496 36308 34524
rect 36372 34496 38200 34524
rect 36188 34468 36216 34496
rect 36170 34416 36176 34468
rect 36228 34416 36234 34468
rect 36372 34388 36400 34496
rect 38194 34484 38200 34496
rect 38252 34484 38258 34536
rect 36096 34360 36400 34388
rect 43073 34391 43131 34397
rect 43073 34357 43085 34391
rect 43119 34388 43131 34391
rect 43254 34388 43260 34400
rect 43119 34360 43260 34388
rect 43119 34357 43131 34360
rect 43073 34351 43131 34357
rect 43254 34348 43260 34360
rect 43312 34348 43318 34400
rect 1104 34298 43884 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 43884 34298
rect 1104 34224 43884 34246
rect 5810 34144 5816 34196
rect 5868 34144 5874 34196
rect 7466 34144 7472 34196
rect 7524 34184 7530 34196
rect 8021 34187 8079 34193
rect 8021 34184 8033 34187
rect 7524 34156 8033 34184
rect 7524 34144 7530 34156
rect 8021 34153 8033 34156
rect 8067 34153 8079 34187
rect 8021 34147 8079 34153
rect 8110 34144 8116 34196
rect 8168 34184 8174 34196
rect 26697 34187 26755 34193
rect 8168 34156 19472 34184
rect 8168 34144 8174 34156
rect 7098 34116 7104 34128
rect 6012 34088 7104 34116
rect 6012 33989 6040 34088
rect 7098 34076 7104 34088
rect 7156 34076 7162 34128
rect 10778 34076 10784 34128
rect 10836 34116 10842 34128
rect 10836 34088 11100 34116
rect 10836 34076 10842 34088
rect 6181 34051 6239 34057
rect 6181 34017 6193 34051
rect 6227 34048 6239 34051
rect 6638 34048 6644 34060
rect 6227 34020 6644 34048
rect 6227 34017 6239 34020
rect 6181 34011 6239 34017
rect 6638 34008 6644 34020
rect 6696 34008 6702 34060
rect 8478 34048 8484 34060
rect 8036 34020 8484 34048
rect 5997 33983 6055 33989
rect 5997 33949 6009 33983
rect 6043 33949 6055 33983
rect 5997 33943 6055 33949
rect 6089 33983 6147 33989
rect 6089 33949 6101 33983
rect 6135 33949 6147 33983
rect 6089 33943 6147 33949
rect 6273 33983 6331 33989
rect 6273 33949 6285 33983
rect 6319 33980 6331 33983
rect 6362 33980 6368 33992
rect 6319 33952 6368 33980
rect 6319 33949 6331 33952
rect 6273 33943 6331 33949
rect 6104 33912 6132 33943
rect 6362 33940 6368 33952
rect 6420 33940 6426 33992
rect 6454 33940 6460 33992
rect 6512 33940 6518 33992
rect 6917 33983 6975 33989
rect 6917 33949 6929 33983
rect 6963 33980 6975 33983
rect 7006 33980 7012 33992
rect 6963 33952 7012 33980
rect 6963 33949 6975 33952
rect 6917 33943 6975 33949
rect 7006 33940 7012 33952
rect 7064 33940 7070 33992
rect 8036 33989 8064 34020
rect 8478 34008 8484 34020
rect 8536 34008 8542 34060
rect 8570 34008 8576 34060
rect 8628 34048 8634 34060
rect 10045 34051 10103 34057
rect 10045 34048 10057 34051
rect 8628 34020 10057 34048
rect 8628 34008 8634 34020
rect 10045 34017 10057 34020
rect 10091 34017 10103 34051
rect 10045 34011 10103 34017
rect 10226 34008 10232 34060
rect 10284 34008 10290 34060
rect 10318 34008 10324 34060
rect 10376 34008 10382 34060
rect 10873 34051 10931 34057
rect 10873 34017 10885 34051
rect 10919 34048 10931 34051
rect 10962 34048 10968 34060
rect 10919 34020 10968 34048
rect 10919 34017 10931 34020
rect 10873 34011 10931 34017
rect 10962 34008 10968 34020
rect 11020 34008 11026 34060
rect 11072 34048 11100 34088
rect 11146 34076 11152 34128
rect 11204 34116 11210 34128
rect 11422 34116 11428 34128
rect 11204 34088 11428 34116
rect 11204 34076 11210 34088
rect 11422 34076 11428 34088
rect 11480 34116 11486 34128
rect 12158 34116 12164 34128
rect 11480 34088 12164 34116
rect 11480 34076 11486 34088
rect 12158 34076 12164 34088
rect 12216 34076 12222 34128
rect 13449 34051 13507 34057
rect 13449 34048 13461 34051
rect 11072 34020 11284 34048
rect 7101 33983 7159 33989
rect 7101 33949 7113 33983
rect 7147 33980 7159 33983
rect 8021 33983 8079 33989
rect 8021 33980 8033 33983
rect 7147 33952 8033 33980
rect 7147 33949 7159 33952
rect 7101 33943 7159 33949
rect 8021 33949 8033 33952
rect 8067 33949 8079 33983
rect 8297 33983 8355 33989
rect 8297 33980 8309 33983
rect 8021 33943 8079 33949
rect 8128 33952 8309 33980
rect 6730 33912 6736 33924
rect 6104 33884 6736 33912
rect 6730 33872 6736 33884
rect 6788 33872 6794 33924
rect 7024 33912 7052 33940
rect 7834 33912 7840 33924
rect 7024 33884 7840 33912
rect 7834 33872 7840 33884
rect 7892 33872 7898 33924
rect 7926 33872 7932 33924
rect 7984 33912 7990 33924
rect 8128 33912 8156 33952
rect 8297 33949 8309 33952
rect 8343 33949 8355 33983
rect 8297 33943 8355 33949
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 11256 33989 11284 34020
rect 12406 34020 13461 34048
rect 10137 33983 10195 33989
rect 10137 33980 10149 33983
rect 9456 33952 10149 33980
rect 9456 33940 9462 33952
rect 10137 33949 10149 33952
rect 10183 33949 10195 33983
rect 10137 33943 10195 33949
rect 11241 33983 11299 33989
rect 11241 33949 11253 33983
rect 11287 33949 11299 33983
rect 11241 33943 11299 33949
rect 11333 33983 11391 33989
rect 11333 33949 11345 33983
rect 11379 33980 11391 33983
rect 12406 33980 12434 34020
rect 13449 34017 13461 34020
rect 13495 34017 13507 34051
rect 13449 34011 13507 34017
rect 11379 33952 12434 33980
rect 13357 33983 13415 33989
rect 11379 33949 11391 33952
rect 11333 33943 11391 33949
rect 13357 33949 13369 33983
rect 13403 33949 13415 33983
rect 13357 33943 13415 33949
rect 13541 33983 13599 33989
rect 13541 33949 13553 33983
rect 13587 33980 13599 33983
rect 13814 33980 13820 33992
rect 13587 33952 13820 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 7984 33884 8156 33912
rect 8205 33915 8263 33921
rect 7984 33872 7990 33884
rect 8205 33881 8217 33915
rect 8251 33912 8263 33915
rect 9674 33912 9680 33924
rect 8251 33884 9680 33912
rect 8251 33881 8263 33884
rect 8205 33875 8263 33881
rect 9674 33872 9680 33884
rect 9732 33872 9738 33924
rect 7006 33804 7012 33856
rect 7064 33804 7070 33856
rect 9858 33804 9864 33856
rect 9916 33804 9922 33856
rect 10152 33844 10180 33943
rect 11054 33921 11060 33924
rect 11031 33915 11060 33921
rect 11031 33881 11043 33915
rect 11031 33875 11060 33881
rect 11054 33872 11060 33875
rect 11112 33872 11118 33924
rect 11146 33872 11152 33924
rect 11204 33872 11210 33924
rect 12158 33872 12164 33924
rect 12216 33872 12222 33924
rect 12894 33872 12900 33924
rect 12952 33872 12958 33924
rect 13372 33912 13400 33943
rect 13814 33940 13820 33952
rect 13872 33940 13878 33992
rect 16942 33940 16948 33992
rect 17000 33980 17006 33992
rect 19444 33989 19472 34156
rect 26697 34153 26709 34187
rect 26743 34184 26755 34187
rect 26786 34184 26792 34196
rect 26743 34156 26792 34184
rect 26743 34153 26755 34156
rect 26697 34147 26755 34153
rect 26786 34144 26792 34156
rect 26844 34144 26850 34196
rect 28169 34187 28227 34193
rect 28169 34153 28181 34187
rect 28215 34184 28227 34187
rect 28258 34184 28264 34196
rect 28215 34156 28264 34184
rect 28215 34153 28227 34156
rect 28169 34147 28227 34153
rect 28258 34144 28264 34156
rect 28316 34144 28322 34196
rect 28442 34144 28448 34196
rect 28500 34184 28506 34196
rect 28500 34156 30696 34184
rect 28500 34144 28506 34156
rect 21637 34119 21695 34125
rect 21637 34085 21649 34119
rect 21683 34116 21695 34119
rect 23014 34116 23020 34128
rect 21683 34088 23020 34116
rect 21683 34085 21695 34088
rect 21637 34079 21695 34085
rect 23014 34076 23020 34088
rect 23072 34076 23078 34128
rect 25866 34076 25872 34128
rect 25924 34116 25930 34128
rect 27982 34116 27988 34128
rect 25924 34088 27988 34116
rect 25924 34076 25930 34088
rect 27982 34076 27988 34088
rect 28040 34116 28046 34128
rect 30190 34116 30196 34128
rect 28040 34088 30196 34116
rect 28040 34076 28046 34088
rect 30190 34076 30196 34088
rect 30248 34076 30254 34128
rect 30668 34125 30696 34156
rect 31662 34144 31668 34196
rect 31720 34184 31726 34196
rect 31941 34187 31999 34193
rect 31941 34184 31953 34187
rect 31720 34156 31953 34184
rect 31720 34144 31726 34156
rect 31941 34153 31953 34156
rect 31987 34184 31999 34187
rect 32766 34184 32772 34196
rect 31987 34156 32772 34184
rect 31987 34153 31999 34156
rect 31941 34147 31999 34153
rect 32766 34144 32772 34156
rect 32824 34144 32830 34196
rect 33778 34144 33784 34196
rect 33836 34144 33842 34196
rect 35897 34187 35955 34193
rect 35897 34184 35909 34187
rect 34624 34156 35909 34184
rect 30653 34119 30711 34125
rect 30653 34085 30665 34119
rect 30699 34116 30711 34119
rect 31018 34116 31024 34128
rect 30699 34088 31024 34116
rect 30699 34085 30711 34088
rect 30653 34079 30711 34085
rect 31018 34076 31024 34088
rect 31076 34076 31082 34128
rect 34514 34116 34520 34128
rect 31128 34088 34520 34116
rect 20346 34048 20352 34060
rect 19536 34020 20352 34048
rect 19536 33992 19564 34020
rect 20346 34008 20352 34020
rect 20404 34008 20410 34060
rect 23106 34048 23112 34060
rect 22664 34020 23112 34048
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 17000 33952 17049 33980
rect 17000 33940 17006 33952
rect 17037 33949 17049 33952
rect 17083 33980 17095 33983
rect 19429 33983 19487 33989
rect 17083 33952 18368 33980
rect 17083 33949 17095 33952
rect 17037 33943 17095 33949
rect 14274 33912 14280 33924
rect 13372 33884 14280 33912
rect 14274 33872 14280 33884
rect 14332 33872 14338 33924
rect 16792 33915 16850 33921
rect 16792 33881 16804 33915
rect 16838 33912 16850 33915
rect 17402 33912 17408 33924
rect 16838 33884 17408 33912
rect 16838 33881 16850 33884
rect 16792 33875 16850 33881
rect 17402 33872 17408 33884
rect 17460 33872 17466 33924
rect 17494 33872 17500 33924
rect 17552 33872 17558 33924
rect 18340 33921 18368 33952
rect 19429 33949 19441 33983
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 19518 33940 19524 33992
rect 19576 33940 19582 33992
rect 19705 33983 19763 33989
rect 19705 33949 19717 33983
rect 19751 33980 19763 33983
rect 20254 33980 20260 33992
rect 19751 33952 20260 33980
rect 19751 33949 19763 33952
rect 19705 33943 19763 33949
rect 20254 33940 20260 33952
rect 20312 33940 20318 33992
rect 22664 33989 22692 34020
rect 23106 34008 23112 34020
rect 23164 34008 23170 34060
rect 25498 34048 25504 34060
rect 23400 34020 25504 34048
rect 21453 33983 21511 33989
rect 21453 33949 21465 33983
rect 21499 33949 21511 33983
rect 21453 33943 21511 33949
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33949 21603 33983
rect 21545 33943 21603 33949
rect 21729 33983 21787 33989
rect 21729 33949 21741 33983
rect 21775 33980 21787 33983
rect 22649 33983 22707 33989
rect 22649 33980 22661 33983
rect 21775 33952 22661 33980
rect 21775 33949 21787 33952
rect 21729 33943 21787 33949
rect 22649 33949 22661 33952
rect 22695 33949 22707 33983
rect 22649 33943 22707 33949
rect 18325 33915 18383 33921
rect 18325 33881 18337 33915
rect 18371 33912 18383 33915
rect 19242 33912 19248 33924
rect 18371 33884 19248 33912
rect 18371 33881 18383 33884
rect 18325 33875 18383 33881
rect 19242 33872 19248 33884
rect 19300 33872 19306 33924
rect 21468 33912 21496 33943
rect 19352 33884 21496 33912
rect 21560 33912 21588 33943
rect 23014 33940 23020 33992
rect 23072 33940 23078 33992
rect 23400 33989 23428 34020
rect 25498 34008 25504 34020
rect 25556 34008 25562 34060
rect 26605 34051 26663 34057
rect 26605 34017 26617 34051
rect 26651 34048 26663 34051
rect 27433 34051 27491 34057
rect 27433 34048 27445 34051
rect 26651 34020 27445 34048
rect 26651 34017 26663 34020
rect 26605 34011 26663 34017
rect 27433 34017 27445 34020
rect 27479 34017 27491 34051
rect 28994 34048 29000 34060
rect 27433 34011 27491 34017
rect 28000 34020 29000 34048
rect 23385 33983 23443 33989
rect 23385 33949 23397 33983
rect 23431 33949 23443 33983
rect 23385 33943 23443 33949
rect 23753 33983 23811 33989
rect 23753 33949 23765 33983
rect 23799 33949 23811 33983
rect 23753 33943 23811 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 24854 33980 24860 33992
rect 24811 33952 24860 33980
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 22922 33912 22928 33924
rect 21560 33884 22928 33912
rect 11330 33844 11336 33856
rect 10152 33816 11336 33844
rect 11330 33804 11336 33816
rect 11388 33804 11394 33856
rect 11517 33847 11575 33853
rect 11517 33813 11529 33847
rect 11563 33844 11575 33847
rect 15102 33844 15108 33856
rect 11563 33816 15108 33844
rect 11563 33813 11575 33816
rect 11517 33807 11575 33813
rect 15102 33804 15108 33816
rect 15160 33804 15166 33856
rect 15657 33847 15715 33853
rect 15657 33813 15669 33847
rect 15703 33844 15715 33847
rect 17862 33844 17868 33856
rect 15703 33816 17868 33844
rect 15703 33813 15715 33816
rect 15657 33807 15715 33813
rect 17862 33804 17868 33816
rect 17920 33844 17926 33856
rect 19352 33844 19380 33884
rect 22922 33872 22928 33884
rect 22980 33912 22986 33924
rect 23400 33912 23428 33943
rect 22980 33884 23428 33912
rect 23768 33912 23796 33943
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 26234 33940 26240 33992
rect 26292 33980 26298 33992
rect 26513 33983 26571 33989
rect 26513 33980 26525 33983
rect 26292 33952 26525 33980
rect 26292 33940 26298 33952
rect 26513 33949 26525 33952
rect 26559 33980 26571 33983
rect 26878 33980 26884 33992
rect 26559 33952 26884 33980
rect 26559 33949 26571 33952
rect 26513 33943 26571 33949
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 27154 33940 27160 33992
rect 27212 33980 27218 33992
rect 27341 33983 27399 33989
rect 27341 33980 27353 33983
rect 27212 33952 27353 33980
rect 27212 33940 27218 33952
rect 27341 33949 27353 33952
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 27522 33940 27528 33992
rect 27580 33940 27586 33992
rect 28000 33989 28028 34020
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 29270 34008 29276 34060
rect 29328 34048 29334 34060
rect 30101 34051 30159 34057
rect 30101 34048 30113 34051
rect 29328 34020 30113 34048
rect 29328 34008 29334 34020
rect 30101 34017 30113 34020
rect 30147 34017 30159 34051
rect 30101 34011 30159 34017
rect 27985 33983 28043 33989
rect 27985 33949 27997 33983
rect 28031 33949 28043 33983
rect 27985 33943 28043 33949
rect 23842 33912 23848 33924
rect 23768 33884 23848 33912
rect 22980 33872 22986 33884
rect 23842 33872 23848 33884
rect 23900 33912 23906 33924
rect 25777 33915 25835 33921
rect 25777 33912 25789 33915
rect 23900 33884 25789 33912
rect 23900 33872 23906 33884
rect 25777 33881 25789 33884
rect 25823 33912 25835 33915
rect 25958 33912 25964 33924
rect 25823 33884 25964 33912
rect 25823 33881 25835 33884
rect 25777 33875 25835 33881
rect 25958 33872 25964 33884
rect 26016 33872 26022 33924
rect 26050 33872 26056 33924
rect 26108 33912 26114 33924
rect 28000 33912 28028 33943
rect 28074 33940 28080 33992
rect 28132 33980 28138 33992
rect 28169 33983 28227 33989
rect 28169 33980 28181 33983
rect 28132 33952 28181 33980
rect 28132 33940 28138 33952
rect 28169 33949 28181 33952
rect 28215 33949 28227 33983
rect 28169 33943 28227 33949
rect 29914 33940 29920 33992
rect 29972 33940 29978 33992
rect 30558 33940 30564 33992
rect 30616 33940 30622 33992
rect 30834 33940 30840 33992
rect 30892 33940 30898 33992
rect 31128 33980 31156 34088
rect 33686 34048 33692 34060
rect 32784 34020 33692 34048
rect 30944 33952 31156 33980
rect 30944 33912 30972 33952
rect 31754 33940 31760 33992
rect 31812 33980 31818 33992
rect 32784 33989 32812 34020
rect 33686 34008 33692 34020
rect 33744 34008 33750 34060
rect 32585 33983 32643 33989
rect 32585 33980 32597 33983
rect 31812 33952 32597 33980
rect 31812 33940 31818 33952
rect 32585 33949 32597 33952
rect 32631 33949 32643 33983
rect 32585 33943 32643 33949
rect 32769 33983 32827 33989
rect 32769 33949 32781 33983
rect 32815 33949 32827 33983
rect 32769 33943 32827 33949
rect 32861 33983 32919 33989
rect 32861 33949 32873 33983
rect 32907 33949 32919 33983
rect 32861 33943 32919 33949
rect 32953 33983 33011 33989
rect 32953 33949 32965 33983
rect 32999 33980 33011 33983
rect 33796 33980 33824 34088
rect 34514 34076 34520 34088
rect 34572 34076 34578 34128
rect 34624 34048 34652 34156
rect 35897 34153 35909 34156
rect 35943 34184 35955 34187
rect 35986 34184 35992 34196
rect 35943 34156 35992 34184
rect 35943 34153 35955 34156
rect 35897 34147 35955 34153
rect 35986 34144 35992 34156
rect 36044 34184 36050 34196
rect 36630 34184 36636 34196
rect 36044 34156 36636 34184
rect 36044 34144 36050 34156
rect 36630 34144 36636 34156
rect 36688 34144 36694 34196
rect 34072 34020 34652 34048
rect 32999 33952 33824 33980
rect 32999 33949 33011 33952
rect 32953 33943 33011 33949
rect 31478 33912 31484 33924
rect 26108 33884 28028 33912
rect 28092 33884 30972 33912
rect 31036 33884 31484 33912
rect 26108 33872 26114 33884
rect 17920 33816 19380 33844
rect 19889 33847 19947 33853
rect 17920 33804 17926 33816
rect 19889 33813 19901 33847
rect 19935 33844 19947 33847
rect 19978 33844 19984 33856
rect 19935 33816 19984 33844
rect 19935 33813 19947 33816
rect 19889 33807 19947 33813
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 21913 33847 21971 33853
rect 21913 33813 21925 33847
rect 21959 33844 21971 33847
rect 22278 33844 22284 33856
rect 21959 33816 22284 33844
rect 21959 33813 21971 33816
rect 21913 33807 21971 33813
rect 22278 33804 22284 33816
rect 22336 33804 22342 33856
rect 22462 33804 22468 33856
rect 22520 33804 22526 33856
rect 26878 33804 26884 33856
rect 26936 33804 26942 33856
rect 27522 33804 27528 33856
rect 27580 33844 27586 33856
rect 27890 33844 27896 33856
rect 27580 33816 27896 33844
rect 27580 33804 27586 33816
rect 27890 33804 27896 33816
rect 27948 33844 27954 33856
rect 28092 33844 28120 33884
rect 27948 33816 28120 33844
rect 29733 33847 29791 33853
rect 27948 33804 27954 33816
rect 29733 33813 29745 33847
rect 29779 33844 29791 33847
rect 30098 33844 30104 33856
rect 29779 33816 30104 33844
rect 29779 33813 29791 33816
rect 29733 33807 29791 33813
rect 30098 33804 30104 33816
rect 30156 33804 30162 33856
rect 30558 33804 30564 33856
rect 30616 33844 30622 33856
rect 31036 33853 31064 33884
rect 31478 33872 31484 33884
rect 31536 33912 31542 33924
rect 32125 33915 32183 33921
rect 32125 33912 32137 33915
rect 31536 33884 32137 33912
rect 31536 33872 31542 33884
rect 32125 33881 32137 33884
rect 32171 33881 32183 33915
rect 32125 33875 32183 33881
rect 32398 33872 32404 33924
rect 32456 33912 32462 33924
rect 32876 33912 32904 33943
rect 33962 33940 33968 33992
rect 34020 33940 34026 33992
rect 34072 33989 34100 34020
rect 35434 34008 35440 34060
rect 35492 34048 35498 34060
rect 35805 34051 35863 34057
rect 35805 34048 35817 34051
rect 35492 34020 35817 34048
rect 35492 34008 35498 34020
rect 35805 34017 35817 34020
rect 35851 34017 35863 34051
rect 35805 34011 35863 34017
rect 41782 34008 41788 34060
rect 41840 34048 41846 34060
rect 41877 34051 41935 34057
rect 41877 34048 41889 34051
rect 41840 34020 41889 34048
rect 41840 34008 41846 34020
rect 41877 34017 41889 34020
rect 41923 34017 41935 34051
rect 41877 34011 41935 34017
rect 34057 33983 34115 33989
rect 34057 33949 34069 33983
rect 34103 33949 34115 33983
rect 34057 33943 34115 33949
rect 34146 33940 34152 33992
rect 34204 33980 34210 33992
rect 35069 33983 35127 33989
rect 35069 33980 35081 33983
rect 34204 33952 35081 33980
rect 34204 33940 34210 33952
rect 35069 33949 35081 33952
rect 35115 33980 35127 33983
rect 35115 33952 35388 33980
rect 35115 33949 35127 33952
rect 35069 33943 35127 33949
rect 32456 33884 32904 33912
rect 33781 33915 33839 33921
rect 32456 33872 32462 33884
rect 33781 33881 33793 33915
rect 33827 33912 33839 33915
rect 34422 33912 34428 33924
rect 33827 33884 34428 33912
rect 33827 33881 33839 33884
rect 33781 33875 33839 33881
rect 34422 33872 34428 33884
rect 34480 33872 34486 33924
rect 34885 33915 34943 33921
rect 34885 33881 34897 33915
rect 34931 33881 34943 33915
rect 34885 33875 34943 33881
rect 31021 33847 31079 33853
rect 31021 33844 31033 33847
rect 30616 33816 31033 33844
rect 30616 33804 30622 33816
rect 31021 33813 31033 33816
rect 31067 33813 31079 33847
rect 31021 33807 31079 33813
rect 31386 33804 31392 33856
rect 31444 33844 31450 33856
rect 31938 33853 31944 33856
rect 31757 33847 31815 33853
rect 31757 33844 31769 33847
rect 31444 33816 31769 33844
rect 31444 33804 31450 33816
rect 31757 33813 31769 33816
rect 31803 33813 31815 33847
rect 31757 33807 31815 33813
rect 31925 33847 31944 33853
rect 31925 33813 31937 33847
rect 31925 33807 31944 33813
rect 31938 33804 31944 33807
rect 31996 33804 32002 33856
rect 33229 33847 33287 33853
rect 33229 33813 33241 33847
rect 33275 33844 33287 33847
rect 33594 33844 33600 33856
rect 33275 33816 33600 33844
rect 33275 33813 33287 33816
rect 33229 33807 33287 33813
rect 33594 33804 33600 33816
rect 33652 33804 33658 33856
rect 34241 33847 34299 33853
rect 34241 33813 34253 33847
rect 34287 33844 34299 33847
rect 34514 33844 34520 33856
rect 34287 33816 34520 33844
rect 34287 33813 34299 33816
rect 34241 33807 34299 33813
rect 34514 33804 34520 33816
rect 34572 33804 34578 33856
rect 34900 33844 34928 33875
rect 35250 33872 35256 33924
rect 35308 33872 35314 33924
rect 35360 33912 35388 33952
rect 35710 33940 35716 33992
rect 35768 33940 35774 33992
rect 37550 33912 37556 33924
rect 35360 33884 37556 33912
rect 37550 33872 37556 33884
rect 37608 33872 37614 33924
rect 42144 33915 42202 33921
rect 42144 33881 42156 33915
rect 42190 33912 42202 33915
rect 42610 33912 42616 33924
rect 42190 33884 42616 33912
rect 42190 33881 42202 33884
rect 42144 33875 42202 33881
rect 42610 33872 42616 33884
rect 42668 33872 42674 33924
rect 35710 33844 35716 33856
rect 34900 33816 35716 33844
rect 35710 33804 35716 33816
rect 35768 33804 35774 33856
rect 35802 33804 35808 33856
rect 35860 33844 35866 33856
rect 36081 33847 36139 33853
rect 36081 33844 36093 33847
rect 35860 33816 36093 33844
rect 35860 33804 35866 33816
rect 36081 33813 36093 33816
rect 36127 33813 36139 33847
rect 36081 33807 36139 33813
rect 42978 33804 42984 33856
rect 43036 33844 43042 33856
rect 43257 33847 43315 33853
rect 43257 33844 43269 33847
rect 43036 33816 43269 33844
rect 43036 33804 43042 33816
rect 43257 33813 43269 33816
rect 43303 33813 43315 33847
rect 43257 33807 43315 33813
rect 1104 33754 43884 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 43884 33754
rect 1104 33680 43884 33702
rect 7101 33643 7159 33649
rect 7101 33609 7113 33643
rect 7147 33640 7159 33643
rect 8110 33640 8116 33652
rect 7147 33612 8116 33640
rect 7147 33609 7159 33612
rect 7101 33603 7159 33609
rect 8110 33600 8116 33612
rect 8168 33600 8174 33652
rect 8941 33643 8999 33649
rect 8941 33609 8953 33643
rect 8987 33640 8999 33643
rect 10226 33640 10232 33652
rect 8987 33612 10232 33640
rect 8987 33609 8999 33612
rect 8941 33603 8999 33609
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 20162 33600 20168 33652
rect 20220 33640 20226 33652
rect 25958 33640 25964 33652
rect 20220 33612 25964 33640
rect 20220 33600 20226 33612
rect 25958 33600 25964 33612
rect 26016 33600 26022 33652
rect 26053 33643 26111 33649
rect 26053 33609 26065 33643
rect 26099 33640 26111 33643
rect 26418 33640 26424 33652
rect 26099 33612 26424 33640
rect 26099 33609 26111 33612
rect 26053 33603 26111 33609
rect 26418 33600 26424 33612
rect 26476 33600 26482 33652
rect 27985 33643 28043 33649
rect 27985 33609 27997 33643
rect 28031 33609 28043 33643
rect 27985 33603 28043 33609
rect 6362 33532 6368 33584
rect 6420 33572 6426 33584
rect 6420 33544 7144 33572
rect 6420 33532 6426 33544
rect 5077 33507 5135 33513
rect 5077 33473 5089 33507
rect 5123 33504 5135 33507
rect 6270 33504 6276 33516
rect 5123 33476 6276 33504
rect 5123 33473 5135 33476
rect 5077 33467 5135 33473
rect 6270 33464 6276 33476
rect 6328 33464 6334 33516
rect 6822 33464 6828 33516
rect 6880 33464 6886 33516
rect 6917 33507 6975 33513
rect 6917 33473 6929 33507
rect 6963 33504 6975 33507
rect 7006 33504 7012 33516
rect 6963 33476 7012 33504
rect 6963 33473 6975 33476
rect 6917 33467 6975 33473
rect 7006 33464 7012 33476
rect 7064 33464 7070 33516
rect 5350 33396 5356 33448
rect 5408 33396 5414 33448
rect 6638 33396 6644 33448
rect 6696 33396 6702 33448
rect 6733 33439 6791 33445
rect 6733 33405 6745 33439
rect 6779 33405 6791 33439
rect 7116 33436 7144 33544
rect 9490 33532 9496 33584
rect 9548 33572 9554 33584
rect 9953 33575 10011 33581
rect 9953 33572 9965 33575
rect 9548 33544 9965 33572
rect 9548 33532 9554 33544
rect 9953 33541 9965 33544
rect 9999 33541 10011 33575
rect 9953 33535 10011 33541
rect 10686 33532 10692 33584
rect 10744 33572 10750 33584
rect 10744 33544 12020 33572
rect 10744 33532 10750 33544
rect 9306 33464 9312 33516
rect 9364 33504 9370 33516
rect 9766 33504 9772 33516
rect 9364 33476 9772 33504
rect 9364 33464 9370 33476
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 10045 33507 10103 33513
rect 10045 33473 10057 33507
rect 10091 33504 10103 33507
rect 10410 33504 10416 33516
rect 10091 33476 10416 33504
rect 10091 33473 10103 33476
rect 10045 33467 10103 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10597 33507 10655 33513
rect 10597 33473 10609 33507
rect 10643 33504 10655 33507
rect 10778 33504 10784 33516
rect 10643 33476 10784 33504
rect 10643 33473 10655 33476
rect 10597 33467 10655 33473
rect 10778 33464 10784 33476
rect 10836 33464 10842 33516
rect 10873 33507 10931 33513
rect 10873 33473 10885 33507
rect 10919 33504 10931 33507
rect 10962 33504 10968 33516
rect 10919 33476 10968 33504
rect 10919 33473 10931 33476
rect 10873 33467 10931 33473
rect 10962 33464 10968 33476
rect 11020 33464 11026 33516
rect 11992 33504 12020 33544
rect 12066 33532 12072 33584
rect 12124 33532 12130 33584
rect 12894 33532 12900 33584
rect 12952 33572 12958 33584
rect 17494 33572 17500 33584
rect 12952 33544 17500 33572
rect 12952 33532 12958 33544
rect 17494 33532 17500 33544
rect 17552 33532 17558 33584
rect 19604 33575 19662 33581
rect 19604 33541 19616 33575
rect 19650 33572 19662 33575
rect 19978 33572 19984 33584
rect 19650 33544 19984 33572
rect 19650 33541 19662 33544
rect 19604 33535 19662 33541
rect 19978 33532 19984 33544
rect 20036 33532 20042 33584
rect 23842 33572 23848 33584
rect 22112 33544 23848 33572
rect 13538 33504 13544 33516
rect 11992 33476 13544 33504
rect 13538 33464 13544 33476
rect 13596 33464 13602 33516
rect 13817 33507 13875 33513
rect 13817 33473 13829 33507
rect 13863 33504 13875 33507
rect 14182 33504 14188 33516
rect 13863 33476 14188 33504
rect 13863 33473 13875 33476
rect 13817 33467 13875 33473
rect 14182 33464 14188 33476
rect 14240 33464 14246 33516
rect 14277 33507 14335 33513
rect 14277 33473 14289 33507
rect 14323 33473 14335 33507
rect 14277 33467 14335 33473
rect 14461 33507 14519 33513
rect 14461 33473 14473 33507
rect 14507 33504 14519 33507
rect 14550 33504 14556 33516
rect 14507 33476 14556 33504
rect 14507 33473 14519 33476
rect 14461 33467 14519 33473
rect 7116 33408 12434 33436
rect 6733 33399 6791 33405
rect 6748 33368 6776 33399
rect 7558 33368 7564 33380
rect 6748 33340 7564 33368
rect 7558 33328 7564 33340
rect 7616 33328 7622 33380
rect 7926 33328 7932 33380
rect 7984 33368 7990 33380
rect 10781 33371 10839 33377
rect 10781 33368 10793 33371
rect 7984 33340 9076 33368
rect 7984 33328 7990 33340
rect 4890 33260 4896 33312
rect 4948 33260 4954 33312
rect 5258 33260 5264 33312
rect 5316 33260 5322 33312
rect 8754 33260 8760 33312
rect 8812 33260 8818 33312
rect 8846 33260 8852 33312
rect 8904 33300 8910 33312
rect 8941 33303 8999 33309
rect 8941 33300 8953 33303
rect 8904 33272 8953 33300
rect 8904 33260 8910 33272
rect 8941 33269 8953 33272
rect 8987 33269 8999 33303
rect 9048 33300 9076 33340
rect 9407 33340 10793 33368
rect 9407 33300 9435 33340
rect 10781 33337 10793 33340
rect 10827 33337 10839 33371
rect 12406 33368 12434 33408
rect 13354 33396 13360 33448
rect 13412 33436 13418 33448
rect 13633 33439 13691 33445
rect 13633 33436 13645 33439
rect 13412 33408 13645 33436
rect 13412 33396 13418 33408
rect 13633 33405 13645 33408
rect 13679 33405 13691 33439
rect 13633 33399 13691 33405
rect 13722 33396 13728 33448
rect 13780 33436 13786 33448
rect 14292 33436 14320 33467
rect 14550 33464 14556 33476
rect 14608 33464 14614 33516
rect 16853 33507 16911 33513
rect 16853 33473 16865 33507
rect 16899 33504 16911 33507
rect 16942 33504 16948 33516
rect 16899 33476 16948 33504
rect 16899 33473 16911 33476
rect 16853 33467 16911 33473
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 17126 33513 17132 33516
rect 17120 33467 17132 33513
rect 17126 33464 17132 33467
rect 17184 33464 17190 33516
rect 22112 33513 22140 33544
rect 23842 33532 23848 33544
rect 23900 33532 23906 33584
rect 24949 33575 25007 33581
rect 24949 33541 24961 33575
rect 24995 33572 25007 33575
rect 25498 33572 25504 33584
rect 24995 33544 25504 33572
rect 24995 33541 25007 33544
rect 24949 33535 25007 33541
rect 25498 33532 25504 33544
rect 25556 33532 25562 33584
rect 26145 33575 26203 33581
rect 26145 33541 26157 33575
rect 26191 33572 26203 33575
rect 26786 33572 26792 33584
rect 26191 33544 26792 33572
rect 26191 33541 26203 33544
rect 26145 33535 26203 33541
rect 26786 33532 26792 33544
rect 26844 33532 26850 33584
rect 26878 33532 26884 33584
rect 26936 33572 26942 33584
rect 27525 33575 27583 33581
rect 27525 33572 27537 33575
rect 26936 33544 27537 33572
rect 26936 33532 26942 33544
rect 27525 33541 27537 33544
rect 27571 33541 27583 33575
rect 28000 33572 28028 33603
rect 28442 33600 28448 33652
rect 28500 33640 28506 33652
rect 30650 33640 30656 33652
rect 28500 33612 30656 33640
rect 28500 33600 28506 33612
rect 30650 33600 30656 33612
rect 30708 33640 30714 33652
rect 31110 33640 31116 33652
rect 30708 33612 31116 33640
rect 30708 33600 30714 33612
rect 31110 33600 31116 33612
rect 31168 33600 31174 33652
rect 31754 33600 31760 33652
rect 31812 33600 31818 33652
rect 32950 33600 32956 33652
rect 33008 33640 33014 33652
rect 36446 33640 36452 33652
rect 33008 33612 36452 33640
rect 33008 33600 33014 33612
rect 36446 33600 36452 33612
rect 36504 33600 36510 33652
rect 37090 33600 37096 33652
rect 37148 33640 37154 33652
rect 37148 33612 39436 33640
rect 37148 33600 37154 33612
rect 32490 33572 32496 33584
rect 28000 33544 32496 33572
rect 27525 33535 27583 33541
rect 32490 33532 32496 33544
rect 32548 33532 32554 33584
rect 33042 33532 33048 33584
rect 33100 33572 33106 33584
rect 33137 33575 33195 33581
rect 33137 33572 33149 33575
rect 33100 33544 33149 33572
rect 33100 33532 33106 33544
rect 33137 33541 33149 33544
rect 33183 33541 33195 33575
rect 33137 33535 33195 33541
rect 34790 33532 34796 33584
rect 34848 33572 34854 33584
rect 35526 33572 35532 33584
rect 34848 33544 35532 33572
rect 34848 33532 34854 33544
rect 35526 33532 35532 33544
rect 35584 33532 35590 33584
rect 36170 33532 36176 33584
rect 36228 33572 36234 33584
rect 36228 33544 39160 33572
rect 36228 33532 36234 33544
rect 22097 33507 22155 33513
rect 22097 33473 22109 33507
rect 22143 33473 22155 33507
rect 22097 33467 22155 33473
rect 22189 33507 22247 33513
rect 22189 33473 22201 33507
rect 22235 33473 22247 33507
rect 22189 33467 22247 33473
rect 13780 33408 14320 33436
rect 13780 33396 13786 33408
rect 19242 33396 19248 33448
rect 19300 33436 19306 33448
rect 19337 33439 19395 33445
rect 19337 33436 19349 33439
rect 19300 33408 19349 33436
rect 19300 33396 19306 33408
rect 19337 33405 19349 33408
rect 19383 33405 19395 33439
rect 19337 33399 19395 33405
rect 16482 33368 16488 33380
rect 12406 33340 16488 33368
rect 10781 33331 10839 33337
rect 16482 33328 16488 33340
rect 16540 33328 16546 33380
rect 20622 33328 20628 33380
rect 20680 33368 20686 33380
rect 20717 33371 20775 33377
rect 20717 33368 20729 33371
rect 20680 33340 20729 33368
rect 20680 33328 20686 33340
rect 20717 33337 20729 33340
rect 20763 33368 20775 33371
rect 22204 33368 22232 33467
rect 22278 33464 22284 33516
rect 22336 33504 22342 33516
rect 22557 33507 22615 33513
rect 22557 33504 22569 33507
rect 22336 33476 22569 33504
rect 22336 33464 22342 33476
rect 22557 33473 22569 33476
rect 22603 33473 22615 33507
rect 22557 33467 22615 33473
rect 24302 33464 24308 33516
rect 24360 33464 24366 33516
rect 24765 33507 24823 33513
rect 24765 33473 24777 33507
rect 24811 33504 24823 33507
rect 24854 33504 24860 33516
rect 24811 33476 24860 33504
rect 24811 33473 24823 33476
rect 24765 33467 24823 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 25406 33464 25412 33516
rect 25464 33464 25470 33516
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33473 26019 33507
rect 25961 33467 26019 33473
rect 22462 33396 22468 33448
rect 22520 33396 22526 33448
rect 23658 33396 23664 33448
rect 23716 33436 23722 33448
rect 25593 33439 25651 33445
rect 25593 33436 25605 33439
rect 23716 33408 25605 33436
rect 23716 33396 23722 33408
rect 25593 33405 25605 33408
rect 25639 33405 25651 33439
rect 25976 33436 26004 33467
rect 26602 33464 26608 33516
rect 26660 33504 26666 33516
rect 27246 33504 27252 33516
rect 26660 33476 27252 33504
rect 26660 33464 26666 33476
rect 27246 33464 27252 33476
rect 27304 33504 27310 33516
rect 27794 33507 27852 33513
rect 27794 33504 27806 33507
rect 27304 33476 27806 33504
rect 27304 33464 27310 33476
rect 27794 33473 27806 33476
rect 27840 33473 27852 33507
rect 27794 33467 27852 33473
rect 28534 33464 28540 33516
rect 28592 33504 28598 33516
rect 28629 33507 28687 33513
rect 28629 33504 28641 33507
rect 28592 33476 28641 33504
rect 28592 33464 28598 33476
rect 28629 33473 28641 33476
rect 28675 33473 28687 33507
rect 28629 33467 28687 33473
rect 28902 33464 28908 33516
rect 28960 33464 28966 33516
rect 30285 33507 30343 33513
rect 30285 33504 30297 33507
rect 30024 33476 30297 33504
rect 27522 33436 27528 33448
rect 25976 33408 27528 33436
rect 25593 33399 25651 33405
rect 27522 33396 27528 33408
rect 27580 33396 27586 33448
rect 27614 33396 27620 33448
rect 27672 33396 27678 33448
rect 28721 33439 28779 33445
rect 28721 33436 28733 33439
rect 27724 33408 28733 33436
rect 20763 33340 22232 33368
rect 20763 33337 20775 33340
rect 20717 33331 20775 33337
rect 22370 33328 22376 33380
rect 22428 33368 22434 33380
rect 27724 33368 27752 33408
rect 28721 33405 28733 33408
rect 28767 33405 28779 33439
rect 28721 33399 28779 33405
rect 28810 33396 28816 33448
rect 28868 33436 28874 33448
rect 30024 33436 30052 33476
rect 30285 33473 30297 33476
rect 30331 33504 30343 33507
rect 30558 33504 30564 33516
rect 30331 33476 30564 33504
rect 30331 33473 30343 33476
rect 30285 33467 30343 33473
rect 30558 33464 30564 33476
rect 30616 33464 30622 33516
rect 30653 33507 30711 33513
rect 30653 33473 30665 33507
rect 30699 33504 30711 33507
rect 30742 33504 30748 33516
rect 30699 33476 30748 33504
rect 30699 33473 30711 33476
rect 30653 33467 30711 33473
rect 30742 33464 30748 33476
rect 30800 33464 30806 33516
rect 31113 33507 31171 33513
rect 31113 33473 31125 33507
rect 31159 33504 31171 33507
rect 31202 33504 31208 33516
rect 31159 33476 31208 33504
rect 31159 33473 31171 33476
rect 31113 33467 31171 33473
rect 31202 33464 31208 33476
rect 31260 33464 31266 33516
rect 31294 33464 31300 33516
rect 31352 33464 31358 33516
rect 31386 33464 31392 33516
rect 31444 33464 31450 33516
rect 31481 33507 31539 33513
rect 31481 33473 31493 33507
rect 31527 33504 31539 33507
rect 31570 33504 31576 33516
rect 31527 33476 31576 33504
rect 31527 33473 31539 33476
rect 31481 33467 31539 33473
rect 31570 33464 31576 33476
rect 31628 33504 31634 33516
rect 36469 33507 36527 33513
rect 31628 33476 33088 33504
rect 31628 33464 31634 33476
rect 28868 33408 30052 33436
rect 28868 33396 28874 33408
rect 30190 33396 30196 33448
rect 30248 33396 30254 33448
rect 33060 33436 33088 33476
rect 36469 33473 36481 33507
rect 36515 33504 36527 33507
rect 37734 33504 37740 33516
rect 36515 33476 37740 33504
rect 36515 33473 36527 33476
rect 36469 33467 36527 33473
rect 37734 33464 37740 33476
rect 37792 33464 37798 33516
rect 39132 33513 39160 33544
rect 39298 33532 39304 33584
rect 39356 33532 39362 33584
rect 39408 33581 39436 33612
rect 42610 33600 42616 33652
rect 42668 33600 42674 33652
rect 39393 33575 39451 33581
rect 39393 33541 39405 33575
rect 39439 33541 39451 33575
rect 39393 33535 39451 33541
rect 40310 33532 40316 33584
rect 40368 33572 40374 33584
rect 40773 33575 40831 33581
rect 40773 33572 40785 33575
rect 40368 33544 40785 33572
rect 40368 33532 40374 33544
rect 40773 33541 40785 33544
rect 40819 33541 40831 33575
rect 42978 33572 42984 33584
rect 40773 33535 40831 33541
rect 41386 33544 42984 33572
rect 39117 33507 39175 33513
rect 39117 33473 39129 33507
rect 39163 33473 39175 33507
rect 39117 33467 39175 33473
rect 33410 33436 33416 33448
rect 33060 33408 33416 33436
rect 33410 33396 33416 33408
rect 33468 33396 33474 33448
rect 36722 33396 36728 33448
rect 36780 33396 36786 33448
rect 38654 33396 38660 33448
rect 38712 33436 38718 33448
rect 39316 33436 39344 33532
rect 39485 33507 39543 33513
rect 39485 33473 39497 33507
rect 39531 33473 39543 33507
rect 40405 33507 40463 33513
rect 40405 33504 40417 33507
rect 39485 33467 39543 33473
rect 39684 33476 40417 33504
rect 38712 33408 39344 33436
rect 38712 33396 38718 33408
rect 39390 33396 39396 33448
rect 39448 33436 39454 33448
rect 39500 33436 39528 33467
rect 39448 33408 39528 33436
rect 39448 33396 39454 33408
rect 22428 33340 27752 33368
rect 22428 33328 22434 33340
rect 28442 33328 28448 33380
rect 28500 33328 28506 33380
rect 31662 33368 31668 33380
rect 28552 33340 31668 33368
rect 9048 33272 9435 33300
rect 8941 33263 8999 33269
rect 9766 33260 9772 33312
rect 9824 33260 9830 33312
rect 12986 33260 12992 33312
rect 13044 33300 13050 33312
rect 13357 33303 13415 33309
rect 13357 33300 13369 33303
rect 13044 33272 13369 33300
rect 13044 33260 13050 33272
rect 13357 33269 13369 33272
rect 13403 33269 13415 33303
rect 13357 33263 13415 33269
rect 13538 33260 13544 33312
rect 13596 33260 13602 33312
rect 13906 33260 13912 33312
rect 13964 33300 13970 33312
rect 14277 33303 14335 33309
rect 14277 33300 14289 33303
rect 13964 33272 14289 33300
rect 13964 33260 13970 33272
rect 14277 33269 14289 33272
rect 14323 33269 14335 33303
rect 14277 33263 14335 33269
rect 18233 33303 18291 33309
rect 18233 33269 18245 33303
rect 18279 33300 18291 33303
rect 20070 33300 20076 33312
rect 18279 33272 20076 33300
rect 18279 33269 18291 33272
rect 18233 33263 18291 33269
rect 20070 33260 20076 33272
rect 20128 33260 20134 33312
rect 22278 33260 22284 33312
rect 22336 33300 22342 33312
rect 23109 33303 23167 33309
rect 23109 33300 23121 33303
rect 22336 33272 23121 33300
rect 22336 33260 22342 33272
rect 23109 33269 23121 33272
rect 23155 33269 23167 33303
rect 23109 33263 23167 33269
rect 24854 33260 24860 33312
rect 24912 33300 24918 33312
rect 27154 33300 27160 33312
rect 24912 33272 27160 33300
rect 24912 33260 24918 33272
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 27798 33260 27804 33312
rect 27856 33260 27862 33312
rect 28074 33260 28080 33312
rect 28132 33300 28138 33312
rect 28552 33300 28580 33340
rect 31662 33328 31668 33340
rect 31720 33328 31726 33380
rect 39684 33377 39712 33476
rect 40405 33473 40417 33476
rect 40451 33473 40463 33507
rect 40405 33467 40463 33473
rect 40498 33507 40556 33513
rect 40498 33473 40510 33507
rect 40544 33473 40556 33507
rect 40498 33467 40556 33473
rect 40512 33436 40540 33467
rect 40586 33464 40592 33516
rect 40644 33504 40650 33516
rect 40681 33507 40739 33513
rect 40681 33504 40693 33507
rect 40644 33476 40693 33504
rect 40644 33464 40650 33476
rect 40681 33473 40693 33476
rect 40727 33473 40739 33507
rect 40681 33467 40739 33473
rect 40911 33507 40969 33513
rect 40911 33473 40923 33507
rect 40957 33504 40969 33507
rect 41138 33504 41144 33516
rect 40957 33476 41144 33504
rect 40957 33473 40969 33476
rect 40911 33467 40969 33473
rect 41138 33464 41144 33476
rect 41196 33464 41202 33516
rect 41386 33436 41414 33544
rect 42978 33532 42984 33544
rect 43036 33532 43042 33584
rect 40512 33408 41414 33436
rect 43073 33439 43131 33445
rect 39669 33371 39727 33377
rect 39669 33337 39681 33371
rect 39715 33337 39727 33371
rect 39669 33331 39727 33337
rect 28132 33272 28580 33300
rect 28132 33260 28138 33272
rect 28626 33260 28632 33312
rect 28684 33260 28690 33312
rect 30561 33303 30619 33309
rect 30561 33269 30573 33303
rect 30607 33300 30619 33303
rect 30742 33300 30748 33312
rect 30607 33272 30748 33300
rect 30607 33269 30619 33272
rect 30561 33263 30619 33269
rect 30742 33260 30748 33272
rect 30800 33260 30806 33312
rect 34422 33260 34428 33312
rect 34480 33260 34486 33312
rect 35342 33260 35348 33312
rect 35400 33260 35406 33312
rect 36446 33260 36452 33312
rect 36504 33300 36510 33312
rect 40512 33300 40540 33408
rect 43073 33405 43085 33439
rect 43119 33405 43131 33439
rect 43073 33399 43131 33405
rect 41049 33371 41107 33377
rect 41049 33337 41061 33371
rect 41095 33368 41107 33371
rect 42886 33368 42892 33380
rect 41095 33340 42892 33368
rect 41095 33337 41107 33340
rect 41049 33331 41107 33337
rect 42886 33328 42892 33340
rect 42944 33368 42950 33380
rect 43088 33368 43116 33399
rect 43254 33396 43260 33448
rect 43312 33396 43318 33448
rect 42944 33340 43116 33368
rect 42944 33328 42950 33340
rect 36504 33272 40540 33300
rect 36504 33260 36510 33272
rect 1104 33210 43884 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 43884 33210
rect 1104 33136 43884 33158
rect 6270 33056 6276 33108
rect 6328 33056 6334 33108
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 7745 33099 7803 33105
rect 7745 33096 7757 33099
rect 7616 33068 7757 33096
rect 7616 33056 7622 33068
rect 7745 33065 7757 33068
rect 7791 33065 7803 33099
rect 7745 33059 7803 33065
rect 7834 33056 7840 33108
rect 7892 33056 7898 33108
rect 7929 33099 7987 33105
rect 7929 33065 7941 33099
rect 7975 33096 7987 33099
rect 9306 33096 9312 33108
rect 7975 33068 9312 33096
rect 7975 33065 7987 33068
rect 7929 33059 7987 33065
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 10410 33056 10416 33108
rect 10468 33096 10474 33108
rect 10594 33096 10600 33108
rect 10468 33068 10600 33096
rect 10468 33056 10474 33068
rect 10594 33056 10600 33068
rect 10652 33096 10658 33108
rect 10781 33099 10839 33105
rect 10781 33096 10793 33099
rect 10652 33068 10793 33096
rect 10652 33056 10658 33068
rect 10781 33065 10793 33068
rect 10827 33065 10839 33099
rect 10781 33059 10839 33065
rect 10962 33056 10968 33108
rect 11020 33056 11026 33108
rect 12250 33056 12256 33108
rect 12308 33056 12314 33108
rect 12406 33068 17264 33096
rect 5350 32988 5356 33040
rect 5408 33028 5414 33040
rect 5445 33031 5503 33037
rect 5445 33028 5457 33031
rect 5408 33000 5457 33028
rect 5408 32988 5414 33000
rect 5445 32997 5457 33000
rect 5491 33028 5503 33031
rect 12406 33028 12434 33068
rect 5491 33000 12434 33028
rect 17236 33028 17264 33068
rect 17402 33056 17408 33108
rect 17460 33096 17466 33108
rect 17497 33099 17555 33105
rect 17497 33096 17509 33099
rect 17460 33068 17509 33096
rect 17460 33056 17466 33068
rect 17497 33065 17509 33068
rect 17543 33065 17555 33099
rect 17497 33059 17555 33065
rect 18046 33056 18052 33108
rect 18104 33096 18110 33108
rect 18690 33096 18696 33108
rect 18104 33068 18696 33096
rect 18104 33056 18110 33068
rect 18690 33056 18696 33068
rect 18748 33096 18754 33108
rect 19150 33096 19156 33108
rect 18748 33068 19156 33096
rect 18748 33056 18754 33068
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 19978 33096 19984 33108
rect 19392 33068 19984 33096
rect 19392 33056 19398 33068
rect 19978 33056 19984 33068
rect 20036 33056 20042 33108
rect 21358 33056 21364 33108
rect 21416 33096 21422 33108
rect 21416 33068 22232 33096
rect 21416 33056 21422 33068
rect 22204 33028 22232 33068
rect 23198 33056 23204 33108
rect 23256 33096 23262 33108
rect 23256 33068 25176 33096
rect 23256 33056 23262 33068
rect 23658 33028 23664 33040
rect 17236 33000 22094 33028
rect 22204 33000 23664 33028
rect 5491 32997 5503 33000
rect 5445 32991 5503 32997
rect 6457 32963 6515 32969
rect 6457 32929 6469 32963
rect 6503 32960 6515 32963
rect 7006 32960 7012 32972
rect 6503 32932 7012 32960
rect 6503 32929 6515 32932
rect 6457 32923 6515 32929
rect 7006 32920 7012 32932
rect 7064 32920 7070 32972
rect 9125 32963 9183 32969
rect 9125 32960 9137 32963
rect 7300 32932 9137 32960
rect 4065 32895 4123 32901
rect 4065 32861 4077 32895
rect 4111 32892 4123 32895
rect 4154 32892 4160 32904
rect 4111 32864 4160 32892
rect 4111 32861 4123 32864
rect 4065 32855 4123 32861
rect 4154 32852 4160 32864
rect 4212 32852 4218 32904
rect 4332 32895 4390 32901
rect 4332 32861 4344 32895
rect 4378 32892 4390 32895
rect 4890 32892 4896 32904
rect 4378 32864 4896 32892
rect 4378 32861 4390 32864
rect 4332 32855 4390 32861
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 6549 32895 6607 32901
rect 6549 32861 6561 32895
rect 6595 32861 6607 32895
rect 6549 32855 6607 32861
rect 6641 32895 6699 32901
rect 6641 32861 6653 32895
rect 6687 32861 6699 32895
rect 6641 32855 6699 32861
rect 6564 32756 6592 32855
rect 6656 32824 6684 32855
rect 6730 32852 6736 32904
rect 6788 32892 6794 32904
rect 7300 32892 7328 32932
rect 9125 32929 9137 32932
rect 9171 32929 9183 32963
rect 9125 32923 9183 32929
rect 9309 32963 9367 32969
rect 9309 32929 9321 32963
rect 9355 32960 9367 32963
rect 9766 32960 9772 32972
rect 9355 32932 9772 32960
rect 9355 32929 9367 32932
rect 9309 32923 9367 32929
rect 9766 32920 9772 32932
rect 9824 32920 9830 32972
rect 15102 32920 15108 32972
rect 15160 32960 15166 32972
rect 17957 32963 18015 32969
rect 17957 32960 17969 32963
rect 15160 32932 17969 32960
rect 15160 32920 15166 32932
rect 17957 32929 17969 32932
rect 18003 32929 18015 32963
rect 17957 32923 18015 32929
rect 18046 32920 18052 32972
rect 18104 32920 18110 32972
rect 20993 32963 21051 32969
rect 20993 32960 21005 32963
rect 18156 32932 21005 32960
rect 8018 32892 8024 32904
rect 6788 32864 7328 32892
rect 7392 32864 8024 32892
rect 6788 32852 6794 32864
rect 7006 32824 7012 32836
rect 6656 32796 7012 32824
rect 7006 32784 7012 32796
rect 7064 32784 7070 32836
rect 7392 32756 7420 32864
rect 8018 32852 8024 32864
rect 8076 32852 8082 32904
rect 8110 32852 8116 32904
rect 8168 32892 8174 32904
rect 8205 32895 8263 32901
rect 8205 32892 8217 32895
rect 8168 32864 8217 32892
rect 8168 32852 8174 32864
rect 8205 32861 8217 32864
rect 8251 32861 8263 32895
rect 8205 32855 8263 32861
rect 9398 32852 9404 32904
rect 9456 32852 9462 32904
rect 9493 32895 9551 32901
rect 9493 32861 9505 32895
rect 9539 32861 9551 32895
rect 9493 32855 9551 32861
rect 9585 32895 9643 32901
rect 9585 32861 9597 32895
rect 9631 32892 9643 32895
rect 10962 32892 10968 32904
rect 9631 32864 10968 32892
rect 9631 32861 9643 32864
rect 9585 32855 9643 32861
rect 7650 32784 7656 32836
rect 7708 32824 7714 32836
rect 9508 32824 9536 32855
rect 10962 32852 10968 32864
rect 11020 32852 11026 32904
rect 11698 32852 11704 32904
rect 11756 32892 11762 32904
rect 11756 32864 12204 32892
rect 11756 32852 11762 32864
rect 7708 32796 9536 32824
rect 7708 32784 7714 32796
rect 9950 32784 9956 32836
rect 10008 32824 10014 32836
rect 10597 32827 10655 32833
rect 10597 32824 10609 32827
rect 10008 32796 10609 32824
rect 10008 32784 10014 32796
rect 10597 32793 10609 32796
rect 10643 32824 10655 32827
rect 10686 32824 10692 32836
rect 10643 32796 10692 32824
rect 10643 32793 10655 32796
rect 10597 32787 10655 32793
rect 10686 32784 10692 32796
rect 10744 32784 10750 32836
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 12069 32827 12127 32833
rect 12069 32824 12081 32827
rect 12032 32796 12081 32824
rect 12032 32784 12038 32796
rect 12069 32793 12081 32796
rect 12115 32793 12127 32827
rect 12176 32824 12204 32864
rect 12250 32852 12256 32904
rect 12308 32892 12314 32904
rect 16390 32892 16396 32904
rect 12308 32864 16396 32892
rect 12308 32852 12314 32864
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 18156 32892 18184 32932
rect 20993 32929 21005 32932
rect 21039 32929 21051 32963
rect 20993 32923 21051 32929
rect 16540 32864 18184 32892
rect 16540 32852 16546 32864
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 18380 32864 19625 32892
rect 18380 32852 18386 32864
rect 19613 32861 19625 32864
rect 19659 32861 19671 32895
rect 19613 32855 19671 32861
rect 19797 32895 19855 32901
rect 19797 32861 19809 32895
rect 19843 32892 19855 32895
rect 19886 32892 19892 32904
rect 19843 32864 19892 32892
rect 19843 32861 19855 32864
rect 19797 32855 19855 32861
rect 19886 32852 19892 32864
rect 19944 32852 19950 32904
rect 19978 32852 19984 32904
rect 20036 32852 20042 32904
rect 21358 32852 21364 32904
rect 21416 32852 21422 32904
rect 22066 32901 22094 33000
rect 23658 32988 23664 33000
rect 23716 32988 23722 33040
rect 22646 32920 22652 32972
rect 22704 32920 22710 32972
rect 24118 32920 24124 32972
rect 24176 32960 24182 32972
rect 24581 32963 24639 32969
rect 24581 32960 24593 32963
rect 24176 32932 24593 32960
rect 24176 32920 24182 32932
rect 24581 32929 24593 32932
rect 24627 32929 24639 32963
rect 24581 32923 24639 32929
rect 24762 32920 24768 32972
rect 24820 32960 24826 32972
rect 25041 32963 25099 32969
rect 25041 32960 25053 32963
rect 24820 32932 25053 32960
rect 24820 32920 24826 32932
rect 25041 32929 25053 32932
rect 25087 32929 25099 32963
rect 25148 32960 25176 33068
rect 25222 33056 25228 33108
rect 25280 33096 25286 33108
rect 25777 33099 25835 33105
rect 25777 33096 25789 33099
rect 25280 33068 25789 33096
rect 25280 33056 25286 33068
rect 25777 33065 25789 33068
rect 25823 33065 25835 33099
rect 25777 33059 25835 33065
rect 27157 33099 27215 33105
rect 27157 33065 27169 33099
rect 27203 33065 27215 33099
rect 27157 33059 27215 33065
rect 27341 33099 27399 33105
rect 27341 33065 27353 33099
rect 27387 33096 27399 33099
rect 27614 33096 27620 33108
rect 27387 33068 27620 33096
rect 27387 33065 27399 33068
rect 27341 33059 27399 33065
rect 25961 33031 26019 33037
rect 25961 32997 25973 33031
rect 26007 33028 26019 33031
rect 26970 33028 26976 33040
rect 26007 33000 26976 33028
rect 26007 32997 26019 33000
rect 25961 32991 26019 32997
rect 26970 32988 26976 33000
rect 27028 32988 27034 33040
rect 27172 33028 27200 33059
rect 27614 33056 27620 33068
rect 27672 33056 27678 33108
rect 28258 33056 28264 33108
rect 28316 33056 28322 33108
rect 28721 33099 28779 33105
rect 28721 33065 28733 33099
rect 28767 33096 28779 33099
rect 28902 33096 28908 33108
rect 28767 33068 28908 33096
rect 28767 33065 28779 33068
rect 28721 33059 28779 33065
rect 28902 33056 28908 33068
rect 28960 33056 28966 33108
rect 38933 33099 38991 33105
rect 38933 33096 38945 33099
rect 38304 33068 38945 33096
rect 30469 33031 30527 33037
rect 30469 33028 30481 33031
rect 27172 33000 30481 33028
rect 30469 32997 30481 33000
rect 30515 33028 30527 33031
rect 35526 33028 35532 33040
rect 30515 33000 35532 33028
rect 30515 32997 30527 33000
rect 30469 32991 30527 32997
rect 35526 32988 35532 33000
rect 35584 32988 35590 33040
rect 37366 32988 37372 33040
rect 37424 33028 37430 33040
rect 37424 33000 38153 33028
rect 37424 32988 37430 33000
rect 25148 32932 26188 32960
rect 25041 32923 25099 32929
rect 22030 32895 22094 32901
rect 22030 32861 22042 32895
rect 22076 32864 22094 32895
rect 22076 32861 22088 32864
rect 22030 32855 22088 32861
rect 22830 32852 22836 32904
rect 22888 32852 22894 32904
rect 23017 32895 23075 32901
rect 23017 32861 23029 32895
rect 23063 32861 23075 32895
rect 23017 32855 23075 32861
rect 15470 32824 15476 32836
rect 12176 32796 15476 32824
rect 12069 32787 12127 32793
rect 15470 32784 15476 32796
rect 15528 32784 15534 32836
rect 17862 32784 17868 32836
rect 17920 32784 17926 32836
rect 19334 32824 19340 32836
rect 17972 32796 19340 32824
rect 6564 32728 7420 32756
rect 7469 32759 7527 32765
rect 7469 32725 7481 32759
rect 7515 32756 7527 32759
rect 7742 32756 7748 32768
rect 7515 32728 7748 32756
rect 7515 32725 7527 32728
rect 7469 32719 7527 32725
rect 7742 32716 7748 32728
rect 7800 32716 7806 32768
rect 8662 32716 8668 32768
rect 8720 32756 8726 32768
rect 10042 32756 10048 32768
rect 8720 32728 10048 32756
rect 8720 32716 8726 32728
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 10318 32716 10324 32768
rect 10376 32756 10382 32768
rect 10797 32759 10855 32765
rect 10797 32756 10809 32759
rect 10376 32728 10809 32756
rect 10376 32716 10382 32728
rect 10797 32725 10809 32728
rect 10843 32725 10855 32759
rect 10797 32719 10855 32725
rect 11330 32716 11336 32768
rect 11388 32756 11394 32768
rect 12269 32759 12327 32765
rect 12269 32756 12281 32759
rect 11388 32728 12281 32756
rect 11388 32716 11394 32728
rect 12269 32725 12281 32728
rect 12315 32725 12327 32759
rect 12269 32719 12327 32725
rect 12437 32759 12495 32765
rect 12437 32725 12449 32759
rect 12483 32756 12495 32759
rect 12802 32756 12808 32768
rect 12483 32728 12808 32756
rect 12483 32725 12495 32728
rect 12437 32719 12495 32725
rect 12802 32716 12808 32728
rect 12860 32716 12866 32768
rect 14182 32716 14188 32768
rect 14240 32756 14246 32768
rect 17972 32756 18000 32796
rect 19334 32784 19340 32796
rect 19392 32784 19398 32836
rect 19705 32827 19763 32833
rect 19705 32793 19717 32827
rect 19751 32793 19763 32827
rect 19904 32824 19932 32852
rect 20438 32824 20444 32836
rect 19904 32796 20444 32824
rect 19705 32787 19763 32793
rect 14240 32728 18000 32756
rect 14240 32716 14246 32728
rect 18414 32716 18420 32768
rect 18472 32756 18478 32768
rect 19429 32759 19487 32765
rect 19429 32756 19441 32759
rect 18472 32728 19441 32756
rect 18472 32716 18478 32728
rect 19429 32725 19441 32728
rect 19475 32725 19487 32759
rect 19720 32756 19748 32787
rect 20438 32784 20444 32796
rect 20496 32784 20502 32836
rect 21269 32827 21327 32833
rect 21269 32793 21281 32827
rect 21315 32824 21327 32827
rect 22462 32824 22468 32836
rect 21315 32796 22468 32824
rect 21315 32793 21327 32796
rect 21269 32787 21327 32793
rect 22462 32784 22468 32796
rect 22520 32824 22526 32836
rect 23032 32824 23060 32855
rect 23658 32852 23664 32904
rect 23716 32852 23722 32904
rect 24302 32852 24308 32904
rect 24360 32892 24366 32904
rect 25133 32895 25191 32901
rect 25133 32892 25145 32895
rect 24360 32864 25145 32892
rect 24360 32852 24366 32864
rect 25133 32861 25145 32864
rect 25179 32861 25191 32895
rect 26160 32892 26188 32932
rect 26694 32920 26700 32972
rect 26752 32960 26758 32972
rect 27065 32963 27123 32969
rect 27065 32960 27077 32963
rect 26752 32932 27077 32960
rect 26752 32920 26758 32932
rect 27065 32929 27077 32932
rect 27111 32929 27123 32963
rect 29730 32960 29736 32972
rect 27065 32923 27123 32929
rect 28460 32932 29736 32960
rect 26160 32864 26832 32892
rect 25133 32855 25191 32861
rect 22520 32796 23060 32824
rect 22520 32784 22526 32796
rect 26142 32784 26148 32836
rect 26200 32824 26206 32836
rect 26237 32827 26295 32833
rect 26237 32824 26249 32827
rect 26200 32796 26249 32824
rect 26200 32784 26206 32796
rect 26237 32793 26249 32796
rect 26283 32793 26295 32827
rect 26804 32824 26832 32864
rect 26878 32852 26884 32904
rect 26936 32892 26942 32904
rect 28460 32901 28488 32932
rect 29730 32920 29736 32932
rect 29788 32920 29794 32972
rect 30190 32920 30196 32972
rect 30248 32960 30254 32972
rect 33502 32960 33508 32972
rect 30248 32932 33508 32960
rect 30248 32920 30254 32932
rect 26973 32895 27031 32901
rect 26973 32892 26985 32895
rect 26936 32864 26985 32892
rect 26936 32852 26942 32864
rect 26973 32861 26985 32864
rect 27019 32861 27031 32895
rect 28445 32895 28503 32901
rect 28445 32892 28457 32895
rect 26973 32855 27031 32861
rect 27080 32864 28457 32892
rect 27080 32824 27108 32864
rect 28445 32861 28457 32864
rect 28491 32861 28503 32895
rect 28445 32855 28503 32861
rect 28537 32895 28595 32901
rect 28537 32861 28549 32895
rect 28583 32892 28595 32895
rect 29822 32892 29828 32904
rect 28583 32864 29828 32892
rect 28583 32861 28595 32864
rect 28537 32855 28595 32861
rect 29822 32852 29828 32864
rect 29880 32852 29886 32904
rect 30282 32852 30288 32904
rect 30340 32852 30346 32904
rect 30466 32852 30472 32904
rect 30524 32892 30530 32904
rect 30834 32892 30840 32904
rect 30524 32864 30840 32892
rect 30524 32852 30530 32864
rect 30834 32852 30840 32864
rect 30892 32892 30898 32904
rect 31220 32901 31248 32932
rect 33502 32920 33508 32932
rect 33560 32920 33566 32972
rect 33962 32920 33968 32972
rect 34020 32960 34026 32972
rect 34977 32963 35035 32969
rect 34977 32960 34989 32963
rect 34020 32932 34989 32960
rect 34020 32920 34026 32932
rect 34977 32929 34989 32932
rect 35023 32960 35035 32963
rect 35250 32960 35256 32972
rect 35023 32932 35256 32960
rect 35023 32929 35035 32932
rect 34977 32923 35035 32929
rect 35250 32920 35256 32932
rect 35308 32920 35314 32972
rect 35342 32920 35348 32972
rect 35400 32960 35406 32972
rect 35400 32932 36216 32960
rect 35400 32920 35406 32932
rect 36188 32904 36216 32932
rect 38010 32920 38016 32972
rect 38068 32920 38074 32972
rect 30929 32895 30987 32901
rect 30929 32892 30941 32895
rect 30892 32864 30941 32892
rect 30892 32852 30898 32864
rect 30929 32861 30941 32864
rect 30975 32861 30987 32895
rect 30929 32855 30987 32861
rect 31205 32895 31263 32901
rect 31205 32861 31217 32895
rect 31251 32861 31263 32895
rect 31205 32855 31263 32861
rect 33318 32852 33324 32904
rect 33376 32852 33382 32904
rect 33410 32852 33416 32904
rect 33468 32892 33474 32904
rect 34057 32895 34115 32901
rect 34057 32892 34069 32895
rect 33468 32864 34069 32892
rect 33468 32852 33474 32864
rect 34057 32861 34069 32864
rect 34103 32892 34115 32895
rect 34422 32892 34428 32904
rect 34103 32864 34428 32892
rect 34103 32861 34115 32864
rect 34057 32855 34115 32861
rect 34422 32852 34428 32864
rect 34480 32852 34486 32904
rect 35529 32895 35587 32901
rect 35529 32861 35541 32895
rect 35575 32892 35587 32895
rect 35710 32892 35716 32904
rect 35575 32864 35716 32892
rect 35575 32861 35587 32864
rect 35529 32855 35587 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 35894 32852 35900 32904
rect 35952 32892 35958 32904
rect 36081 32895 36139 32901
rect 36081 32892 36093 32895
rect 35952 32864 36093 32892
rect 35952 32852 35958 32864
rect 36081 32861 36093 32864
rect 36127 32861 36139 32895
rect 36081 32855 36139 32861
rect 36170 32852 36176 32904
rect 36228 32852 36234 32904
rect 36546 32895 36604 32901
rect 36546 32861 36558 32895
rect 36592 32892 36604 32895
rect 37366 32892 37372 32904
rect 36592 32864 37372 32892
rect 36592 32861 36604 32864
rect 36546 32855 36604 32861
rect 37366 32852 37372 32864
rect 37424 32852 37430 32904
rect 37458 32852 37464 32904
rect 37516 32892 37522 32904
rect 37645 32895 37703 32901
rect 37645 32892 37657 32895
rect 37516 32864 37657 32892
rect 37516 32852 37522 32864
rect 37645 32861 37657 32864
rect 37691 32861 37703 32895
rect 37645 32855 37703 32861
rect 37793 32895 37851 32901
rect 37793 32861 37805 32895
rect 37839 32892 37851 32895
rect 38028 32892 38056 32920
rect 38125 32901 38153 33000
rect 37839 32864 38056 32892
rect 38110 32895 38168 32901
rect 37839 32861 37851 32864
rect 37793 32855 37851 32861
rect 38110 32861 38122 32895
rect 38156 32861 38168 32895
rect 38110 32855 38168 32861
rect 26804 32796 27108 32824
rect 28261 32827 28319 32833
rect 26237 32787 26295 32793
rect 28261 32793 28273 32827
rect 28307 32824 28319 32827
rect 28718 32824 28724 32836
rect 28307 32796 28724 32824
rect 28307 32793 28319 32796
rect 28261 32787 28319 32793
rect 28718 32784 28724 32796
rect 28776 32784 28782 32836
rect 28810 32784 28816 32836
rect 28868 32824 28874 32836
rect 32398 32824 32404 32836
rect 28868 32796 32404 32824
rect 28868 32784 28874 32796
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 34974 32784 34980 32836
rect 35032 32824 35038 32836
rect 36357 32827 36415 32833
rect 36357 32824 36369 32827
rect 35032 32796 36369 32824
rect 35032 32784 35038 32796
rect 36096 32768 36124 32796
rect 36357 32793 36369 32796
rect 36403 32793 36415 32827
rect 36357 32787 36415 32793
rect 19978 32756 19984 32768
rect 19720 32728 19984 32756
rect 19429 32719 19487 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 21174 32716 21180 32768
rect 21232 32716 21238 32768
rect 21545 32759 21603 32765
rect 21545 32725 21557 32759
rect 21591 32756 21603 32759
rect 23382 32756 23388 32768
rect 21591 32728 23388 32756
rect 21591 32725 21603 32728
rect 21545 32719 21603 32725
rect 23382 32716 23388 32728
rect 23440 32716 23446 32768
rect 24762 32716 24768 32768
rect 24820 32716 24826 32768
rect 26970 32716 26976 32768
rect 27028 32756 27034 32768
rect 29638 32756 29644 32768
rect 27028 32728 29644 32756
rect 27028 32716 27034 32728
rect 29638 32716 29644 32728
rect 29696 32716 29702 32768
rect 34057 32759 34115 32765
rect 34057 32725 34069 32759
rect 34103 32756 34115 32759
rect 34330 32756 34336 32768
rect 34103 32728 34336 32756
rect 34103 32725 34115 32728
rect 34057 32719 34115 32725
rect 34330 32716 34336 32728
rect 34388 32716 34394 32768
rect 36078 32716 36084 32768
rect 36136 32716 36142 32768
rect 36372 32756 36400 32787
rect 36446 32784 36452 32836
rect 36504 32784 36510 32836
rect 37921 32827 37979 32833
rect 37921 32824 37933 32827
rect 36648 32796 37933 32824
rect 36648 32756 36676 32796
rect 37921 32793 37933 32796
rect 37967 32793 37979 32827
rect 37921 32787 37979 32793
rect 38010 32784 38016 32836
rect 38068 32784 38074 32836
rect 38304 32824 38332 33068
rect 38933 33065 38945 33068
rect 38979 33065 38991 33099
rect 38933 33059 38991 33065
rect 38378 32852 38384 32904
rect 38436 32892 38442 32904
rect 38436 32864 39160 32892
rect 38436 32852 38442 32864
rect 38212 32796 38332 32824
rect 38749 32827 38807 32833
rect 36372 32728 36676 32756
rect 36725 32759 36783 32765
rect 36725 32725 36737 32759
rect 36771 32756 36783 32759
rect 37826 32756 37832 32768
rect 36771 32728 37832 32756
rect 36771 32725 36783 32728
rect 36725 32719 36783 32725
rect 37826 32716 37832 32728
rect 37884 32756 37890 32768
rect 38212 32756 38240 32796
rect 38749 32793 38761 32827
rect 38795 32824 38807 32827
rect 38838 32824 38844 32836
rect 38795 32796 38844 32824
rect 38795 32793 38807 32796
rect 38749 32787 38807 32793
rect 38838 32784 38844 32796
rect 38896 32784 38902 32836
rect 37884 32728 38240 32756
rect 38289 32759 38347 32765
rect 37884 32716 37890 32728
rect 38289 32725 38301 32759
rect 38335 32756 38347 32759
rect 38930 32756 38936 32768
rect 38335 32728 38936 32756
rect 38335 32725 38347 32728
rect 38289 32719 38347 32725
rect 38930 32716 38936 32728
rect 38988 32716 38994 32768
rect 39132 32765 39160 32864
rect 41414 32852 41420 32904
rect 41472 32892 41478 32904
rect 41874 32892 41880 32904
rect 41472 32864 41880 32892
rect 41472 32852 41478 32864
rect 41874 32852 41880 32864
rect 41932 32852 41938 32904
rect 42886 32852 42892 32904
rect 42944 32852 42950 32904
rect 39574 32784 39580 32836
rect 39632 32824 39638 32836
rect 41150 32827 41208 32833
rect 41150 32824 41162 32827
rect 39632 32796 41162 32824
rect 39632 32784 39638 32796
rect 41150 32793 41162 32796
rect 41196 32793 41208 32827
rect 41150 32787 41208 32793
rect 43162 32784 43168 32836
rect 43220 32784 43226 32836
rect 39117 32759 39175 32765
rect 39117 32725 39129 32759
rect 39163 32756 39175 32759
rect 39482 32756 39488 32768
rect 39163 32728 39488 32756
rect 39163 32725 39175 32728
rect 39117 32719 39175 32725
rect 39482 32716 39488 32728
rect 39540 32716 39546 32768
rect 40034 32716 40040 32768
rect 40092 32716 40098 32768
rect 1104 32666 43884 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 43884 32666
rect 1104 32592 43884 32614
rect 6638 32512 6644 32564
rect 6696 32552 6702 32564
rect 7101 32555 7159 32561
rect 7101 32552 7113 32555
rect 6696 32524 7113 32552
rect 6696 32512 6702 32524
rect 7101 32521 7113 32524
rect 7147 32521 7159 32555
rect 7101 32515 7159 32521
rect 7742 32512 7748 32564
rect 7800 32512 7806 32564
rect 9217 32555 9275 32561
rect 9217 32521 9229 32555
rect 9263 32552 9275 32555
rect 9398 32552 9404 32564
rect 9263 32524 9404 32552
rect 9263 32521 9275 32524
rect 9217 32515 9275 32521
rect 9398 32512 9404 32524
rect 9456 32512 9462 32564
rect 11330 32512 11336 32564
rect 11388 32552 11394 32564
rect 11885 32555 11943 32561
rect 11885 32552 11897 32555
rect 11388 32524 11897 32552
rect 11388 32512 11394 32524
rect 11885 32521 11897 32524
rect 11931 32521 11943 32555
rect 11885 32515 11943 32521
rect 12710 32512 12716 32564
rect 12768 32552 12774 32564
rect 13354 32552 13360 32564
rect 12768 32524 13360 32552
rect 12768 32512 12774 32524
rect 13354 32512 13360 32524
rect 13412 32512 13418 32564
rect 13630 32512 13636 32564
rect 13688 32552 13694 32564
rect 14369 32555 14427 32561
rect 13688 32524 14228 32552
rect 13688 32512 13694 32524
rect 8665 32487 8723 32493
rect 8665 32484 8677 32487
rect 7668 32456 8677 32484
rect 7668 32428 7696 32456
rect 8665 32453 8677 32456
rect 8711 32453 8723 32487
rect 8665 32447 8723 32453
rect 9306 32444 9312 32496
rect 9364 32484 9370 32496
rect 9582 32484 9588 32496
rect 9364 32456 9588 32484
rect 9364 32444 9370 32456
rect 9582 32444 9588 32456
rect 9640 32444 9646 32496
rect 10778 32444 10784 32496
rect 10836 32484 10842 32496
rect 11701 32487 11759 32493
rect 11701 32484 11713 32487
rect 10836 32456 11713 32484
rect 10836 32444 10842 32456
rect 11701 32453 11713 32456
rect 11747 32484 11759 32487
rect 12434 32484 12440 32496
rect 11747 32456 12440 32484
rect 11747 32453 11759 32456
rect 11701 32447 11759 32453
rect 12434 32444 12440 32456
rect 12492 32444 12498 32496
rect 12989 32487 13047 32493
rect 12989 32453 13001 32487
rect 13035 32484 13047 32487
rect 13035 32456 13860 32484
rect 13035 32453 13047 32456
rect 12989 32447 13047 32453
rect 4240 32419 4298 32425
rect 4240 32385 4252 32419
rect 4286 32416 4298 32419
rect 4706 32416 4712 32428
rect 4286 32388 4712 32416
rect 4286 32385 4298 32388
rect 4240 32379 4298 32385
rect 4706 32376 4712 32388
rect 4764 32376 4770 32428
rect 7282 32376 7288 32428
rect 7340 32376 7346 32428
rect 7377 32419 7435 32425
rect 7377 32385 7389 32419
rect 7423 32416 7435 32419
rect 7650 32416 7656 32428
rect 7423 32388 7656 32416
rect 7423 32385 7435 32388
rect 7377 32379 7435 32385
rect 7650 32376 7656 32388
rect 7708 32376 7714 32428
rect 8570 32376 8576 32428
rect 8628 32376 8634 32428
rect 8757 32419 8815 32425
rect 8757 32385 8769 32419
rect 8803 32385 8815 32419
rect 8757 32379 8815 32385
rect 9401 32419 9459 32425
rect 9401 32385 9413 32419
rect 9447 32416 9459 32419
rect 9490 32416 9496 32428
rect 9447 32388 9496 32416
rect 9447 32385 9459 32388
rect 9401 32379 9459 32385
rect 3973 32351 4031 32357
rect 3973 32317 3985 32351
rect 4019 32317 4031 32351
rect 3973 32311 4031 32317
rect 3988 32212 4016 32311
rect 7006 32308 7012 32360
rect 7064 32348 7070 32360
rect 7558 32348 7564 32360
rect 7064 32320 7564 32348
rect 7064 32308 7070 32320
rect 7558 32308 7564 32320
rect 7616 32348 7622 32360
rect 8772 32348 8800 32379
rect 9490 32376 9496 32388
rect 9548 32376 9554 32428
rect 9674 32376 9680 32428
rect 9732 32416 9738 32428
rect 12161 32419 12219 32425
rect 9732 32388 11744 32416
rect 9732 32376 9738 32388
rect 11716 32360 11744 32388
rect 12161 32385 12173 32419
rect 12207 32385 12219 32419
rect 12161 32379 12219 32385
rect 10778 32348 10784 32360
rect 7616 32320 10784 32348
rect 7616 32308 7622 32320
rect 10778 32308 10784 32320
rect 10836 32308 10842 32360
rect 11698 32308 11704 32360
rect 11756 32308 11762 32360
rect 12066 32308 12072 32360
rect 12124 32348 12130 32360
rect 12176 32348 12204 32379
rect 12802 32376 12808 32428
rect 12860 32376 12866 32428
rect 13078 32376 13084 32428
rect 13136 32376 13142 32428
rect 13173 32419 13231 32425
rect 13173 32385 13185 32419
rect 13219 32416 13231 32419
rect 13630 32416 13636 32428
rect 13219 32388 13636 32416
rect 13219 32385 13231 32388
rect 13173 32379 13231 32385
rect 13630 32376 13636 32388
rect 13688 32376 13694 32428
rect 13832 32425 13860 32456
rect 13817 32419 13875 32425
rect 13817 32385 13829 32419
rect 13863 32416 13875 32419
rect 13906 32416 13912 32428
rect 13863 32388 13912 32416
rect 13863 32385 13875 32388
rect 13817 32379 13875 32385
rect 13906 32376 13912 32388
rect 13964 32376 13970 32428
rect 14200 32425 14228 32524
rect 14369 32521 14381 32555
rect 14415 32521 14427 32555
rect 14369 32515 14427 32521
rect 14384 32484 14412 32515
rect 16390 32512 16396 32564
rect 16448 32552 16454 32564
rect 16448 32524 19380 32552
rect 16448 32512 16454 32524
rect 15074 32487 15132 32493
rect 15074 32484 15086 32487
rect 14384 32456 15086 32484
rect 15074 32453 15086 32456
rect 15120 32453 15132 32487
rect 15074 32447 15132 32453
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 14093 32419 14151 32425
rect 14093 32385 14105 32419
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 14185 32419 14243 32425
rect 14185 32385 14197 32419
rect 14231 32416 14243 32419
rect 14734 32416 14740 32428
rect 14231 32388 14740 32416
rect 14231 32385 14243 32388
rect 14185 32379 14243 32385
rect 14016 32348 14044 32379
rect 12124 32320 14044 32348
rect 12124 32308 12130 32320
rect 5350 32240 5356 32292
rect 5408 32280 5414 32292
rect 12250 32280 12256 32292
rect 5408 32252 12256 32280
rect 5408 32240 5414 32252
rect 12250 32240 12256 32252
rect 12308 32240 12314 32292
rect 14108 32280 14136 32379
rect 14734 32376 14740 32388
rect 14792 32416 14798 32428
rect 14792 32388 15976 32416
rect 14792 32376 14798 32388
rect 14274 32308 14280 32360
rect 14332 32348 14338 32360
rect 14829 32351 14887 32357
rect 14829 32348 14841 32351
rect 14332 32320 14841 32348
rect 14332 32308 14338 32320
rect 14829 32317 14841 32320
rect 14875 32317 14887 32351
rect 15948 32348 15976 32388
rect 18138 32376 18144 32428
rect 18196 32416 18202 32428
rect 19242 32416 19248 32428
rect 18196 32388 19248 32416
rect 18196 32376 18202 32388
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 18322 32348 18328 32360
rect 15948 32320 18328 32348
rect 14829 32311 14887 32317
rect 18322 32308 18328 32320
rect 18380 32308 18386 32360
rect 18414 32308 18420 32360
rect 18472 32308 18478 32360
rect 19352 32348 19380 32524
rect 20254 32512 20260 32564
rect 20312 32512 20318 32564
rect 20622 32512 20628 32564
rect 20680 32512 20686 32564
rect 21174 32512 21180 32564
rect 21232 32552 21238 32564
rect 22830 32552 22836 32564
rect 21232 32524 22836 32552
rect 21232 32512 21238 32524
rect 22830 32512 22836 32524
rect 22888 32552 22894 32564
rect 25314 32552 25320 32564
rect 22888 32524 25320 32552
rect 22888 32512 22894 32524
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 25958 32512 25964 32564
rect 26016 32552 26022 32564
rect 26145 32555 26203 32561
rect 26145 32552 26157 32555
rect 26016 32524 26157 32552
rect 26016 32512 26022 32524
rect 26145 32521 26157 32524
rect 26191 32521 26203 32555
rect 26145 32515 26203 32521
rect 27249 32555 27307 32561
rect 27249 32521 27261 32555
rect 27295 32552 27307 32555
rect 27338 32552 27344 32564
rect 27295 32524 27344 32552
rect 27295 32521 27307 32524
rect 27249 32515 27307 32521
rect 27338 32512 27344 32524
rect 27396 32512 27402 32564
rect 27522 32512 27528 32564
rect 27580 32552 27586 32564
rect 27706 32552 27712 32564
rect 27580 32524 27712 32552
rect 27580 32512 27586 32524
rect 27706 32512 27712 32524
rect 27764 32552 27770 32564
rect 29457 32555 29515 32561
rect 27764 32524 29408 32552
rect 27764 32512 27770 32524
rect 19426 32444 19432 32496
rect 19484 32484 19490 32496
rect 24762 32484 24768 32496
rect 19484 32456 24768 32484
rect 19484 32444 19490 32456
rect 24762 32444 24768 32456
rect 24820 32444 24826 32496
rect 25774 32484 25780 32496
rect 25516 32456 25780 32484
rect 20438 32376 20444 32428
rect 20496 32376 20502 32428
rect 20717 32419 20775 32425
rect 20717 32385 20729 32419
rect 20763 32416 20775 32419
rect 22186 32416 22192 32428
rect 20763 32388 22192 32416
rect 20763 32385 20775 32388
rect 20717 32379 20775 32385
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32416 22891 32419
rect 22922 32416 22928 32428
rect 22879 32388 22928 32416
rect 22879 32385 22891 32388
rect 22833 32379 22891 32385
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23198 32376 23204 32428
rect 23256 32376 23262 32428
rect 23382 32376 23388 32428
rect 23440 32376 23446 32428
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 22204 32348 22232 32376
rect 23014 32348 23020 32360
rect 19352 32320 22094 32348
rect 22204 32320 23020 32348
rect 22066 32280 22094 32320
rect 23014 32308 23020 32320
rect 23072 32308 23078 32360
rect 23584 32280 23612 32379
rect 23658 32376 23664 32428
rect 23716 32416 23722 32428
rect 23842 32416 23848 32428
rect 23716 32388 23848 32416
rect 23716 32376 23722 32388
rect 23842 32376 23848 32388
rect 23900 32376 23906 32428
rect 25222 32376 25228 32428
rect 25280 32416 25286 32428
rect 25516 32425 25544 32456
rect 25774 32444 25780 32456
rect 25832 32444 25838 32496
rect 28258 32484 28264 32496
rect 26344 32456 28264 32484
rect 25501 32419 25559 32425
rect 25501 32416 25513 32419
rect 25280 32388 25513 32416
rect 25280 32376 25286 32388
rect 25501 32385 25513 32388
rect 25547 32385 25559 32419
rect 25501 32379 25559 32385
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32416 25743 32419
rect 26050 32416 26056 32428
rect 25731 32388 26056 32416
rect 25731 32385 25743 32388
rect 25685 32379 25743 32385
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26344 32425 26372 32456
rect 28258 32444 28264 32456
rect 28316 32444 28322 32496
rect 28552 32493 28580 32524
rect 28537 32487 28595 32493
rect 28537 32453 28549 32487
rect 28583 32453 28595 32487
rect 28537 32447 28595 32453
rect 28721 32487 28779 32493
rect 28721 32453 28733 32487
rect 28767 32484 28779 32487
rect 28810 32484 28816 32496
rect 28767 32456 28816 32484
rect 28767 32453 28779 32456
rect 28721 32447 28779 32453
rect 26329 32419 26387 32425
rect 26329 32385 26341 32419
rect 26375 32385 26387 32419
rect 26329 32379 26387 32385
rect 26510 32376 26516 32428
rect 26568 32376 26574 32428
rect 26605 32419 26663 32425
rect 26605 32385 26617 32419
rect 26651 32385 26663 32419
rect 26605 32379 26663 32385
rect 27433 32419 27491 32425
rect 27433 32385 27445 32419
rect 27479 32416 27491 32419
rect 27522 32416 27528 32428
rect 27479 32388 27528 32416
rect 27479 32385 27491 32388
rect 27433 32379 27491 32385
rect 26620 32348 26648 32379
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 27709 32419 27767 32425
rect 27709 32385 27721 32419
rect 27755 32385 27767 32419
rect 27709 32379 27767 32385
rect 27893 32419 27951 32425
rect 27893 32385 27905 32419
rect 27939 32416 27951 32419
rect 28353 32419 28411 32425
rect 28353 32416 28365 32419
rect 27939 32388 28365 32416
rect 27939 32385 27951 32388
rect 27893 32379 27951 32385
rect 28353 32385 28365 32388
rect 28399 32416 28411 32419
rect 28442 32416 28448 32428
rect 28399 32388 28448 32416
rect 28399 32385 28411 32388
rect 28353 32379 28411 32385
rect 27617 32351 27675 32357
rect 27617 32348 27629 32351
rect 14108 32252 14688 32280
rect 4154 32212 4160 32224
rect 3988 32184 4160 32212
rect 4154 32172 4160 32184
rect 4212 32212 4218 32224
rect 4614 32212 4620 32224
rect 4212 32184 4620 32212
rect 4212 32172 4218 32184
rect 4614 32172 4620 32184
rect 4672 32172 4678 32224
rect 8018 32172 8024 32224
rect 8076 32212 8082 32224
rect 10318 32212 10324 32224
rect 8076 32184 10324 32212
rect 8076 32172 8082 32184
rect 10318 32172 10324 32184
rect 10376 32212 10382 32224
rect 11606 32212 11612 32224
rect 10376 32184 11612 32212
rect 10376 32172 10382 32184
rect 11606 32172 11612 32184
rect 11664 32212 11670 32224
rect 11885 32215 11943 32221
rect 11885 32212 11897 32215
rect 11664 32184 11897 32212
rect 11664 32172 11670 32184
rect 11885 32181 11897 32184
rect 11931 32181 11943 32215
rect 11885 32175 11943 32181
rect 13357 32215 13415 32221
rect 13357 32181 13369 32215
rect 13403 32212 13415 32215
rect 14550 32212 14556 32224
rect 13403 32184 14556 32212
rect 13403 32181 13415 32184
rect 13357 32175 13415 32181
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 14660 32212 14688 32252
rect 19076 32252 20116 32280
rect 22066 32252 23612 32280
rect 23676 32320 27629 32348
rect 16206 32212 16212 32224
rect 14660 32184 16212 32212
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 16298 32172 16304 32224
rect 16356 32212 16362 32224
rect 19076 32212 19104 32252
rect 16356 32184 19104 32212
rect 19705 32215 19763 32221
rect 16356 32172 16362 32184
rect 19705 32181 19717 32215
rect 19751 32212 19763 32215
rect 19978 32212 19984 32224
rect 19751 32184 19984 32212
rect 19751 32181 19763 32184
rect 19705 32175 19763 32181
rect 19978 32172 19984 32184
rect 20036 32172 20042 32224
rect 20088 32212 20116 32252
rect 23106 32212 23112 32224
rect 20088 32184 23112 32212
rect 23106 32172 23112 32184
rect 23164 32172 23170 32224
rect 23474 32172 23480 32224
rect 23532 32212 23538 32224
rect 23676 32212 23704 32320
rect 27617 32317 27629 32320
rect 27663 32317 27675 32351
rect 27617 32311 27675 32317
rect 27724 32292 27752 32379
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 28258 32308 28264 32360
rect 28316 32348 28322 32360
rect 28552 32348 28580 32447
rect 28810 32444 28816 32456
rect 28868 32444 28874 32496
rect 29086 32376 29092 32428
rect 29144 32416 29150 32428
rect 29273 32419 29331 32425
rect 29273 32416 29285 32419
rect 29144 32388 29285 32416
rect 29144 32376 29150 32388
rect 29273 32385 29285 32388
rect 29319 32385 29331 32419
rect 29380 32416 29408 32524
rect 29457 32521 29469 32555
rect 29503 32552 29515 32555
rect 29822 32552 29828 32564
rect 29503 32524 29828 32552
rect 29503 32521 29515 32524
rect 29457 32515 29515 32521
rect 29822 32512 29828 32524
rect 29880 32512 29886 32564
rect 31726 32524 33364 32552
rect 31570 32484 31576 32496
rect 31128 32456 31576 32484
rect 31128 32425 31156 32456
rect 31570 32444 31576 32456
rect 31628 32444 31634 32496
rect 29457 32419 29515 32425
rect 29457 32416 29469 32419
rect 29380 32388 29469 32416
rect 29273 32379 29331 32385
rect 29457 32385 29469 32388
rect 29503 32416 29515 32419
rect 31113 32419 31171 32425
rect 31113 32416 31125 32419
rect 29503 32388 31125 32416
rect 29503 32385 29515 32388
rect 29457 32379 29515 32385
rect 31113 32385 31125 32388
rect 31159 32385 31171 32419
rect 31113 32379 31171 32385
rect 31478 32376 31484 32428
rect 31536 32376 31542 32428
rect 28316 32320 28580 32348
rect 28316 32308 28322 32320
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 30929 32351 30987 32357
rect 30929 32348 30941 32351
rect 30432 32320 30941 32348
rect 30432 32308 30438 32320
rect 30929 32317 30941 32320
rect 30975 32348 30987 32351
rect 31726 32348 31754 32524
rect 32490 32444 32496 32496
rect 32548 32444 32554 32496
rect 33336 32484 33364 32524
rect 34330 32512 34336 32564
rect 34388 32552 34394 32564
rect 34388 32524 36308 32552
rect 34388 32512 34394 32524
rect 34514 32484 34520 32496
rect 33336 32456 34520 32484
rect 34514 32444 34520 32456
rect 34572 32444 34578 32496
rect 36280 32484 36308 32524
rect 36354 32512 36360 32564
rect 36412 32552 36418 32564
rect 36412 32524 36584 32552
rect 36412 32512 36418 32524
rect 36556 32493 36584 32524
rect 36906 32512 36912 32564
rect 36964 32512 36970 32564
rect 39574 32512 39580 32564
rect 39632 32512 39638 32564
rect 36541 32487 36599 32493
rect 36280 32456 36492 32484
rect 33502 32376 33508 32428
rect 33560 32376 33566 32428
rect 34422 32376 34428 32428
rect 34480 32416 34486 32428
rect 34609 32419 34667 32425
rect 34609 32416 34621 32419
rect 34480 32388 34621 32416
rect 34480 32376 34486 32388
rect 34609 32385 34621 32388
rect 34655 32385 34667 32419
rect 34609 32379 34667 32385
rect 34974 32376 34980 32428
rect 35032 32376 35038 32428
rect 35250 32376 35256 32428
rect 35308 32376 35314 32428
rect 35986 32376 35992 32428
rect 36044 32416 36050 32428
rect 36265 32419 36323 32425
rect 36265 32416 36277 32419
rect 36044 32388 36277 32416
rect 36044 32376 36050 32388
rect 36265 32385 36277 32388
rect 36311 32385 36323 32419
rect 36265 32379 36323 32385
rect 36358 32419 36416 32425
rect 36358 32385 36370 32419
rect 36404 32385 36416 32419
rect 36464 32416 36492 32456
rect 36541 32453 36553 32487
rect 36587 32453 36599 32487
rect 36541 32447 36599 32453
rect 36633 32487 36691 32493
rect 36633 32453 36645 32487
rect 36679 32484 36691 32487
rect 37918 32484 37924 32496
rect 36679 32456 37924 32484
rect 36679 32453 36691 32456
rect 36633 32447 36691 32453
rect 37918 32444 37924 32456
rect 37976 32444 37982 32496
rect 38120 32456 38884 32484
rect 38120 32425 38148 32456
rect 38856 32428 38884 32456
rect 38930 32444 38936 32496
rect 38988 32484 38994 32496
rect 39025 32487 39083 32493
rect 39025 32484 39037 32487
rect 38988 32456 39037 32484
rect 38988 32444 38994 32456
rect 39025 32453 39037 32456
rect 39071 32453 39083 32487
rect 39942 32484 39948 32496
rect 39025 32447 39083 32453
rect 39132 32456 39948 32484
rect 36730 32419 36788 32425
rect 36730 32416 36742 32419
rect 36464 32388 36742 32416
rect 36358 32379 36416 32385
rect 30975 32320 31754 32348
rect 30975 32317 30987 32320
rect 30929 32311 30987 32317
rect 25409 32283 25467 32289
rect 25409 32249 25421 32283
rect 25455 32280 25467 32283
rect 26786 32280 26792 32292
rect 25455 32252 26792 32280
rect 25455 32249 25467 32252
rect 25409 32243 25467 32249
rect 26786 32240 26792 32252
rect 26844 32240 26850 32292
rect 27525 32283 27583 32289
rect 27525 32249 27537 32283
rect 27571 32249 27583 32283
rect 27525 32243 27583 32249
rect 23532 32184 23704 32212
rect 23532 32172 23538 32184
rect 23750 32172 23756 32224
rect 23808 32212 23814 32224
rect 24213 32215 24271 32221
rect 24213 32212 24225 32215
rect 23808 32184 24225 32212
rect 23808 32172 23814 32184
rect 24213 32181 24225 32184
rect 24259 32181 24271 32215
rect 27540 32212 27568 32243
rect 27706 32240 27712 32292
rect 27764 32280 27770 32292
rect 31294 32280 31300 32292
rect 27764 32252 31300 32280
rect 27764 32240 27770 32252
rect 31294 32240 31300 32252
rect 31352 32240 31358 32292
rect 31846 32240 31852 32292
rect 31904 32280 31910 32292
rect 36372 32280 36400 32379
rect 36648 32360 36676 32388
rect 36730 32385 36742 32388
rect 36776 32385 36788 32419
rect 36730 32379 36788 32385
rect 38105 32419 38163 32425
rect 38105 32385 38117 32419
rect 38151 32385 38163 32419
rect 38105 32379 38163 32385
rect 38749 32419 38807 32425
rect 38749 32385 38761 32419
rect 38795 32385 38807 32419
rect 38749 32379 38807 32385
rect 36630 32308 36636 32360
rect 36688 32308 36694 32360
rect 37734 32308 37740 32360
rect 37792 32308 37798 32360
rect 37826 32308 37832 32360
rect 37884 32348 37890 32360
rect 38013 32351 38071 32357
rect 38013 32348 38025 32351
rect 37884 32320 38025 32348
rect 37884 32308 37890 32320
rect 38013 32317 38025 32320
rect 38059 32348 38071 32351
rect 38764 32348 38792 32379
rect 38838 32376 38844 32428
rect 38896 32416 38902 32428
rect 39132 32416 39160 32456
rect 39942 32444 39948 32456
rect 40000 32444 40006 32496
rect 38896 32388 39160 32416
rect 38896 32376 38902 32388
rect 39482 32376 39488 32428
rect 39540 32376 39546 32428
rect 39669 32419 39727 32425
rect 39669 32385 39681 32419
rect 39715 32385 39727 32419
rect 39669 32379 39727 32385
rect 39684 32348 39712 32379
rect 42978 32376 42984 32428
rect 43036 32376 43042 32428
rect 38059 32320 38792 32348
rect 39040 32320 39712 32348
rect 38059 32317 38071 32320
rect 38013 32311 38071 32317
rect 39040 32289 39068 32320
rect 40954 32308 40960 32360
rect 41012 32348 41018 32360
rect 42886 32348 42892 32360
rect 41012 32320 42892 32348
rect 41012 32308 41018 32320
rect 42886 32308 42892 32320
rect 42944 32348 42950 32360
rect 43073 32351 43131 32357
rect 43073 32348 43085 32351
rect 42944 32320 43085 32348
rect 42944 32308 42950 32320
rect 43073 32317 43085 32320
rect 43119 32317 43131 32351
rect 43073 32311 43131 32317
rect 43254 32308 43260 32360
rect 43312 32308 43318 32360
rect 39025 32283 39083 32289
rect 31904 32252 38976 32280
rect 31904 32240 31910 32252
rect 28074 32212 28080 32224
rect 27540 32184 28080 32212
rect 24213 32175 24271 32181
rect 28074 32172 28080 32184
rect 28132 32172 28138 32224
rect 34606 32172 34612 32224
rect 34664 32212 34670 32224
rect 34790 32212 34796 32224
rect 34664 32184 34796 32212
rect 34664 32172 34670 32184
rect 34790 32172 34796 32184
rect 34848 32172 34854 32224
rect 35710 32172 35716 32224
rect 35768 32212 35774 32224
rect 37734 32212 37740 32224
rect 35768 32184 37740 32212
rect 35768 32172 35774 32184
rect 37734 32172 37740 32184
rect 37792 32172 37798 32224
rect 38948 32212 38976 32252
rect 39025 32249 39037 32283
rect 39071 32249 39083 32283
rect 39025 32243 39083 32249
rect 40402 32212 40408 32224
rect 38948 32184 40408 32212
rect 40402 32172 40408 32184
rect 40460 32172 40466 32224
rect 42610 32172 42616 32224
rect 42668 32172 42674 32224
rect 1104 32122 43884 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 43884 32122
rect 1104 32048 43884 32070
rect 4617 32011 4675 32017
rect 4617 31977 4629 32011
rect 4663 32008 4675 32011
rect 4706 32008 4712 32020
rect 4663 31980 4712 32008
rect 4663 31977 4675 31980
rect 4617 31971 4675 31977
rect 4706 31968 4712 31980
rect 4764 31968 4770 32020
rect 9674 32008 9680 32020
rect 6196 31980 9680 32008
rect 5258 31832 5264 31884
rect 5316 31872 5322 31884
rect 6196 31872 6224 31980
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 10318 31968 10324 32020
rect 10376 31968 10382 32020
rect 11146 32008 11152 32020
rect 10428 31980 11152 32008
rect 8018 31900 8024 31952
rect 8076 31940 8082 31952
rect 8076 31912 9628 31940
rect 8076 31900 8082 31912
rect 7374 31872 7380 31884
rect 5316 31844 6224 31872
rect 6412 31844 7380 31872
rect 5316 31832 5322 31844
rect 6412 31813 6440 31844
rect 7374 31832 7380 31844
rect 7432 31832 7438 31884
rect 7466 31832 7472 31884
rect 7524 31872 7530 31884
rect 8202 31872 8208 31884
rect 7524 31844 8208 31872
rect 7524 31832 7530 31844
rect 8202 31832 8208 31844
rect 8260 31872 8266 31884
rect 9600 31872 9628 31912
rect 10428 31872 10456 31980
rect 11146 31968 11152 31980
rect 11204 31968 11210 32020
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 13136 31980 15700 32008
rect 13136 31968 13142 31980
rect 10870 31940 10876 31952
rect 10520 31912 10876 31940
rect 10520 31881 10548 31912
rect 10870 31900 10876 31912
rect 10928 31940 10934 31952
rect 11238 31940 11244 31952
rect 10928 31912 11244 31940
rect 10928 31900 10934 31912
rect 11238 31900 11244 31912
rect 11296 31900 11302 31952
rect 13354 31900 13360 31952
rect 13412 31900 13418 31952
rect 13449 31943 13507 31949
rect 13449 31909 13461 31943
rect 13495 31940 13507 31943
rect 13906 31940 13912 31952
rect 13495 31912 13912 31940
rect 13495 31909 13507 31912
rect 13449 31903 13507 31909
rect 13906 31900 13912 31912
rect 13964 31900 13970 31952
rect 15672 31949 15700 31980
rect 16206 31968 16212 32020
rect 16264 32008 16270 32020
rect 16264 31980 20392 32008
rect 16264 31968 16270 31980
rect 15657 31943 15715 31949
rect 15657 31909 15669 31943
rect 15703 31940 15715 31943
rect 16298 31940 16304 31952
rect 15703 31912 16304 31940
rect 15703 31909 15715 31912
rect 15657 31903 15715 31909
rect 16298 31900 16304 31912
rect 16356 31900 16362 31952
rect 17773 31943 17831 31949
rect 17773 31909 17785 31943
rect 17819 31940 17831 31943
rect 20364 31940 20392 31980
rect 22738 31968 22744 32020
rect 22796 32008 22802 32020
rect 23382 32008 23388 32020
rect 22796 31980 23388 32008
rect 22796 31968 22802 31980
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 26881 32011 26939 32017
rect 26881 31977 26893 32011
rect 26927 32008 26939 32011
rect 27706 32008 27712 32020
rect 26927 31980 27712 32008
rect 26927 31977 26939 31980
rect 26881 31971 26939 31977
rect 27706 31968 27712 31980
rect 27764 31968 27770 32020
rect 30834 32008 30840 32020
rect 28644 31980 30840 32008
rect 23201 31943 23259 31949
rect 23201 31940 23213 31943
rect 17819 31912 20300 31940
rect 20364 31912 23213 31940
rect 17819 31909 17831 31912
rect 17773 31903 17831 31909
rect 8260 31844 9435 31872
rect 8260 31832 8266 31844
rect 5077 31807 5135 31813
rect 5077 31773 5089 31807
rect 5123 31804 5135 31807
rect 6089 31807 6147 31813
rect 6089 31804 6101 31807
rect 5123 31776 6101 31804
rect 5123 31773 5135 31776
rect 5077 31767 5135 31773
rect 6089 31773 6101 31776
rect 6135 31773 6147 31807
rect 6365 31807 6440 31813
rect 6089 31767 6147 31773
rect 6265 31785 6323 31791
rect 6265 31751 6277 31785
rect 6311 31751 6323 31785
rect 6365 31773 6377 31807
rect 6411 31773 6440 31807
rect 6365 31770 6440 31773
rect 6365 31767 6423 31770
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 6641 31807 6699 31813
rect 6641 31773 6653 31807
rect 6687 31804 6699 31807
rect 7006 31804 7012 31816
rect 6687 31776 7012 31804
rect 6687 31773 6699 31776
rect 6641 31767 6699 31773
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 7098 31764 7104 31816
rect 7156 31764 7162 31816
rect 7285 31807 7343 31813
rect 7285 31773 7297 31807
rect 7331 31804 7343 31807
rect 7484 31804 7512 31832
rect 7331 31776 7512 31804
rect 7331 31773 7343 31776
rect 7285 31767 7343 31773
rect 8754 31764 8760 31816
rect 8812 31804 8818 31816
rect 9309 31807 9367 31813
rect 9309 31804 9321 31807
rect 8812 31776 9321 31804
rect 8812 31764 8818 31776
rect 9309 31773 9321 31776
rect 9355 31773 9367 31807
rect 9407 31804 9435 31844
rect 9600 31844 10456 31872
rect 10505 31875 10563 31881
rect 9600 31813 9628 31844
rect 10505 31841 10517 31875
rect 10551 31841 10563 31875
rect 11974 31872 11980 31884
rect 10505 31835 10563 31841
rect 10704 31844 11980 31872
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 9407 31776 9505 31804
rect 9309 31767 9367 31773
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 9585 31807 9643 31813
rect 9585 31773 9597 31807
rect 9631 31773 9643 31807
rect 9585 31767 9643 31773
rect 6265 31748 6323 31751
rect 4985 31739 5043 31745
rect 4985 31705 4997 31739
rect 5031 31736 5043 31739
rect 5350 31736 5356 31748
rect 5031 31708 5356 31736
rect 5031 31705 5043 31708
rect 4985 31699 5043 31705
rect 5350 31696 5356 31708
rect 5408 31696 5414 31748
rect 6265 31745 6276 31748
rect 6270 31696 6276 31745
rect 6328 31736 6334 31748
rect 7193 31739 7251 31745
rect 7193 31736 7205 31739
rect 6328 31708 7205 31736
rect 6328 31696 6334 31708
rect 7193 31705 7205 31708
rect 7239 31705 7251 31739
rect 9508 31736 9536 31767
rect 9858 31764 9864 31816
rect 9916 31804 9922 31816
rect 10321 31807 10379 31813
rect 10321 31804 10333 31807
rect 9916 31776 10333 31804
rect 9916 31764 9922 31776
rect 10321 31773 10333 31776
rect 10367 31773 10379 31807
rect 10321 31767 10379 31773
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 10704 31736 10732 31844
rect 11974 31832 11980 31844
rect 12032 31872 12038 31884
rect 13173 31875 13231 31881
rect 13173 31872 13185 31875
rect 12032 31844 13185 31872
rect 12032 31832 12038 31844
rect 12360 31813 12388 31844
rect 13173 31841 13185 31844
rect 13219 31841 13231 31875
rect 14182 31872 14188 31884
rect 13173 31835 13231 31841
rect 13648 31844 14188 31872
rect 12345 31807 12403 31813
rect 12345 31773 12357 31807
rect 12391 31804 12403 31807
rect 13449 31807 13507 31813
rect 12391 31776 12425 31804
rect 12391 31773 12403 31776
rect 12345 31767 12403 31773
rect 13449 31773 13461 31807
rect 13495 31798 13507 31807
rect 13648 31804 13676 31844
rect 14182 31832 14188 31844
rect 14240 31832 14246 31884
rect 14274 31832 14280 31884
rect 14332 31832 14338 31884
rect 14550 31813 14556 31816
rect 14544 31804 14556 31813
rect 13556 31798 13676 31804
rect 13495 31776 13676 31798
rect 14511 31776 14556 31804
rect 13495 31773 13584 31776
rect 13449 31770 13584 31773
rect 13449 31767 13507 31770
rect 14544 31767 14556 31776
rect 14550 31764 14556 31767
rect 14608 31764 14614 31816
rect 16393 31807 16451 31813
rect 16393 31773 16405 31807
rect 16439 31804 16451 31807
rect 18138 31804 18144 31816
rect 16439 31776 18144 31804
rect 16439 31773 16451 31776
rect 16393 31767 16451 31773
rect 18138 31764 18144 31776
rect 18196 31764 18202 31816
rect 20272 31813 20300 31912
rect 23201 31909 23213 31912
rect 23247 31909 23259 31943
rect 23201 31903 23259 31909
rect 25130 31900 25136 31952
rect 25188 31940 25194 31952
rect 26234 31940 26240 31952
rect 25188 31912 26240 31940
rect 25188 31900 25194 31912
rect 26234 31900 26240 31912
rect 26292 31900 26298 31952
rect 23382 31832 23388 31884
rect 23440 31832 23446 31884
rect 27154 31832 27160 31884
rect 27212 31872 27218 31884
rect 28644 31881 28672 31980
rect 30834 31968 30840 31980
rect 30892 31968 30898 32020
rect 31202 31968 31208 32020
rect 31260 32008 31266 32020
rect 32309 32011 32367 32017
rect 32309 32008 32321 32011
rect 31260 31980 32321 32008
rect 31260 31968 31266 31980
rect 32309 31977 32321 31980
rect 32355 32008 32367 32011
rect 35250 32008 35256 32020
rect 32355 31980 35256 32008
rect 32355 31977 32367 31980
rect 32309 31971 32367 31977
rect 35250 31968 35256 31980
rect 35308 31968 35314 32020
rect 35894 31968 35900 32020
rect 35952 31968 35958 32020
rect 36078 31968 36084 32020
rect 36136 32008 36142 32020
rect 36538 32008 36544 32020
rect 36136 31980 36544 32008
rect 36136 31968 36142 31980
rect 36538 31968 36544 31980
rect 36596 31968 36602 32020
rect 37458 31968 37464 32020
rect 37516 31968 37522 32020
rect 40954 31968 40960 32020
rect 41012 31968 41018 32020
rect 41782 32008 41788 32020
rect 41524 31980 41788 32008
rect 33134 31900 33140 31952
rect 33192 31940 33198 31952
rect 33192 31912 33272 31940
rect 33192 31900 33198 31912
rect 28629 31875 28687 31881
rect 28629 31872 28641 31875
rect 27212 31844 28641 31872
rect 27212 31832 27218 31844
rect 28629 31841 28641 31844
rect 28675 31841 28687 31875
rect 32490 31872 32496 31884
rect 28629 31835 28687 31841
rect 32416 31844 32496 31872
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31804 20683 31807
rect 20898 31804 20904 31816
rect 20671 31776 20904 31804
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31804 21143 31807
rect 21131 31776 21864 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 9508 31708 10732 31736
rect 7193 31699 7251 31705
rect 12434 31696 12440 31748
rect 12492 31736 12498 31748
rect 13630 31736 13636 31748
rect 12492 31708 13636 31736
rect 12492 31696 12498 31708
rect 13630 31696 13636 31708
rect 13688 31736 13694 31748
rect 16638 31739 16696 31745
rect 16638 31736 16650 31739
rect 13688 31708 16650 31736
rect 13688 31696 13694 31708
rect 16638 31705 16650 31708
rect 16684 31705 16696 31739
rect 16638 31699 16696 31705
rect 20990 31696 20996 31748
rect 21048 31736 21054 31748
rect 21729 31739 21787 31745
rect 21729 31736 21741 31739
rect 21048 31708 21741 31736
rect 21048 31696 21054 31708
rect 21729 31705 21741 31708
rect 21775 31705 21787 31739
rect 21836 31736 21864 31776
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22002 31764 22008 31816
rect 22060 31764 22066 31816
rect 22112 31776 23060 31804
rect 22112 31736 22140 31776
rect 21836 31708 22140 31736
rect 23032 31736 23060 31776
rect 23106 31764 23112 31816
rect 23164 31764 23170 31816
rect 23290 31764 23296 31816
rect 23348 31764 23354 31816
rect 23474 31804 23480 31816
rect 23400 31776 23480 31804
rect 23400 31736 23428 31776
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 23569 31807 23627 31813
rect 23569 31773 23581 31807
rect 23615 31804 23627 31807
rect 24670 31804 24676 31816
rect 23615 31776 24676 31804
rect 23615 31773 23627 31776
rect 23569 31767 23627 31773
rect 24670 31764 24676 31776
rect 24728 31764 24734 31816
rect 24854 31764 24860 31816
rect 24912 31804 24918 31816
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 24912 31776 24961 31804
rect 24912 31764 24918 31776
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25087 31807 25145 31813
rect 25087 31773 25099 31807
rect 25133 31804 25145 31807
rect 25222 31804 25228 31816
rect 25133 31776 25228 31804
rect 25133 31773 25145 31776
rect 25087 31767 25145 31773
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 25317 31807 25375 31813
rect 25317 31773 25329 31807
rect 25363 31804 25375 31807
rect 25866 31804 25872 31816
rect 25363 31776 25872 31804
rect 25363 31773 25375 31776
rect 25317 31767 25375 31773
rect 25866 31764 25872 31776
rect 25924 31764 25930 31816
rect 26050 31764 26056 31816
rect 26108 31804 26114 31816
rect 26145 31807 26203 31813
rect 26145 31804 26157 31807
rect 26108 31776 26157 31804
rect 26108 31764 26114 31776
rect 26145 31773 26157 31776
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 26234 31764 26240 31816
rect 26292 31804 26298 31816
rect 26789 31807 26847 31813
rect 26789 31804 26801 31807
rect 26292 31776 26801 31804
rect 26292 31764 26298 31776
rect 26789 31773 26801 31776
rect 26835 31773 26847 31807
rect 26789 31767 26847 31773
rect 26970 31764 26976 31816
rect 27028 31764 27034 31816
rect 27890 31764 27896 31816
rect 27948 31804 27954 31816
rect 27948 31776 28120 31804
rect 27948 31764 27954 31776
rect 23032 31708 23428 31736
rect 21729 31699 21787 31705
rect 25682 31696 25688 31748
rect 25740 31736 25746 31748
rect 25777 31739 25835 31745
rect 25777 31736 25789 31739
rect 25740 31708 25789 31736
rect 25740 31696 25746 31708
rect 25777 31705 25789 31708
rect 25823 31705 25835 31739
rect 26329 31739 26387 31745
rect 26329 31736 26341 31739
rect 25777 31699 25835 31705
rect 26252 31708 26341 31736
rect 26252 31680 26280 31708
rect 26329 31705 26341 31708
rect 26375 31736 26387 31739
rect 27062 31736 27068 31748
rect 26375 31708 27068 31736
rect 26375 31705 26387 31708
rect 26329 31699 26387 31705
rect 27062 31696 27068 31708
rect 27120 31696 27126 31748
rect 28092 31736 28120 31776
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28261 31807 28319 31813
rect 28261 31804 28273 31807
rect 28224 31776 28273 31804
rect 28224 31764 28230 31776
rect 28261 31773 28273 31776
rect 28307 31773 28319 31807
rect 28261 31767 28319 31773
rect 28442 31764 28448 31816
rect 28500 31764 28506 31816
rect 28534 31764 28540 31816
rect 28592 31764 28598 31816
rect 28813 31807 28871 31813
rect 28813 31804 28825 31807
rect 28736 31776 28825 31804
rect 28736 31736 28764 31776
rect 28813 31773 28825 31776
rect 28859 31773 28871 31807
rect 28813 31767 28871 31773
rect 29730 31764 29736 31816
rect 29788 31764 29794 31816
rect 29822 31764 29828 31816
rect 29880 31804 29886 31816
rect 29917 31807 29975 31813
rect 29917 31804 29929 31807
rect 29880 31776 29929 31804
rect 29880 31764 29886 31776
rect 29917 31773 29929 31776
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 32416 31813 32444 31844
rect 32490 31832 32496 31844
rect 32548 31872 32554 31884
rect 33244 31872 33272 31912
rect 33502 31900 33508 31952
rect 33560 31900 33566 31952
rect 34790 31900 34796 31952
rect 34848 31940 34854 31952
rect 35434 31940 35440 31952
rect 34848 31912 35440 31940
rect 34848 31900 34854 31912
rect 35434 31900 35440 31912
rect 35492 31900 35498 31952
rect 35710 31900 35716 31952
rect 35768 31900 35774 31952
rect 36630 31940 36636 31952
rect 35820 31912 36636 31940
rect 33367 31875 33425 31881
rect 33367 31872 33379 31875
rect 32548 31844 33180 31872
rect 33244 31844 33379 31872
rect 32548 31832 32554 31844
rect 31297 31807 31355 31813
rect 31297 31804 31309 31807
rect 31076 31776 31309 31804
rect 31076 31764 31082 31776
rect 31297 31773 31309 31776
rect 31343 31773 31355 31807
rect 31297 31767 31355 31773
rect 32401 31807 32459 31813
rect 32401 31773 32413 31807
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 28092 31708 28764 31736
rect 33152 31736 33180 31844
rect 33367 31841 33379 31844
rect 33413 31841 33425 31875
rect 35728 31872 35756 31900
rect 33367 31835 33425 31841
rect 35636 31844 35756 31872
rect 33226 31764 33232 31816
rect 33284 31764 33290 31816
rect 33597 31807 33655 31813
rect 33597 31773 33609 31807
rect 33643 31804 33655 31807
rect 33686 31804 33692 31816
rect 33643 31776 33692 31804
rect 33643 31773 33655 31776
rect 33597 31767 33655 31773
rect 33686 31764 33692 31776
rect 33744 31764 33750 31816
rect 35158 31764 35164 31816
rect 35216 31804 35222 31816
rect 35636 31813 35664 31844
rect 35253 31807 35311 31813
rect 35253 31804 35265 31807
rect 35216 31776 35265 31804
rect 35216 31764 35222 31776
rect 35253 31773 35265 31776
rect 35299 31773 35311 31807
rect 35253 31767 35311 31773
rect 35401 31807 35459 31813
rect 35401 31773 35413 31807
rect 35447 31773 35459 31807
rect 35401 31767 35459 31773
rect 35529 31807 35587 31813
rect 35529 31773 35541 31807
rect 35575 31773 35587 31807
rect 35529 31767 35587 31773
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31773 35679 31807
rect 35621 31767 35679 31773
rect 35718 31807 35776 31813
rect 35718 31773 35730 31807
rect 35764 31804 35776 31807
rect 35820 31804 35848 31912
rect 36630 31900 36636 31912
rect 36688 31900 36694 31952
rect 36354 31872 36360 31884
rect 35764 31776 35848 31804
rect 35912 31844 36360 31872
rect 35764 31773 35776 31776
rect 35718 31767 35776 31773
rect 33318 31736 33324 31748
rect 33152 31708 33324 31736
rect 33318 31696 33324 31708
rect 33376 31696 33382 31748
rect 8294 31628 8300 31680
rect 8352 31668 8358 31680
rect 9125 31671 9183 31677
rect 9125 31668 9137 31671
rect 8352 31640 9137 31668
rect 8352 31628 8358 31640
rect 9125 31637 9137 31640
rect 9171 31637 9183 31671
rect 9125 31631 9183 31637
rect 9214 31628 9220 31680
rect 9272 31668 9278 31680
rect 10318 31668 10324 31680
rect 9272 31640 10324 31668
rect 9272 31628 9278 31640
rect 10318 31628 10324 31640
rect 10376 31628 10382 31680
rect 10686 31628 10692 31680
rect 10744 31668 10750 31680
rect 10781 31671 10839 31677
rect 10781 31668 10793 31671
rect 10744 31640 10793 31668
rect 10744 31628 10750 31640
rect 10781 31637 10793 31640
rect 10827 31637 10839 31671
rect 10781 31631 10839 31637
rect 11422 31628 11428 31680
rect 11480 31668 11486 31680
rect 13814 31668 13820 31680
rect 11480 31640 13820 31668
rect 11480 31628 11486 31640
rect 13814 31628 13820 31640
rect 13872 31628 13878 31680
rect 22922 31628 22928 31680
rect 22980 31628 22986 31680
rect 24946 31628 24952 31680
rect 25004 31668 25010 31680
rect 25225 31671 25283 31677
rect 25225 31668 25237 31671
rect 25004 31640 25237 31668
rect 25004 31628 25010 31640
rect 25225 31637 25237 31640
rect 25271 31668 25283 31671
rect 25314 31668 25320 31680
rect 25271 31640 25320 31668
rect 25271 31637 25283 31640
rect 25225 31631 25283 31637
rect 25314 31628 25320 31640
rect 25372 31628 25378 31680
rect 26234 31628 26240 31680
rect 26292 31628 26298 31680
rect 28994 31628 29000 31680
rect 29052 31628 29058 31680
rect 29086 31628 29092 31680
rect 29144 31668 29150 31680
rect 29825 31671 29883 31677
rect 29825 31668 29837 31671
rect 29144 31640 29837 31668
rect 29144 31628 29150 31640
rect 29825 31637 29837 31640
rect 29871 31637 29883 31671
rect 35416 31668 35444 31767
rect 35544 31736 35572 31767
rect 35912 31736 35940 31844
rect 36354 31832 36360 31844
rect 36412 31872 36418 31884
rect 37090 31872 37096 31884
rect 36412 31844 37096 31872
rect 36412 31832 36418 31844
rect 37090 31832 37096 31844
rect 37148 31872 37154 31884
rect 37921 31875 37979 31881
rect 37921 31872 37933 31875
rect 37148 31844 37933 31872
rect 37148 31832 37154 31844
rect 37921 31841 37933 31844
rect 37967 31841 37979 31875
rect 37921 31835 37979 31841
rect 38102 31832 38108 31884
rect 38160 31872 38166 31884
rect 40034 31872 40040 31884
rect 38160 31844 40040 31872
rect 38160 31832 38166 31844
rect 40034 31832 40040 31844
rect 40092 31832 40098 31884
rect 41524 31881 41552 31980
rect 41782 31968 41788 31980
rect 41840 31968 41846 32020
rect 42889 31943 42947 31949
rect 42889 31940 42901 31943
rect 42720 31912 42901 31940
rect 41509 31875 41567 31881
rect 40512 31844 41414 31872
rect 35986 31764 35992 31816
rect 36044 31804 36050 31816
rect 36817 31807 36875 31813
rect 36817 31804 36829 31807
rect 36044 31776 36829 31804
rect 36044 31764 36050 31776
rect 36817 31773 36829 31776
rect 36863 31773 36875 31807
rect 36817 31767 36875 31773
rect 36906 31764 36912 31816
rect 36964 31764 36970 31816
rect 37282 31807 37340 31813
rect 37282 31804 37294 31807
rect 37016 31776 37294 31804
rect 35544 31708 35940 31736
rect 36630 31696 36636 31748
rect 36688 31736 36694 31748
rect 37016 31736 37044 31776
rect 37282 31773 37294 31776
rect 37328 31773 37340 31807
rect 37282 31767 37340 31773
rect 37550 31764 37556 31816
rect 37608 31804 37614 31816
rect 38289 31807 38347 31813
rect 38289 31804 38301 31807
rect 37608 31776 38301 31804
rect 37608 31764 37614 31776
rect 38289 31773 38301 31776
rect 38335 31773 38347 31807
rect 38289 31767 38347 31773
rect 38470 31764 38476 31816
rect 38528 31764 38534 31816
rect 38654 31764 38660 31816
rect 38712 31804 38718 31816
rect 40313 31807 40371 31813
rect 40313 31804 40325 31807
rect 38712 31776 40325 31804
rect 38712 31764 38718 31776
rect 40313 31773 40325 31776
rect 40359 31773 40371 31807
rect 40313 31767 40371 31773
rect 40402 31764 40408 31816
rect 40460 31804 40466 31816
rect 40512 31804 40540 31844
rect 40460 31776 40540 31804
rect 40819 31807 40877 31813
rect 40460 31764 40466 31776
rect 40819 31773 40831 31807
rect 40865 31804 40877 31807
rect 41386 31804 41414 31844
rect 41509 31841 41521 31875
rect 41555 31841 41567 31875
rect 41509 31835 41567 31841
rect 41776 31807 41834 31813
rect 40865 31776 41092 31804
rect 41386 31776 41736 31804
rect 40865 31773 40877 31776
rect 40819 31767 40877 31773
rect 41064 31748 41092 31776
rect 36688 31708 37044 31736
rect 36688 31696 36694 31708
rect 37090 31696 37096 31748
rect 37148 31696 37154 31748
rect 37185 31739 37243 31745
rect 37185 31705 37197 31739
rect 37231 31705 37243 31739
rect 37185 31699 37243 31705
rect 35894 31668 35900 31680
rect 35416 31640 35900 31668
rect 29825 31631 29883 31637
rect 35894 31628 35900 31640
rect 35952 31628 35958 31680
rect 35986 31628 35992 31680
rect 36044 31668 36050 31680
rect 37200 31668 37228 31699
rect 37458 31696 37464 31748
rect 37516 31736 37522 31748
rect 38010 31736 38016 31748
rect 37516 31708 38016 31736
rect 37516 31696 37522 31708
rect 38010 31696 38016 31708
rect 38068 31696 38074 31748
rect 38562 31696 38568 31748
rect 38620 31736 38626 31748
rect 38746 31736 38752 31748
rect 38620 31708 38752 31736
rect 38620 31696 38626 31708
rect 38746 31696 38752 31708
rect 38804 31696 38810 31748
rect 39574 31696 39580 31748
rect 39632 31736 39638 31748
rect 40586 31736 40592 31748
rect 39632 31708 40592 31736
rect 39632 31696 39638 31708
rect 40586 31696 40592 31708
rect 40644 31696 40650 31748
rect 40681 31739 40739 31745
rect 40681 31705 40693 31739
rect 40727 31736 40739 31739
rect 40727 31708 40816 31736
rect 40727 31705 40739 31708
rect 40681 31699 40739 31705
rect 40788 31680 40816 31708
rect 41046 31696 41052 31748
rect 41104 31696 41110 31748
rect 41708 31736 41736 31776
rect 41776 31773 41788 31807
rect 41822 31804 41834 31807
rect 42610 31804 42616 31816
rect 41822 31776 42616 31804
rect 41822 31773 41834 31776
rect 41776 31767 41834 31773
rect 42610 31764 42616 31776
rect 42668 31764 42674 31816
rect 42720 31736 42748 31912
rect 42889 31909 42901 31912
rect 42935 31940 42947 31943
rect 42978 31940 42984 31952
rect 42935 31912 42984 31940
rect 42935 31909 42947 31912
rect 42889 31903 42947 31909
rect 42978 31900 42984 31912
rect 43036 31900 43042 31952
rect 41708 31708 42748 31736
rect 39298 31668 39304 31680
rect 36044 31640 39304 31668
rect 36044 31628 36050 31640
rect 39298 31628 39304 31640
rect 39356 31628 39362 31680
rect 40770 31628 40776 31680
rect 40828 31628 40834 31680
rect 1104 31578 43884 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 43884 31578
rect 1104 31504 43884 31526
rect 6917 31467 6975 31473
rect 6917 31433 6929 31467
rect 6963 31464 6975 31467
rect 7558 31464 7564 31476
rect 6963 31436 7564 31464
rect 6963 31433 6975 31436
rect 6917 31427 6975 31433
rect 7558 31424 7564 31436
rect 7616 31424 7622 31476
rect 9306 31424 9312 31476
rect 9364 31464 9370 31476
rect 9401 31467 9459 31473
rect 9401 31464 9413 31467
rect 9364 31436 9413 31464
rect 9364 31424 9370 31436
rect 9401 31433 9413 31436
rect 9447 31433 9459 31467
rect 9401 31427 9459 31433
rect 9490 31424 9496 31476
rect 9548 31424 9554 31476
rect 10226 31464 10232 31476
rect 9600 31436 10232 31464
rect 8018 31396 8024 31408
rect 6840 31368 8024 31396
rect 6840 31337 6868 31368
rect 8018 31356 8024 31368
rect 8076 31356 8082 31408
rect 8665 31399 8723 31405
rect 8665 31365 8677 31399
rect 8711 31396 8723 31399
rect 9214 31396 9220 31408
rect 8711 31368 9220 31396
rect 8711 31365 8723 31368
rect 8665 31359 8723 31365
rect 9214 31356 9220 31368
rect 9272 31356 9278 31408
rect 6825 31331 6883 31337
rect 6825 31297 6837 31331
rect 6871 31297 6883 31331
rect 6825 31291 6883 31297
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31328 7159 31331
rect 7282 31328 7288 31340
rect 7147 31300 7288 31328
rect 7147 31297 7159 31300
rect 7101 31291 7159 31297
rect 7282 31288 7288 31300
rect 7340 31288 7346 31340
rect 8205 31331 8263 31337
rect 8205 31297 8217 31331
rect 8251 31297 8263 31331
rect 8205 31291 8263 31297
rect 7190 31220 7196 31272
rect 7248 31260 7254 31272
rect 8220 31260 8248 31291
rect 8294 31288 8300 31340
rect 8352 31288 8358 31340
rect 8481 31331 8539 31337
rect 8481 31297 8493 31331
rect 8527 31297 8539 31331
rect 8481 31291 8539 31297
rect 7248 31232 8248 31260
rect 8496 31260 8524 31291
rect 9306 31288 9312 31340
rect 9364 31328 9370 31340
rect 9600 31328 9628 31436
rect 10226 31424 10232 31436
rect 10284 31464 10290 31476
rect 10284 31436 10456 31464
rect 10284 31424 10290 31436
rect 10428 31396 10456 31436
rect 10594 31424 10600 31476
rect 10652 31464 10658 31476
rect 10781 31467 10839 31473
rect 10781 31464 10793 31467
rect 10652 31436 10793 31464
rect 10652 31424 10658 31436
rect 10781 31433 10793 31436
rect 10827 31433 10839 31467
rect 13354 31464 13360 31476
rect 10781 31427 10839 31433
rect 12820 31436 13360 31464
rect 11977 31399 12035 31405
rect 11977 31396 11989 31399
rect 9364 31300 9628 31328
rect 10060 31368 10364 31396
rect 10428 31368 11989 31396
rect 9364 31288 9370 31300
rect 10060 31260 10088 31368
rect 10336 31337 10364 31368
rect 11977 31365 11989 31368
rect 12023 31365 12035 31399
rect 11977 31359 12035 31365
rect 10137 31331 10195 31337
rect 10137 31297 10149 31331
rect 10183 31297 10195 31331
rect 10137 31291 10195 31297
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 8496 31232 10088 31260
rect 7248 31220 7254 31232
rect 6178 31152 6184 31204
rect 6236 31192 6242 31204
rect 6236 31164 8248 31192
rect 6236 31152 6242 31164
rect 7190 31084 7196 31136
rect 7248 31124 7254 31136
rect 7285 31127 7343 31133
rect 7285 31124 7297 31127
rect 7248 31096 7297 31124
rect 7248 31084 7254 31096
rect 7285 31093 7297 31096
rect 7331 31093 7343 31127
rect 7285 31087 7343 31093
rect 8110 31084 8116 31136
rect 8168 31124 8174 31136
rect 8220 31124 8248 31164
rect 8294 31152 8300 31204
rect 8352 31192 8358 31204
rect 8389 31195 8447 31201
rect 8389 31192 8401 31195
rect 8352 31164 8401 31192
rect 8352 31152 8358 31164
rect 8389 31161 8401 31164
rect 8435 31161 8447 31195
rect 8389 31155 8447 31161
rect 8496 31124 8524 31232
rect 8662 31152 8668 31204
rect 8720 31192 8726 31204
rect 9125 31195 9183 31201
rect 9125 31192 9137 31195
rect 8720 31164 9137 31192
rect 8720 31152 8726 31164
rect 9125 31161 9137 31164
rect 9171 31192 9183 31195
rect 9858 31192 9864 31204
rect 9171 31164 9864 31192
rect 9171 31161 9183 31164
rect 9125 31155 9183 31161
rect 9858 31152 9864 31164
rect 9916 31192 9922 31204
rect 10152 31192 10180 31291
rect 10336 31260 10364 31291
rect 10410 31288 10416 31340
rect 10468 31288 10474 31340
rect 10502 31288 10508 31340
rect 10560 31288 10566 31340
rect 11698 31288 11704 31340
rect 11756 31288 11762 31340
rect 12713 31331 12771 31337
rect 12713 31297 12725 31331
rect 12759 31328 12771 31331
rect 12820 31328 12848 31436
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 19978 31424 19984 31476
rect 20036 31464 20042 31476
rect 32306 31464 32312 31476
rect 20036 31436 32312 31464
rect 20036 31424 20042 31436
rect 32306 31424 32312 31436
rect 32364 31424 32370 31476
rect 34146 31424 34152 31476
rect 34204 31424 34210 31476
rect 34330 31424 34336 31476
rect 34388 31464 34394 31476
rect 34388 31436 36216 31464
rect 34388 31424 34394 31436
rect 13725 31399 13783 31405
rect 13725 31396 13737 31399
rect 12912 31368 13737 31396
rect 12912 31337 12940 31368
rect 13725 31365 13737 31368
rect 13771 31365 13783 31399
rect 13725 31359 13783 31365
rect 13906 31356 13912 31408
rect 13964 31405 13970 31408
rect 13964 31399 13983 31405
rect 13971 31365 13983 31399
rect 13964 31359 13983 31365
rect 13964 31356 13970 31359
rect 23106 31356 23112 31408
rect 23164 31396 23170 31408
rect 25685 31399 25743 31405
rect 23164 31368 23980 31396
rect 23164 31356 23170 31368
rect 12759 31300 12848 31328
rect 12897 31331 12955 31337
rect 12759 31297 12771 31300
rect 12713 31291 12771 31297
rect 12897 31297 12909 31331
rect 12943 31297 12955 31331
rect 12897 31291 12955 31297
rect 11422 31260 11428 31272
rect 10336 31232 11428 31260
rect 11422 31220 11428 31232
rect 11480 31220 11486 31272
rect 12912 31192 12940 31291
rect 18230 31288 18236 31340
rect 18288 31328 18294 31340
rect 19061 31331 19119 31337
rect 19061 31328 19073 31331
rect 18288 31300 19073 31328
rect 18288 31288 18294 31300
rect 19061 31297 19073 31300
rect 19107 31297 19119 31331
rect 19061 31291 19119 31297
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 23017 31331 23075 31337
rect 23017 31328 23029 31331
rect 22980 31300 23029 31328
rect 22980 31288 22986 31300
rect 23017 31297 23029 31300
rect 23063 31297 23075 31331
rect 23017 31291 23075 31297
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31328 23351 31331
rect 23842 31328 23848 31340
rect 23339 31300 23848 31328
rect 23339 31297 23351 31300
rect 23293 31291 23351 31297
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 23952 31337 23980 31368
rect 25685 31365 25697 31399
rect 25731 31396 25743 31399
rect 25731 31368 29960 31396
rect 25731 31365 25743 31368
rect 25685 31359 25743 31365
rect 23937 31331 23995 31337
rect 23937 31297 23949 31331
rect 23983 31297 23995 31331
rect 23937 31291 23995 31297
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 23109 31263 23167 31269
rect 23109 31229 23121 31263
rect 23155 31260 23167 31263
rect 24854 31260 24860 31272
rect 23155 31232 24860 31260
rect 23155 31229 23167 31232
rect 23109 31223 23167 31229
rect 24854 31220 24860 31232
rect 24912 31220 24918 31272
rect 9916 31164 12940 31192
rect 23201 31195 23259 31201
rect 9916 31152 9922 31164
rect 23201 31161 23213 31195
rect 23247 31161 23259 31195
rect 23201 31155 23259 31161
rect 23477 31195 23535 31201
rect 23477 31161 23489 31195
rect 23523 31192 23535 31195
rect 24486 31192 24492 31204
rect 23523 31164 24492 31192
rect 23523 31161 23535 31164
rect 23477 31155 23535 31161
rect 8168 31096 8524 31124
rect 9677 31127 9735 31133
rect 8168 31084 8174 31096
rect 9677 31093 9689 31127
rect 9723 31124 9735 31127
rect 10686 31124 10692 31136
rect 9723 31096 10692 31124
rect 9723 31093 9735 31096
rect 9677 31087 9735 31093
rect 10686 31084 10692 31096
rect 10744 31084 10750 31136
rect 12713 31127 12771 31133
rect 12713 31093 12725 31127
rect 12759 31124 12771 31127
rect 12802 31124 12808 31136
rect 12759 31096 12808 31124
rect 12759 31093 12771 31096
rect 12713 31087 12771 31093
rect 12802 31084 12808 31096
rect 12860 31084 12866 31136
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 13909 31127 13967 31133
rect 13909 31124 13921 31127
rect 13872 31096 13921 31124
rect 13872 31084 13878 31096
rect 13909 31093 13921 31096
rect 13955 31093 13967 31127
rect 13909 31087 13967 31093
rect 14093 31127 14151 31133
rect 14093 31093 14105 31127
rect 14139 31124 14151 31127
rect 15010 31124 15016 31136
rect 14139 31096 15016 31124
rect 14139 31093 14151 31096
rect 14093 31087 14151 31093
rect 15010 31084 15016 31096
rect 15068 31084 15074 31136
rect 19153 31127 19211 31133
rect 19153 31093 19165 31127
rect 19199 31124 19211 31127
rect 19334 31124 19340 31136
rect 19199 31096 19340 31124
rect 19199 31093 19211 31096
rect 19153 31087 19211 31093
rect 19334 31084 19340 31096
rect 19392 31084 19398 31136
rect 23216 31124 23244 31155
rect 24486 31152 24492 31164
rect 24544 31152 24550 31204
rect 25240 31192 25268 31291
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 26605 31331 26663 31337
rect 26605 31297 26617 31331
rect 26651 31328 26663 31331
rect 26970 31328 26976 31340
rect 26651 31300 26976 31328
rect 26651 31297 26663 31300
rect 26605 31291 26663 31297
rect 26970 31288 26976 31300
rect 27028 31288 27034 31340
rect 28074 31288 28080 31340
rect 28132 31288 28138 31340
rect 28258 31288 28264 31340
rect 28316 31328 28322 31340
rect 28445 31331 28503 31337
rect 28445 31328 28457 31331
rect 28316 31300 28457 31328
rect 28316 31288 28322 31300
rect 28445 31297 28457 31300
rect 28491 31297 28503 31331
rect 29932 31328 29960 31368
rect 30006 31356 30012 31408
rect 30064 31396 30070 31408
rect 30650 31396 30656 31408
rect 30064 31368 30656 31396
rect 30064 31356 30070 31368
rect 30650 31356 30656 31368
rect 30708 31396 30714 31408
rect 32585 31399 32643 31405
rect 30708 31368 31064 31396
rect 30708 31356 30714 31368
rect 30098 31328 30104 31340
rect 29932 31300 30104 31328
rect 28445 31291 28503 31297
rect 30098 31288 30104 31300
rect 30156 31288 30162 31340
rect 30834 31288 30840 31340
rect 30892 31288 30898 31340
rect 31036 31337 31064 31368
rect 32585 31365 32597 31399
rect 32631 31396 32643 31399
rect 33410 31396 33416 31408
rect 32631 31368 33416 31396
rect 32631 31365 32643 31368
rect 32585 31359 32643 31365
rect 33410 31356 33416 31368
rect 33468 31356 33474 31408
rect 34422 31356 34428 31408
rect 34480 31396 34486 31408
rect 36078 31396 36084 31408
rect 34480 31368 36084 31396
rect 34480 31356 34486 31368
rect 36078 31356 36084 31368
rect 36136 31356 36142 31408
rect 31021 31331 31079 31337
rect 31021 31297 31033 31331
rect 31067 31297 31079 31331
rect 31021 31291 31079 31297
rect 32398 31288 32404 31340
rect 32456 31288 32462 31340
rect 33318 31288 33324 31340
rect 33376 31288 33382 31340
rect 34238 31288 34244 31340
rect 34296 31288 34302 31340
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 35222 31331 35280 31337
rect 35222 31328 35234 31331
rect 34756 31300 35234 31328
rect 34756 31288 34762 31300
rect 35222 31297 35234 31300
rect 35268 31297 35280 31331
rect 35222 31291 35280 31297
rect 35345 31331 35403 31337
rect 35345 31297 35357 31331
rect 35391 31297 35403 31331
rect 35986 31328 35992 31340
rect 35345 31291 35403 31297
rect 35636 31300 35992 31328
rect 26418 31220 26424 31272
rect 26476 31220 26482 31272
rect 26510 31220 26516 31272
rect 26568 31260 26574 31272
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 26568 31232 27721 31260
rect 26568 31220 26574 31232
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 32769 31263 32827 31269
rect 32769 31229 32781 31263
rect 32815 31260 32827 31263
rect 32950 31260 32956 31272
rect 32815 31232 32956 31260
rect 32815 31229 32827 31232
rect 32769 31223 32827 31229
rect 32950 31220 32956 31232
rect 33008 31260 33014 31272
rect 35360 31260 35388 31291
rect 33008 31232 35388 31260
rect 33008 31220 33014 31232
rect 35434 31220 35440 31272
rect 35492 31260 35498 31272
rect 35636 31269 35664 31300
rect 35986 31288 35992 31300
rect 36044 31288 36050 31340
rect 35621 31263 35679 31269
rect 35621 31260 35633 31263
rect 35492 31232 35633 31260
rect 35492 31220 35498 31232
rect 35621 31229 35633 31232
rect 35667 31229 35679 31263
rect 35621 31223 35679 31229
rect 35713 31263 35771 31269
rect 35713 31229 35725 31263
rect 35759 31229 35771 31263
rect 36188 31260 36216 31436
rect 38010 31424 38016 31476
rect 38068 31464 38074 31476
rect 38473 31467 38531 31473
rect 38068 31436 38424 31464
rect 38068 31424 38074 31436
rect 38396 31396 38424 31436
rect 38473 31433 38485 31467
rect 38519 31464 38531 31467
rect 38654 31464 38660 31476
rect 38519 31436 38660 31464
rect 38519 31433 38531 31436
rect 38473 31427 38531 31433
rect 38654 31424 38660 31436
rect 38712 31424 38718 31476
rect 41046 31424 41052 31476
rect 41104 31424 41110 31476
rect 38746 31396 38752 31408
rect 36372 31368 38332 31396
rect 38396 31368 38752 31396
rect 36372 31337 36400 31368
rect 36357 31331 36415 31337
rect 36357 31297 36369 31331
rect 36403 31297 36415 31331
rect 36357 31291 36415 31297
rect 36446 31288 36452 31340
rect 36504 31288 36510 31340
rect 36538 31288 36544 31340
rect 36596 31337 36602 31340
rect 36596 31331 36645 31337
rect 36596 31297 36599 31331
rect 36633 31297 36645 31331
rect 36596 31291 36645 31297
rect 36725 31331 36783 31337
rect 36725 31297 36737 31331
rect 36771 31297 36783 31331
rect 36725 31291 36783 31297
rect 36596 31288 36602 31291
rect 36464 31260 36492 31288
rect 36188 31232 36492 31260
rect 35713 31223 35771 31229
rect 29362 31192 29368 31204
rect 25240 31164 29368 31192
rect 29362 31152 29368 31164
rect 29420 31152 29426 31204
rect 30006 31152 30012 31204
rect 30064 31192 30070 31204
rect 30064 31164 31754 31192
rect 30064 31152 30070 31164
rect 23566 31124 23572 31136
rect 23216 31096 23572 31124
rect 23566 31084 23572 31096
rect 23624 31084 23630 31136
rect 23658 31084 23664 31136
rect 23716 31124 23722 31136
rect 24029 31127 24087 31133
rect 24029 31124 24041 31127
rect 23716 31096 24041 31124
rect 23716 31084 23722 31096
rect 24029 31093 24041 31096
rect 24075 31093 24087 31127
rect 24029 31087 24087 31093
rect 24118 31084 24124 31136
rect 24176 31124 24182 31136
rect 25041 31127 25099 31133
rect 25041 31124 25053 31127
rect 24176 31096 25053 31124
rect 24176 31084 24182 31096
rect 25041 31093 25053 31096
rect 25087 31093 25099 31127
rect 25041 31087 25099 31093
rect 25222 31084 25228 31136
rect 25280 31084 25286 31136
rect 26418 31084 26424 31136
rect 26476 31124 26482 31136
rect 27062 31124 27068 31136
rect 26476 31096 27068 31124
rect 26476 31084 26482 31096
rect 27062 31084 27068 31096
rect 27120 31084 27126 31136
rect 31110 31084 31116 31136
rect 31168 31084 31174 31136
rect 31726 31124 31754 31164
rect 35342 31152 35348 31204
rect 35400 31192 35406 31204
rect 35728 31192 35756 31223
rect 35802 31192 35808 31204
rect 35400 31164 35808 31192
rect 35400 31152 35406 31164
rect 35802 31152 35808 31164
rect 35860 31152 35866 31204
rect 35894 31152 35900 31204
rect 35952 31192 35958 31204
rect 36630 31192 36636 31204
rect 35952 31164 36636 31192
rect 35952 31152 35958 31164
rect 36630 31152 36636 31164
rect 36688 31192 36694 31204
rect 36740 31192 36768 31291
rect 37274 31288 37280 31340
rect 37332 31328 37338 31340
rect 37332 31300 37872 31328
rect 37332 31288 37338 31300
rect 37844 31260 37872 31300
rect 37918 31288 37924 31340
rect 37976 31288 37982 31340
rect 38010 31288 38016 31340
rect 38068 31328 38074 31340
rect 38304 31337 38332 31368
rect 38746 31356 38752 31368
rect 38804 31356 38810 31408
rect 38105 31331 38163 31337
rect 38105 31328 38117 31331
rect 38068 31300 38117 31328
rect 38068 31288 38074 31300
rect 38105 31297 38117 31300
rect 38151 31297 38163 31331
rect 38105 31291 38163 31297
rect 38197 31331 38255 31337
rect 38197 31297 38209 31331
rect 38243 31297 38255 31331
rect 38197 31291 38255 31297
rect 38289 31331 38347 31337
rect 38289 31297 38301 31331
rect 38335 31328 38347 31331
rect 39114 31328 39120 31340
rect 38335 31300 39120 31328
rect 38335 31297 38347 31300
rect 38289 31291 38347 31297
rect 38212 31260 38240 31291
rect 39114 31288 39120 31300
rect 39172 31328 39178 31340
rect 39390 31328 39396 31340
rect 39172 31300 39396 31328
rect 39172 31288 39178 31300
rect 39390 31288 39396 31300
rect 39448 31288 39454 31340
rect 39482 31288 39488 31340
rect 39540 31328 39546 31340
rect 40865 31331 40923 31337
rect 40865 31328 40877 31331
rect 39540 31300 40877 31328
rect 39540 31288 39546 31300
rect 40865 31297 40877 31300
rect 40911 31297 40923 31331
rect 40865 31291 40923 31297
rect 42889 31331 42947 31337
rect 42889 31297 42901 31331
rect 42935 31328 42947 31331
rect 43070 31328 43076 31340
rect 42935 31300 43076 31328
rect 42935 31297 42947 31300
rect 42889 31291 42947 31297
rect 43070 31288 43076 31300
rect 43128 31288 43134 31340
rect 37844 31232 38240 31260
rect 38838 31220 38844 31272
rect 38896 31260 38902 31272
rect 39206 31260 39212 31272
rect 38896 31232 39212 31260
rect 38896 31220 38902 31232
rect 39206 31220 39212 31232
rect 39264 31220 39270 31272
rect 43162 31220 43168 31272
rect 43220 31220 43226 31272
rect 36688 31164 36768 31192
rect 36688 31152 36694 31164
rect 34330 31124 34336 31136
rect 31726 31096 34336 31124
rect 34330 31084 34336 31096
rect 34388 31084 34394 31136
rect 34514 31084 34520 31136
rect 34572 31124 34578 31136
rect 35069 31127 35127 31133
rect 35069 31124 35081 31127
rect 34572 31096 35081 31124
rect 34572 31084 34578 31096
rect 35069 31093 35081 31096
rect 35115 31093 35127 31127
rect 35069 31087 35127 31093
rect 36078 31084 36084 31136
rect 36136 31124 36142 31136
rect 36173 31127 36231 31133
rect 36173 31124 36185 31127
rect 36136 31096 36185 31124
rect 36136 31084 36142 31096
rect 36173 31093 36185 31096
rect 36219 31093 36231 31127
rect 36173 31087 36231 31093
rect 36906 31084 36912 31136
rect 36964 31124 36970 31136
rect 38746 31124 38752 31136
rect 36964 31096 38752 31124
rect 36964 31084 36970 31096
rect 38746 31084 38752 31096
rect 38804 31124 38810 31136
rect 39206 31124 39212 31136
rect 38804 31096 39212 31124
rect 38804 31084 38810 31096
rect 39206 31084 39212 31096
rect 39264 31084 39270 31136
rect 1104 31034 43884 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 43884 31034
rect 1104 30960 43884 30982
rect 7006 30880 7012 30932
rect 7064 30880 7070 30932
rect 7282 30880 7288 30932
rect 7340 30920 7346 30932
rect 7377 30923 7435 30929
rect 7377 30920 7389 30923
rect 7340 30892 7389 30920
rect 7340 30880 7346 30892
rect 7377 30889 7389 30892
rect 7423 30889 7435 30923
rect 7377 30883 7435 30889
rect 7466 30880 7472 30932
rect 7524 30920 7530 30932
rect 20254 30920 20260 30932
rect 7524 30892 20260 30920
rect 7524 30880 7530 30892
rect 20254 30880 20260 30892
rect 20312 30880 20318 30932
rect 23566 30880 23572 30932
rect 23624 30920 23630 30932
rect 24946 30920 24952 30932
rect 23624 30892 24952 30920
rect 23624 30880 23630 30892
rect 24946 30880 24952 30892
rect 25004 30880 25010 30932
rect 25041 30923 25099 30929
rect 25041 30889 25053 30923
rect 25087 30920 25099 30923
rect 25130 30920 25136 30932
rect 25087 30892 25136 30920
rect 25087 30889 25099 30892
rect 25041 30883 25099 30889
rect 25130 30880 25136 30892
rect 25188 30880 25194 30932
rect 25406 30880 25412 30932
rect 25464 30920 25470 30932
rect 25464 30892 27844 30920
rect 25464 30880 25470 30892
rect 4614 30812 4620 30864
rect 4672 30852 4678 30864
rect 19705 30855 19763 30861
rect 4672 30824 11652 30852
rect 4672 30812 4678 30824
rect 5445 30787 5503 30793
rect 5445 30753 5457 30787
rect 5491 30784 5503 30787
rect 6454 30784 6460 30796
rect 5491 30756 6460 30784
rect 5491 30753 5503 30756
rect 5445 30747 5503 30753
rect 6454 30744 6460 30756
rect 6512 30784 6518 30796
rect 7374 30784 7380 30796
rect 6512 30756 7380 30784
rect 6512 30744 6518 30756
rect 7374 30744 7380 30756
rect 7432 30744 7438 30796
rect 7469 30787 7527 30793
rect 7469 30753 7481 30787
rect 7515 30784 7527 30787
rect 8294 30784 8300 30796
rect 7515 30756 8300 30784
rect 7515 30753 7527 30756
rect 7469 30747 7527 30753
rect 8294 30744 8300 30756
rect 8352 30744 8358 30796
rect 9490 30744 9496 30796
rect 9548 30784 9554 30796
rect 9677 30787 9735 30793
rect 9677 30784 9689 30787
rect 9548 30756 9689 30784
rect 9548 30744 9554 30756
rect 9677 30753 9689 30756
rect 9723 30753 9735 30787
rect 9677 30747 9735 30753
rect 5261 30719 5319 30725
rect 5261 30685 5273 30719
rect 5307 30716 5319 30719
rect 6270 30716 6276 30728
rect 5307 30688 6276 30716
rect 5307 30685 5319 30688
rect 5261 30679 5319 30685
rect 6270 30676 6276 30688
rect 6328 30676 6334 30728
rect 7098 30676 7104 30728
rect 7156 30716 7162 30728
rect 7193 30719 7251 30725
rect 7193 30716 7205 30719
rect 7156 30688 7205 30716
rect 7156 30676 7162 30688
rect 7193 30685 7205 30688
rect 7239 30685 7251 30719
rect 7193 30679 7251 30685
rect 8110 30676 8116 30728
rect 8168 30676 8174 30728
rect 8202 30676 8208 30728
rect 8260 30676 8266 30728
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30716 8447 30719
rect 8754 30716 8760 30728
rect 8435 30688 8760 30716
rect 8435 30685 8447 30688
rect 8389 30679 8447 30685
rect 8754 30676 8760 30688
rect 8812 30676 8818 30728
rect 7558 30608 7564 30660
rect 7616 30648 7622 30660
rect 9692 30648 9720 30747
rect 9766 30744 9772 30796
rect 9824 30784 9830 30796
rect 10410 30784 10416 30796
rect 9824 30756 10416 30784
rect 9824 30744 9830 30756
rect 10410 30744 10416 30756
rect 10468 30744 10474 30796
rect 10778 30744 10784 30796
rect 10836 30744 10842 30796
rect 11624 30793 11652 30824
rect 19705 30821 19717 30855
rect 19751 30852 19763 30855
rect 19978 30852 19984 30864
rect 19751 30824 19984 30852
rect 19751 30821 19763 30824
rect 19705 30815 19763 30821
rect 19978 30812 19984 30824
rect 20036 30812 20042 30864
rect 24118 30852 24124 30864
rect 20916 30824 24124 30852
rect 11609 30787 11667 30793
rect 11609 30753 11621 30787
rect 11655 30753 11667 30787
rect 11609 30747 11667 30753
rect 9858 30676 9864 30728
rect 9916 30676 9922 30728
rect 9953 30719 10011 30725
rect 9953 30685 9965 30719
rect 9999 30716 10011 30719
rect 10502 30716 10508 30728
rect 9999 30688 10508 30716
rect 9999 30685 10011 30688
rect 9953 30679 10011 30685
rect 10502 30676 10508 30688
rect 10560 30676 10566 30728
rect 10597 30719 10655 30725
rect 10597 30685 10609 30719
rect 10643 30716 10655 30719
rect 10796 30716 10824 30744
rect 10643 30688 10824 30716
rect 10643 30685 10655 30688
rect 10597 30679 10655 30685
rect 10962 30676 10968 30728
rect 11020 30676 11026 30728
rect 11514 30716 11520 30728
rect 11072 30688 11520 30716
rect 7616 30620 9720 30648
rect 7616 30608 7622 30620
rect 10686 30608 10692 30660
rect 10744 30648 10750 30660
rect 10781 30651 10839 30657
rect 10781 30648 10793 30651
rect 10744 30620 10793 30648
rect 10744 30608 10750 30620
rect 10781 30617 10793 30620
rect 10827 30617 10839 30651
rect 10781 30611 10839 30617
rect 10873 30651 10931 30657
rect 10873 30617 10885 30651
rect 10919 30648 10931 30651
rect 11072 30648 11100 30688
rect 11514 30676 11520 30688
rect 11572 30676 11578 30728
rect 11624 30716 11652 30747
rect 17586 30744 17592 30796
rect 17644 30784 17650 30796
rect 17865 30787 17923 30793
rect 17865 30784 17877 30787
rect 17644 30756 17877 30784
rect 17644 30744 17650 30756
rect 17865 30753 17877 30756
rect 17911 30753 17923 30787
rect 17865 30747 17923 30753
rect 18322 30744 18328 30796
rect 18380 30744 18386 30796
rect 20916 30784 20944 30824
rect 24118 30812 24124 30824
rect 24176 30812 24182 30864
rect 24673 30855 24731 30861
rect 24673 30821 24685 30855
rect 24719 30852 24731 30855
rect 25222 30852 25228 30864
rect 24719 30824 25228 30852
rect 24719 30821 24731 30824
rect 24673 30815 24731 30821
rect 25222 30812 25228 30824
rect 25280 30812 25286 30864
rect 26694 30812 26700 30864
rect 26752 30852 26758 30864
rect 26752 30824 27752 30852
rect 26752 30812 26758 30824
rect 19720 30756 20944 30784
rect 21361 30787 21419 30793
rect 12158 30716 12164 30728
rect 11624 30688 12164 30716
rect 12158 30676 12164 30688
rect 12216 30716 12222 30728
rect 14274 30716 14280 30728
rect 12216 30688 14280 30716
rect 12216 30676 12222 30688
rect 14274 30676 14280 30688
rect 14332 30716 14338 30728
rect 14553 30719 14611 30725
rect 14553 30716 14565 30719
rect 14332 30688 14565 30716
rect 14332 30676 14338 30688
rect 14553 30685 14565 30688
rect 14599 30685 14611 30719
rect 14553 30679 14611 30685
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18340 30716 18368 30744
rect 18003 30688 18368 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 19426 30676 19432 30728
rect 19484 30676 19490 30728
rect 19720 30725 19748 30756
rect 21361 30753 21373 30787
rect 21407 30784 21419 30787
rect 22370 30784 22376 30796
rect 21407 30756 22376 30784
rect 21407 30753 21419 30756
rect 21361 30747 21419 30753
rect 22370 30744 22376 30756
rect 22428 30744 22434 30796
rect 23658 30744 23664 30796
rect 23716 30744 23722 30796
rect 23842 30744 23848 30796
rect 23900 30784 23906 30796
rect 25038 30784 25044 30796
rect 23900 30756 25044 30784
rect 23900 30744 23906 30756
rect 25038 30744 25044 30756
rect 25096 30744 25102 30796
rect 25133 30787 25191 30793
rect 25133 30753 25145 30787
rect 25179 30784 25191 30787
rect 26418 30784 26424 30796
rect 25179 30756 26424 30784
rect 25179 30753 25191 30756
rect 25133 30747 25191 30753
rect 26418 30744 26424 30756
rect 26476 30744 26482 30796
rect 27430 30744 27436 30796
rect 27488 30784 27494 30796
rect 27724 30793 27752 30824
rect 27617 30787 27675 30793
rect 27617 30784 27629 30787
rect 27488 30756 27629 30784
rect 27488 30744 27494 30756
rect 27617 30753 27629 30756
rect 27663 30753 27675 30787
rect 27617 30747 27675 30753
rect 27709 30787 27767 30793
rect 27709 30753 27721 30787
rect 27755 30753 27767 30787
rect 27816 30784 27844 30892
rect 31570 30880 31576 30932
rect 31628 30920 31634 30932
rect 31628 30892 34928 30920
rect 31628 30880 31634 30892
rect 32950 30812 32956 30864
rect 33008 30852 33014 30864
rect 33045 30855 33103 30861
rect 33045 30852 33057 30855
rect 33008 30824 33057 30852
rect 33008 30812 33014 30824
rect 33045 30821 33057 30824
rect 33091 30821 33103 30855
rect 33045 30815 33103 30821
rect 33502 30812 33508 30864
rect 33560 30852 33566 30864
rect 33778 30852 33784 30864
rect 33560 30824 33784 30852
rect 33560 30812 33566 30824
rect 33778 30812 33784 30824
rect 33836 30812 33842 30864
rect 33965 30855 34023 30861
rect 33965 30821 33977 30855
rect 34011 30821 34023 30855
rect 33965 30815 34023 30821
rect 28445 30787 28503 30793
rect 28445 30784 28457 30787
rect 27816 30756 28457 30784
rect 27709 30747 27767 30753
rect 28445 30753 28457 30756
rect 28491 30784 28503 30787
rect 29270 30784 29276 30796
rect 28491 30756 29276 30784
rect 28491 30753 28503 30756
rect 28445 30747 28503 30753
rect 29270 30744 29276 30756
rect 29328 30744 29334 30796
rect 33980 30784 34008 30815
rect 32968 30756 34008 30784
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 20254 30676 20260 30728
rect 20312 30716 20318 30728
rect 20349 30719 20407 30725
rect 20349 30716 20361 30719
rect 20312 30688 20361 30716
rect 20312 30676 20318 30688
rect 20349 30685 20361 30688
rect 20395 30716 20407 30719
rect 20395 30688 20944 30716
rect 20395 30685 20407 30688
rect 20349 30679 20407 30685
rect 11854 30651 11912 30657
rect 11854 30648 11866 30651
rect 10919 30620 11100 30648
rect 11624 30620 11866 30648
rect 10919 30617 10931 30620
rect 10873 30611 10931 30617
rect 4798 30540 4804 30592
rect 4856 30540 4862 30592
rect 5169 30583 5227 30589
rect 5169 30549 5181 30583
rect 5215 30580 5227 30583
rect 5534 30580 5540 30592
rect 5215 30552 5540 30580
rect 5215 30549 5227 30552
rect 5169 30543 5227 30549
rect 5534 30540 5540 30552
rect 5592 30540 5598 30592
rect 8570 30540 8576 30592
rect 8628 30540 8634 30592
rect 9490 30540 9496 30592
rect 9548 30540 9554 30592
rect 11149 30583 11207 30589
rect 11149 30549 11161 30583
rect 11195 30580 11207 30583
rect 11624 30580 11652 30620
rect 11854 30617 11866 30620
rect 11900 30617 11912 30651
rect 11854 30611 11912 30617
rect 14642 30608 14648 30660
rect 14700 30648 14706 30660
rect 14798 30651 14856 30657
rect 14798 30648 14810 30651
rect 14700 30620 14810 30648
rect 14700 30608 14706 30620
rect 14798 30617 14810 30620
rect 14844 30617 14856 30651
rect 14798 30611 14856 30617
rect 18230 30608 18236 30660
rect 18288 30608 18294 30660
rect 18325 30651 18383 30657
rect 18325 30617 18337 30651
rect 18371 30648 18383 30651
rect 20162 30648 20168 30660
rect 18371 30620 20168 30648
rect 18371 30617 18383 30620
rect 18325 30611 18383 30617
rect 20162 30608 20168 30620
rect 20220 30608 20226 30660
rect 20806 30608 20812 30660
rect 20864 30608 20870 30660
rect 20916 30648 20944 30688
rect 20990 30676 20996 30728
rect 21048 30676 21054 30728
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30716 24915 30719
rect 25406 30716 25412 30728
rect 24903 30688 25412 30716
rect 24903 30685 24915 30688
rect 24857 30679 24915 30685
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 25866 30676 25872 30728
rect 25924 30676 25930 30728
rect 26145 30719 26203 30725
rect 26145 30685 26157 30719
rect 26191 30716 26203 30719
rect 26234 30716 26240 30728
rect 26191 30688 26240 30716
rect 26191 30685 26203 30688
rect 26145 30679 26203 30685
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 26970 30676 26976 30728
rect 27028 30716 27034 30728
rect 27341 30719 27399 30725
rect 27341 30716 27353 30719
rect 27028 30688 27353 30716
rect 27028 30676 27034 30688
rect 27341 30685 27353 30688
rect 27387 30685 27399 30719
rect 28721 30719 28779 30725
rect 27341 30679 27399 30685
rect 27448 30688 28488 30716
rect 27448 30648 27476 30688
rect 28460 30660 28488 30688
rect 28721 30685 28733 30719
rect 28767 30716 28779 30719
rect 28994 30716 29000 30728
rect 28767 30688 29000 30716
rect 28767 30685 28779 30688
rect 28721 30679 28779 30685
rect 28994 30676 29000 30688
rect 29052 30676 29058 30728
rect 30650 30676 30656 30728
rect 30708 30676 30714 30728
rect 30834 30676 30840 30728
rect 30892 30716 30898 30728
rect 32968 30725 32996 30756
rect 31297 30719 31355 30725
rect 31297 30716 31309 30719
rect 30892 30688 31309 30716
rect 30892 30676 30898 30688
rect 31297 30685 31309 30688
rect 31343 30685 31355 30719
rect 31297 30679 31355 30685
rect 32953 30719 33011 30725
rect 32953 30685 32965 30719
rect 32999 30685 33011 30719
rect 32953 30679 33011 30685
rect 33134 30676 33140 30728
rect 33192 30676 33198 30728
rect 33229 30719 33287 30725
rect 33229 30685 33241 30719
rect 33275 30716 33287 30719
rect 33686 30716 33692 30728
rect 33275 30688 33692 30716
rect 33275 30685 33287 30688
rect 33229 30679 33287 30685
rect 33686 30676 33692 30688
rect 33744 30676 33750 30728
rect 34238 30676 34244 30728
rect 34296 30676 34302 30728
rect 34900 30725 34928 30892
rect 36262 30880 36268 30932
rect 36320 30920 36326 30932
rect 36998 30920 37004 30932
rect 36320 30892 37004 30920
rect 36320 30880 36326 30892
rect 36998 30880 37004 30892
rect 37056 30880 37062 30932
rect 37550 30880 37556 30932
rect 37608 30920 37614 30932
rect 38930 30920 38936 30932
rect 37608 30892 38936 30920
rect 37608 30880 37614 30892
rect 38930 30880 38936 30892
rect 38988 30880 38994 30932
rect 39206 30880 39212 30932
rect 39264 30920 39270 30932
rect 42978 30920 42984 30932
rect 39264 30892 42984 30920
rect 39264 30880 39270 30892
rect 42978 30880 42984 30892
rect 43036 30920 43042 30932
rect 43257 30923 43315 30929
rect 43257 30920 43269 30923
rect 43036 30892 43269 30920
rect 43036 30880 43042 30892
rect 43257 30889 43269 30892
rect 43303 30889 43315 30923
rect 43257 30883 43315 30889
rect 36538 30852 36544 30864
rect 35636 30824 36544 30852
rect 35636 30793 35664 30824
rect 36538 30812 36544 30824
rect 36596 30852 36602 30864
rect 36596 30824 38654 30852
rect 36596 30812 36602 30824
rect 35621 30787 35679 30793
rect 35621 30753 35633 30787
rect 35667 30753 35679 30787
rect 35621 30747 35679 30753
rect 37458 30744 37464 30796
rect 37516 30784 37522 30796
rect 38626 30784 38654 30824
rect 39574 30784 39580 30796
rect 37516 30756 38516 30784
rect 38626 30756 39580 30784
rect 37516 30744 37522 30756
rect 34885 30719 34943 30725
rect 34885 30685 34897 30719
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 34974 30676 34980 30728
rect 35032 30676 35038 30728
rect 35158 30676 35164 30728
rect 35216 30676 35222 30728
rect 36078 30676 36084 30728
rect 36136 30676 36142 30728
rect 36170 30676 36176 30728
rect 36228 30676 36234 30728
rect 36354 30676 36360 30728
rect 36412 30676 36418 30728
rect 36449 30719 36507 30725
rect 36449 30685 36461 30719
rect 36495 30716 36507 30719
rect 37550 30716 37556 30728
rect 36495 30688 37556 30716
rect 36495 30685 36507 30688
rect 36449 30679 36507 30685
rect 37550 30676 37556 30688
rect 37608 30676 37614 30728
rect 37737 30719 37795 30725
rect 37737 30685 37749 30719
rect 37783 30716 37795 30719
rect 38378 30716 38384 30728
rect 37783 30688 38384 30716
rect 37783 30685 37795 30688
rect 37737 30679 37795 30685
rect 38378 30676 38384 30688
rect 38436 30676 38442 30728
rect 20916 30620 27476 30648
rect 27826 30651 27884 30657
rect 27826 30617 27838 30651
rect 27872 30648 27884 30651
rect 27872 30620 28304 30648
rect 27872 30617 27884 30620
rect 27826 30611 27884 30617
rect 11195 30552 11652 30580
rect 11195 30549 11207 30552
rect 11149 30543 11207 30549
rect 11698 30540 11704 30592
rect 11756 30580 11762 30592
rect 12989 30583 13047 30589
rect 12989 30580 13001 30583
rect 11756 30552 13001 30580
rect 11756 30540 11762 30552
rect 12989 30549 13001 30552
rect 13035 30580 13047 30583
rect 14458 30580 14464 30592
rect 13035 30552 14464 30580
rect 13035 30549 13047 30552
rect 12989 30543 13047 30549
rect 14458 30540 14464 30552
rect 14516 30540 14522 30592
rect 15930 30540 15936 30592
rect 15988 30540 15994 30592
rect 17586 30540 17592 30592
rect 17644 30580 17650 30592
rect 17681 30583 17739 30589
rect 17681 30580 17693 30583
rect 17644 30552 17693 30580
rect 17644 30540 17650 30552
rect 17681 30549 17693 30552
rect 17727 30549 17739 30583
rect 17681 30543 17739 30549
rect 18874 30540 18880 30592
rect 18932 30580 18938 30592
rect 19521 30583 19579 30589
rect 19521 30580 19533 30583
rect 18932 30552 19533 30580
rect 18932 30540 18938 30552
rect 19521 30549 19533 30552
rect 19567 30549 19579 30583
rect 19521 30543 19579 30549
rect 20254 30540 20260 30592
rect 20312 30540 20318 30592
rect 23198 30540 23204 30592
rect 23256 30540 23262 30592
rect 23566 30540 23572 30592
rect 23624 30540 23630 30592
rect 24854 30540 24860 30592
rect 24912 30580 24918 30592
rect 25685 30583 25743 30589
rect 25685 30580 25697 30583
rect 24912 30552 25697 30580
rect 24912 30540 24918 30552
rect 25685 30549 25697 30552
rect 25731 30549 25743 30583
rect 25685 30543 25743 30549
rect 27982 30540 27988 30592
rect 28040 30540 28046 30592
rect 28276 30580 28304 30620
rect 28442 30608 28448 30660
rect 28500 30608 28506 30660
rect 28813 30651 28871 30657
rect 28813 30617 28825 30651
rect 28859 30648 28871 30651
rect 29086 30648 29092 30660
rect 28859 30620 29092 30648
rect 28859 30617 28871 30620
rect 28813 30611 28871 30617
rect 29086 30608 29092 30620
rect 29144 30608 29150 30660
rect 29181 30651 29239 30657
rect 29181 30617 29193 30651
rect 29227 30648 29239 30651
rect 30926 30648 30932 30660
rect 29227 30620 30932 30648
rect 29227 30617 29239 30620
rect 29181 30611 29239 30617
rect 30926 30608 30932 30620
rect 30984 30608 30990 30660
rect 32306 30608 32312 30660
rect 32364 30648 32370 30660
rect 32364 30620 33548 30648
rect 32364 30608 32370 30620
rect 28626 30580 28632 30592
rect 28276 30552 28632 30580
rect 28626 30540 28632 30552
rect 28684 30540 28690 30592
rect 31478 30540 31484 30592
rect 31536 30540 31542 30592
rect 33410 30540 33416 30592
rect 33468 30540 33474 30592
rect 33520 30580 33548 30620
rect 33962 30608 33968 30660
rect 34020 30608 34026 30660
rect 37369 30651 37427 30657
rect 37369 30617 37381 30651
rect 37415 30648 37427 30651
rect 38102 30648 38108 30660
rect 37415 30620 38108 30648
rect 37415 30617 37427 30620
rect 37369 30611 37427 30617
rect 38102 30608 38108 30620
rect 38160 30608 38166 30660
rect 38488 30648 38516 30756
rect 38746 30676 38752 30728
rect 38804 30676 38810 30728
rect 38948 30725 38976 30756
rect 39574 30744 39580 30756
rect 39632 30744 39638 30796
rect 40034 30744 40040 30796
rect 40092 30744 40098 30796
rect 40129 30787 40187 30793
rect 40129 30753 40141 30787
rect 40175 30784 40187 30787
rect 40402 30784 40408 30796
rect 40175 30756 40408 30784
rect 40175 30753 40187 30756
rect 40129 30747 40187 30753
rect 40402 30744 40408 30756
rect 40460 30744 40466 30796
rect 41690 30744 41696 30796
rect 41748 30784 41754 30796
rect 41877 30787 41935 30793
rect 41877 30784 41889 30787
rect 41748 30756 41889 30784
rect 41748 30744 41754 30756
rect 41877 30753 41889 30756
rect 41923 30753 41935 30787
rect 41877 30747 41935 30753
rect 38933 30719 38991 30725
rect 38933 30685 38945 30719
rect 38979 30685 38991 30719
rect 38933 30679 38991 30685
rect 39114 30676 39120 30728
rect 39172 30676 39178 30728
rect 40218 30676 40224 30728
rect 40276 30716 40282 30728
rect 40313 30719 40371 30725
rect 40313 30716 40325 30719
rect 40276 30688 40325 30716
rect 40276 30676 40282 30688
rect 40313 30685 40325 30688
rect 40359 30685 40371 30719
rect 40313 30679 40371 30685
rect 39025 30651 39083 30657
rect 39025 30648 39037 30651
rect 38488 30620 39037 30648
rect 39025 30617 39037 30620
rect 39071 30617 39083 30651
rect 39025 30611 39083 30617
rect 42144 30651 42202 30657
rect 42144 30617 42156 30651
rect 42190 30648 42202 30651
rect 42610 30648 42616 30660
rect 42190 30620 42616 30648
rect 42190 30617 42202 30620
rect 42144 30611 42202 30617
rect 42610 30608 42616 30620
rect 42668 30608 42674 30660
rect 34149 30583 34207 30589
rect 34149 30580 34161 30583
rect 33520 30552 34161 30580
rect 34149 30549 34161 30552
rect 34195 30549 34207 30583
rect 34149 30543 34207 30549
rect 36633 30583 36691 30589
rect 36633 30549 36645 30583
rect 36679 30580 36691 30583
rect 37918 30580 37924 30592
rect 36679 30552 37924 30580
rect 36679 30549 36691 30552
rect 36633 30543 36691 30549
rect 37918 30540 37924 30552
rect 37976 30540 37982 30592
rect 39206 30540 39212 30592
rect 39264 30580 39270 30592
rect 39301 30583 39359 30589
rect 39301 30580 39313 30583
rect 39264 30552 39313 30580
rect 39264 30540 39270 30552
rect 39301 30549 39313 30552
rect 39347 30549 39359 30583
rect 39301 30543 39359 30549
rect 40497 30583 40555 30589
rect 40497 30549 40509 30583
rect 40543 30580 40555 30583
rect 43070 30580 43076 30592
rect 40543 30552 43076 30580
rect 40543 30549 40555 30552
rect 40497 30543 40555 30549
rect 43070 30540 43076 30552
rect 43128 30540 43134 30592
rect 1104 30490 43884 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 43884 30490
rect 1104 30416 43884 30438
rect 5534 30336 5540 30388
rect 5592 30376 5598 30388
rect 7466 30376 7472 30388
rect 5592 30348 7472 30376
rect 5592 30336 5598 30348
rect 7466 30336 7472 30348
rect 7524 30336 7530 30388
rect 14553 30379 14611 30385
rect 14553 30345 14565 30379
rect 14599 30376 14611 30379
rect 14642 30376 14648 30388
rect 14599 30348 14648 30376
rect 14599 30345 14611 30348
rect 14553 30339 14611 30345
rect 14642 30336 14648 30348
rect 14700 30336 14706 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 20073 30379 20131 30385
rect 20073 30376 20085 30379
rect 19484 30348 20085 30376
rect 19484 30336 19490 30348
rect 20073 30345 20085 30348
rect 20119 30345 20131 30379
rect 20073 30339 20131 30345
rect 20806 30336 20812 30388
rect 20864 30376 20870 30388
rect 20864 30348 22140 30376
rect 20864 30336 20870 30348
rect 4614 30308 4620 30320
rect 4172 30280 4620 30308
rect 4172 30249 4200 30280
rect 4614 30268 4620 30280
rect 4672 30268 4678 30320
rect 9398 30268 9404 30320
rect 9456 30308 9462 30320
rect 9493 30311 9551 30317
rect 9493 30308 9505 30311
rect 9456 30280 9505 30308
rect 9456 30268 9462 30280
rect 9493 30277 9505 30280
rect 9539 30277 9551 30311
rect 9493 30271 9551 30277
rect 13814 30268 13820 30320
rect 13872 30308 13878 30320
rect 14185 30311 14243 30317
rect 14185 30308 14197 30311
rect 13872 30280 14197 30308
rect 13872 30268 13878 30280
rect 14185 30277 14197 30280
rect 14231 30277 14243 30311
rect 14185 30271 14243 30277
rect 14458 30268 14464 30320
rect 14516 30308 14522 30320
rect 14516 30280 18828 30308
rect 14516 30268 14522 30280
rect 4157 30243 4215 30249
rect 4157 30209 4169 30243
rect 4203 30209 4215 30243
rect 4157 30203 4215 30209
rect 4424 30243 4482 30249
rect 4424 30209 4436 30243
rect 4470 30240 4482 30243
rect 4798 30240 4804 30252
rect 4470 30212 4804 30240
rect 4470 30209 4482 30212
rect 4424 30203 4482 30209
rect 4798 30200 4804 30212
rect 4856 30200 4862 30252
rect 9585 30243 9643 30249
rect 9585 30209 9597 30243
rect 9631 30240 9643 30243
rect 9766 30240 9772 30252
rect 9631 30212 9772 30240
rect 9631 30209 9643 30212
rect 9585 30203 9643 30209
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 10686 30200 10692 30252
rect 10744 30240 10750 30252
rect 10873 30243 10931 30249
rect 10873 30240 10885 30243
rect 10744 30212 10885 30240
rect 10744 30200 10750 30212
rect 10873 30209 10885 30212
rect 10919 30209 10931 30243
rect 10873 30203 10931 30209
rect 11057 30243 11115 30249
rect 11057 30209 11069 30243
rect 11103 30209 11115 30243
rect 11057 30203 11115 30209
rect 11072 30172 11100 30203
rect 11146 30200 11152 30252
rect 11204 30200 11210 30252
rect 12342 30200 12348 30252
rect 12400 30240 12406 30252
rect 12989 30243 13047 30249
rect 12989 30240 13001 30243
rect 12400 30212 13001 30240
rect 12400 30200 12406 30212
rect 12989 30209 13001 30212
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 13262 30200 13268 30252
rect 13320 30200 13326 30252
rect 13906 30200 13912 30252
rect 13964 30240 13970 30252
rect 14001 30243 14059 30249
rect 14001 30240 14013 30243
rect 13964 30212 14013 30240
rect 13964 30200 13970 30212
rect 14001 30209 14013 30212
rect 14047 30209 14059 30243
rect 14001 30203 14059 30209
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30209 14335 30243
rect 14277 30203 14335 30209
rect 11606 30172 11612 30184
rect 11072 30144 11612 30172
rect 11606 30132 11612 30144
rect 11664 30132 11670 30184
rect 14292 30172 14320 30203
rect 14366 30200 14372 30252
rect 14424 30200 14430 30252
rect 17954 30200 17960 30252
rect 18012 30200 18018 30252
rect 18800 30249 18828 30280
rect 18874 30268 18880 30320
rect 18932 30268 18938 30320
rect 19242 30268 19248 30320
rect 19300 30308 19306 30320
rect 22112 30308 22140 30348
rect 23566 30336 23572 30388
rect 23624 30376 23630 30388
rect 25774 30376 25780 30388
rect 23624 30348 25780 30376
rect 23624 30336 23630 30348
rect 25774 30336 25780 30348
rect 25832 30336 25838 30388
rect 29270 30336 29276 30388
rect 29328 30376 29334 30388
rect 29457 30379 29515 30385
rect 29457 30376 29469 30379
rect 29328 30348 29469 30376
rect 29328 30336 29334 30348
rect 29457 30345 29469 30348
rect 29503 30345 29515 30379
rect 29457 30339 29515 30345
rect 29546 30336 29552 30388
rect 29604 30376 29610 30388
rect 30282 30376 30288 30388
rect 29604 30348 30288 30376
rect 29604 30336 29610 30348
rect 30282 30336 30288 30348
rect 30340 30376 30346 30388
rect 30653 30379 30711 30385
rect 30653 30376 30665 30379
rect 30340 30348 30665 30376
rect 30340 30336 30346 30348
rect 30653 30345 30665 30348
rect 30699 30345 30711 30379
rect 30653 30339 30711 30345
rect 31110 30336 31116 30388
rect 31168 30376 31174 30388
rect 35710 30376 35716 30388
rect 31168 30348 32812 30376
rect 31168 30336 31174 30348
rect 19300 30280 22048 30308
rect 22112 30280 25728 30308
rect 19300 30268 19306 30280
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30240 18843 30243
rect 18966 30240 18972 30252
rect 18831 30212 18972 30240
rect 18831 30209 18843 30212
rect 18785 30203 18843 30209
rect 18966 30200 18972 30212
rect 19024 30200 19030 30252
rect 19587 30243 19645 30249
rect 19587 30209 19599 30243
rect 19633 30240 19645 30243
rect 19633 30209 19656 30240
rect 19587 30203 19656 30209
rect 15930 30172 15936 30184
rect 14292 30144 15936 30172
rect 15930 30132 15936 30144
rect 15988 30132 15994 30184
rect 17773 30175 17831 30181
rect 17773 30141 17785 30175
rect 17819 30172 17831 30175
rect 18414 30172 18420 30184
rect 17819 30144 18420 30172
rect 17819 30141 17831 30144
rect 17773 30135 17831 30141
rect 18414 30132 18420 30144
rect 18472 30132 18478 30184
rect 19429 30175 19487 30181
rect 19429 30141 19441 30175
rect 19475 30141 19487 30175
rect 19628 30172 19656 30203
rect 19702 30200 19708 30252
rect 19760 30200 19766 30252
rect 19794 30200 19800 30252
rect 19852 30200 19858 30252
rect 19889 30243 19947 30249
rect 19889 30209 19901 30243
rect 19935 30240 19947 30243
rect 20806 30240 20812 30252
rect 19935 30212 20812 30240
rect 19935 30209 19947 30212
rect 19889 30203 19947 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 21266 30200 21272 30252
rect 21324 30200 21330 30252
rect 21450 30200 21456 30252
rect 21508 30200 21514 30252
rect 22020 30249 22048 30280
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22261 30243 22319 30249
rect 22261 30240 22273 30243
rect 22005 30203 22063 30209
rect 22112 30212 22273 30240
rect 21085 30175 21143 30181
rect 19628 30144 19932 30172
rect 19429 30135 19487 30141
rect 13170 30064 13176 30116
rect 13228 30104 13234 30116
rect 13228 30076 18368 30104
rect 13228 30064 13234 30076
rect 10686 29996 10692 30048
rect 10744 29996 10750 30048
rect 11606 29996 11612 30048
rect 11664 30036 11670 30048
rect 18230 30036 18236 30048
rect 11664 30008 18236 30036
rect 11664 29996 11670 30008
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 18340 30036 18368 30076
rect 19242 30064 19248 30116
rect 19300 30104 19306 30116
rect 19444 30104 19472 30135
rect 19300 30076 19472 30104
rect 19300 30064 19306 30076
rect 19904 30048 19932 30144
rect 21085 30141 21097 30175
rect 21131 30172 21143 30175
rect 22112 30172 22140 30212
rect 22261 30209 22273 30212
rect 22307 30209 22319 30243
rect 22261 30203 22319 30209
rect 24302 30200 24308 30252
rect 24360 30200 24366 30252
rect 25038 30200 25044 30252
rect 25096 30240 25102 30252
rect 25133 30243 25191 30249
rect 25133 30240 25145 30243
rect 25096 30212 25145 30240
rect 25096 30200 25102 30212
rect 25133 30209 25145 30212
rect 25179 30209 25191 30243
rect 25133 30203 25191 30209
rect 21131 30144 22140 30172
rect 21131 30141 21143 30144
rect 21085 30135 21143 30141
rect 23566 30132 23572 30184
rect 23624 30172 23630 30184
rect 24397 30175 24455 30181
rect 24397 30172 24409 30175
rect 23624 30144 24409 30172
rect 23624 30132 23630 30144
rect 24397 30141 24409 30144
rect 24443 30141 24455 30175
rect 24397 30135 24455 30141
rect 24486 30132 24492 30184
rect 24544 30132 24550 30184
rect 23937 30107 23995 30113
rect 23937 30104 23949 30107
rect 22940 30076 23949 30104
rect 19794 30036 19800 30048
rect 18340 30008 19800 30036
rect 19794 29996 19800 30008
rect 19852 29996 19858 30048
rect 19886 29996 19892 30048
rect 19944 30036 19950 30048
rect 20990 30036 20996 30048
rect 19944 30008 20996 30036
rect 19944 29996 19950 30008
rect 20990 29996 20996 30008
rect 21048 29996 21054 30048
rect 21450 29996 21456 30048
rect 21508 30036 21514 30048
rect 22940 30036 22968 30076
rect 23937 30073 23949 30076
rect 23983 30073 23995 30107
rect 23937 30067 23995 30073
rect 24026 30064 24032 30116
rect 24084 30104 24090 30116
rect 25148 30104 25176 30203
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25590 30240 25596 30252
rect 25372 30212 25596 30240
rect 25372 30200 25378 30212
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 25700 30181 25728 30280
rect 25866 30268 25872 30320
rect 25924 30308 25930 30320
rect 25924 30280 26556 30308
rect 25924 30268 25930 30280
rect 26326 30200 26332 30252
rect 26384 30200 26390 30252
rect 26528 30249 26556 30280
rect 26620 30280 32720 30308
rect 26513 30243 26571 30249
rect 26513 30209 26525 30243
rect 26559 30209 26571 30243
rect 26513 30203 26571 30209
rect 25685 30175 25743 30181
rect 25685 30141 25697 30175
rect 25731 30172 25743 30175
rect 26620 30172 26648 30280
rect 28074 30200 28080 30252
rect 28132 30200 28138 30252
rect 28350 30200 28356 30252
rect 28408 30200 28414 30252
rect 28718 30200 28724 30252
rect 28776 30200 28782 30252
rect 29362 30200 29368 30252
rect 29420 30240 29426 30252
rect 29457 30243 29515 30249
rect 29457 30240 29469 30243
rect 29420 30212 29469 30240
rect 29420 30200 29426 30212
rect 29457 30209 29469 30212
rect 29503 30240 29515 30243
rect 29546 30240 29552 30252
rect 29503 30212 29552 30240
rect 29503 30209 29515 30212
rect 29457 30203 29515 30209
rect 29546 30200 29552 30212
rect 29604 30200 29610 30252
rect 29641 30243 29699 30249
rect 29641 30209 29653 30243
rect 29687 30209 29699 30243
rect 29641 30203 29699 30209
rect 28092 30172 28120 30200
rect 25731 30144 26648 30172
rect 27816 30144 28028 30172
rect 28092 30144 28580 30172
rect 25731 30141 25743 30144
rect 25685 30135 25743 30141
rect 26050 30104 26056 30116
rect 24084 30076 25084 30104
rect 25148 30076 26056 30104
rect 24084 30064 24090 30076
rect 21508 30008 22968 30036
rect 23385 30039 23443 30045
rect 21508 29996 21514 30008
rect 23385 30005 23397 30039
rect 23431 30036 23443 30039
rect 24302 30036 24308 30048
rect 23431 30008 24308 30036
rect 23431 30005 23443 30008
rect 23385 29999 23443 30005
rect 24302 29996 24308 30008
rect 24360 29996 24366 30048
rect 25056 30036 25084 30076
rect 26050 30064 26056 30076
rect 26108 30104 26114 30116
rect 26329 30107 26387 30113
rect 26329 30104 26341 30107
rect 26108 30076 26341 30104
rect 26108 30064 26114 30076
rect 26329 30073 26341 30076
rect 26375 30073 26387 30107
rect 26329 30067 26387 30073
rect 27816 30045 27844 30144
rect 28000 30104 28028 30144
rect 28258 30104 28264 30116
rect 28000 30076 28264 30104
rect 28258 30064 28264 30076
rect 28316 30064 28322 30116
rect 27801 30039 27859 30045
rect 27801 30036 27813 30039
rect 25056 30008 27813 30036
rect 27801 30005 27813 30008
rect 27847 30005 27859 30039
rect 28552 30036 28580 30144
rect 28718 30064 28724 30116
rect 28776 30104 28782 30116
rect 29656 30104 29684 30203
rect 30650 30200 30656 30252
rect 30708 30200 30714 30252
rect 31297 30243 31355 30249
rect 31297 30209 31309 30243
rect 31343 30240 31355 30243
rect 32398 30240 32404 30252
rect 31343 30212 32404 30240
rect 31343 30209 31355 30212
rect 31297 30203 31355 30209
rect 32398 30200 32404 30212
rect 32456 30200 32462 30252
rect 31573 30175 31631 30181
rect 31573 30141 31585 30175
rect 31619 30172 31631 30175
rect 31662 30172 31668 30184
rect 31619 30144 31668 30172
rect 31619 30141 31631 30144
rect 31573 30135 31631 30141
rect 31662 30132 31668 30144
rect 31720 30132 31726 30184
rect 32306 30132 32312 30184
rect 32364 30132 32370 30184
rect 28776 30076 29684 30104
rect 28776 30064 28782 30076
rect 30282 30064 30288 30116
rect 30340 30104 30346 30116
rect 32692 30104 32720 30280
rect 32784 30249 32812 30348
rect 35544 30348 35716 30376
rect 35158 30308 35164 30320
rect 34072 30280 35164 30308
rect 34072 30252 34100 30280
rect 35158 30268 35164 30280
rect 35216 30268 35222 30320
rect 32769 30243 32827 30249
rect 32769 30209 32781 30243
rect 32815 30209 32827 30243
rect 32769 30203 32827 30209
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30240 33655 30243
rect 34054 30240 34060 30252
rect 33643 30212 34060 30240
rect 33643 30209 33655 30212
rect 33597 30203 33655 30209
rect 34054 30200 34060 30212
rect 34112 30200 34118 30252
rect 34164 30212 34836 30240
rect 33137 30175 33195 30181
rect 33137 30141 33149 30175
rect 33183 30172 33195 30175
rect 34164 30172 34192 30212
rect 33183 30144 34192 30172
rect 34241 30175 34299 30181
rect 33183 30141 33195 30144
rect 33137 30135 33195 30141
rect 34241 30141 34253 30175
rect 34287 30172 34299 30175
rect 34514 30172 34520 30184
rect 34287 30144 34520 30172
rect 34287 30141 34299 30144
rect 34241 30135 34299 30141
rect 34514 30132 34520 30144
rect 34572 30132 34578 30184
rect 34808 30172 34836 30212
rect 34882 30200 34888 30252
rect 34940 30240 34946 30252
rect 34977 30243 35035 30249
rect 34977 30240 34989 30243
rect 34940 30212 34989 30240
rect 34940 30200 34946 30212
rect 34977 30209 34989 30212
rect 35023 30209 35035 30243
rect 34977 30203 35035 30209
rect 35434 30200 35440 30252
rect 35492 30200 35498 30252
rect 35544 30249 35572 30348
rect 35710 30336 35716 30348
rect 35768 30336 35774 30388
rect 35989 30379 36047 30385
rect 35989 30345 36001 30379
rect 36035 30376 36047 30379
rect 36170 30376 36176 30388
rect 36035 30348 36176 30376
rect 36035 30345 36047 30348
rect 35989 30339 36047 30345
rect 36170 30336 36176 30348
rect 36228 30336 36234 30388
rect 37826 30336 37832 30388
rect 37884 30376 37890 30388
rect 37884 30348 39344 30376
rect 37884 30336 37890 30348
rect 37844 30308 37872 30336
rect 39206 30308 39212 30320
rect 35820 30280 37872 30308
rect 39040 30280 39212 30308
rect 35820 30252 35848 30280
rect 35529 30243 35587 30249
rect 35529 30209 35541 30243
rect 35575 30209 35587 30243
rect 35529 30203 35587 30209
rect 35710 30200 35716 30252
rect 35768 30200 35774 30252
rect 35802 30200 35808 30252
rect 35860 30200 35866 30252
rect 36449 30243 36507 30249
rect 36449 30209 36461 30243
rect 36495 30209 36507 30243
rect 36449 30203 36507 30209
rect 35894 30172 35900 30184
rect 34808 30144 35900 30172
rect 35894 30132 35900 30144
rect 35952 30132 35958 30184
rect 34790 30104 34796 30116
rect 30340 30076 32628 30104
rect 32692 30076 34796 30104
rect 30340 30064 30346 30076
rect 30374 30036 30380 30048
rect 28552 30008 30380 30036
rect 27801 29999 27859 30005
rect 30374 29996 30380 30008
rect 30432 29996 30438 30048
rect 32600 30036 32628 30076
rect 34790 30064 34796 30076
rect 34848 30104 34854 30116
rect 34974 30104 34980 30116
rect 34848 30076 34980 30104
rect 34848 30064 34854 30076
rect 34974 30064 34980 30076
rect 35032 30064 35038 30116
rect 35526 30064 35532 30116
rect 35584 30104 35590 30116
rect 36464 30104 36492 30203
rect 36630 30200 36636 30252
rect 36688 30240 36694 30252
rect 39040 30249 39068 30280
rect 39206 30268 39212 30280
rect 39264 30268 39270 30320
rect 39316 30308 39344 30348
rect 42610 30336 42616 30388
rect 42668 30336 42674 30388
rect 42978 30336 42984 30388
rect 43036 30336 43042 30388
rect 43070 30336 43076 30388
rect 43128 30336 43134 30388
rect 39577 30311 39635 30317
rect 39316 30280 39436 30308
rect 37829 30243 37887 30249
rect 37829 30240 37841 30243
rect 36688 30212 37841 30240
rect 36688 30200 36694 30212
rect 37829 30209 37841 30212
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 39025 30243 39083 30249
rect 39025 30209 39037 30243
rect 39071 30209 39083 30243
rect 39025 30203 39083 30209
rect 39117 30243 39175 30249
rect 39117 30209 39129 30243
rect 39163 30209 39175 30243
rect 39117 30203 39175 30209
rect 36725 30175 36783 30181
rect 36725 30141 36737 30175
rect 36771 30172 36783 30175
rect 37274 30172 37280 30184
rect 36771 30144 37280 30172
rect 36771 30141 36783 30144
rect 36725 30135 36783 30141
rect 37274 30132 37280 30144
rect 37332 30132 37338 30184
rect 37918 30132 37924 30184
rect 37976 30132 37982 30184
rect 38102 30132 38108 30184
rect 38160 30132 38166 30184
rect 38930 30132 38936 30184
rect 38988 30172 38994 30184
rect 39132 30172 39160 30203
rect 39298 30200 39304 30252
rect 39356 30200 39362 30252
rect 39408 30249 39436 30280
rect 39577 30277 39589 30311
rect 39623 30308 39635 30311
rect 40218 30308 40224 30320
rect 39623 30280 40224 30308
rect 39623 30277 39635 30280
rect 39577 30271 39635 30277
rect 40218 30268 40224 30280
rect 40276 30268 40282 30320
rect 39393 30243 39451 30249
rect 39393 30209 39405 30243
rect 39439 30209 39451 30243
rect 39393 30203 39451 30209
rect 39942 30200 39948 30252
rect 40000 30240 40006 30252
rect 40000 30212 40264 30240
rect 40000 30200 40006 30212
rect 38988 30144 39160 30172
rect 38988 30132 38994 30144
rect 40126 30132 40132 30184
rect 40184 30132 40190 30184
rect 40236 30172 40264 30212
rect 40310 30200 40316 30252
rect 40368 30200 40374 30252
rect 40957 30243 41015 30249
rect 40957 30240 40969 30243
rect 40420 30212 40969 30240
rect 40420 30172 40448 30212
rect 40957 30209 40969 30212
rect 41003 30209 41015 30243
rect 40957 30203 41015 30209
rect 41141 30243 41199 30249
rect 41141 30209 41153 30243
rect 41187 30209 41199 30243
rect 41141 30203 41199 30209
rect 40236 30144 40448 30172
rect 40497 30175 40555 30181
rect 40497 30141 40509 30175
rect 40543 30172 40555 30175
rect 41156 30172 41184 30203
rect 40543 30144 41184 30172
rect 43165 30175 43223 30181
rect 40543 30141 40555 30144
rect 40497 30135 40555 30141
rect 43165 30141 43177 30175
rect 43211 30141 43223 30175
rect 43165 30135 43223 30141
rect 35584 30076 36492 30104
rect 38120 30104 38148 30132
rect 43180 30104 43208 30135
rect 43254 30104 43260 30116
rect 38120 30076 43260 30104
rect 35584 30064 35590 30076
rect 43254 30064 43260 30076
rect 43312 30064 43318 30116
rect 34330 30036 34336 30048
rect 32600 30008 34336 30036
rect 34330 29996 34336 30008
rect 34388 29996 34394 30048
rect 36722 29996 36728 30048
rect 36780 30036 36786 30048
rect 37090 30036 37096 30048
rect 36780 30008 37096 30036
rect 36780 29996 36786 30008
rect 37090 29996 37096 30008
rect 37148 29996 37154 30048
rect 37458 29996 37464 30048
rect 37516 29996 37522 30048
rect 37550 29996 37556 30048
rect 37608 30036 37614 30048
rect 41046 30036 41052 30048
rect 37608 30008 41052 30036
rect 37608 29996 37614 30008
rect 41046 29996 41052 30008
rect 41104 29996 41110 30048
rect 41138 29996 41144 30048
rect 41196 29996 41202 30048
rect 1104 29946 43884 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 43884 29946
rect 1104 29872 43884 29894
rect 9214 29792 9220 29844
rect 9272 29832 9278 29844
rect 11514 29832 11520 29844
rect 9272 29804 11520 29832
rect 9272 29792 9278 29804
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 11606 29792 11612 29844
rect 11664 29792 11670 29844
rect 17218 29792 17224 29844
rect 17276 29832 17282 29844
rect 17276 29804 18736 29832
rect 17276 29792 17282 29804
rect 8110 29764 8116 29776
rect 6840 29736 8116 29764
rect 6840 29637 6868 29736
rect 8110 29724 8116 29736
rect 8168 29724 8174 29776
rect 17865 29767 17923 29773
rect 17865 29733 17877 29767
rect 17911 29733 17923 29767
rect 18708 29764 18736 29804
rect 18782 29792 18788 29844
rect 18840 29832 18846 29844
rect 19242 29832 19248 29844
rect 18840 29804 19248 29832
rect 18840 29792 18846 29804
rect 19242 29792 19248 29804
rect 19300 29832 19306 29844
rect 22830 29832 22836 29844
rect 19300 29804 22836 29832
rect 19300 29792 19306 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 23566 29792 23572 29844
rect 23624 29792 23630 29844
rect 24302 29792 24308 29844
rect 24360 29832 24366 29844
rect 32122 29832 32128 29844
rect 24360 29804 32128 29832
rect 24360 29792 24366 29804
rect 32122 29792 32128 29804
rect 32180 29792 32186 29844
rect 32401 29835 32459 29841
rect 32401 29801 32413 29835
rect 32447 29832 32459 29835
rect 33226 29832 33232 29844
rect 32447 29804 33232 29832
rect 32447 29801 32459 29804
rect 32401 29795 32459 29801
rect 33226 29792 33232 29804
rect 33284 29792 33290 29844
rect 33318 29792 33324 29844
rect 33376 29792 33382 29844
rect 33597 29835 33655 29841
rect 33597 29801 33609 29835
rect 33643 29832 33655 29835
rect 33962 29832 33968 29844
rect 33643 29804 33968 29832
rect 33643 29801 33655 29804
rect 33597 29795 33655 29801
rect 33962 29792 33968 29804
rect 34020 29792 34026 29844
rect 34514 29792 34520 29844
rect 34572 29832 34578 29844
rect 35526 29832 35532 29844
rect 34572 29804 35532 29832
rect 34572 29792 34578 29804
rect 35526 29792 35532 29804
rect 35584 29792 35590 29844
rect 36170 29792 36176 29844
rect 36228 29832 36234 29844
rect 36449 29835 36507 29841
rect 36449 29832 36461 29835
rect 36228 29804 36461 29832
rect 36228 29792 36234 29804
rect 36449 29801 36461 29804
rect 36495 29832 36507 29835
rect 36630 29832 36636 29844
rect 36495 29804 36636 29832
rect 36495 29801 36507 29804
rect 36449 29795 36507 29801
rect 36630 29792 36636 29804
rect 36688 29792 36694 29844
rect 41690 29832 41696 29844
rect 37844 29804 41696 29832
rect 25682 29764 25688 29776
rect 18708 29736 22876 29764
rect 17865 29727 17923 29733
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 16853 29699 16911 29705
rect 7156 29668 7972 29696
rect 7156 29656 7162 29668
rect 6825 29631 6883 29637
rect 6825 29597 6837 29631
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29628 6975 29631
rect 6963 29600 7144 29628
rect 6963 29597 6975 29600
rect 6917 29591 6975 29597
rect 7116 29572 7144 29600
rect 7190 29588 7196 29640
rect 7248 29588 7254 29640
rect 7944 29637 7972 29668
rect 16853 29665 16865 29699
rect 16899 29696 16911 29699
rect 17405 29699 17463 29705
rect 17405 29696 17417 29699
rect 16899 29668 17417 29696
rect 16899 29665 16911 29668
rect 16853 29659 16911 29665
rect 17405 29665 17417 29668
rect 17451 29665 17463 29699
rect 17880 29696 17908 29727
rect 18046 29696 18052 29708
rect 17880 29668 18052 29696
rect 17405 29659 17463 29665
rect 18046 29656 18052 29668
rect 18104 29656 18110 29708
rect 18230 29656 18236 29708
rect 18288 29696 18294 29708
rect 18288 29668 18828 29696
rect 18288 29656 18294 29668
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29597 7987 29631
rect 7929 29591 7987 29597
rect 8021 29631 8079 29637
rect 8021 29597 8033 29631
rect 8067 29628 8079 29631
rect 9306 29628 9312 29640
rect 8067 29600 9312 29628
rect 8067 29597 8079 29600
rect 8021 29591 8079 29597
rect 7009 29563 7067 29569
rect 7009 29529 7021 29563
rect 7055 29529 7067 29563
rect 7009 29523 7067 29529
rect 6638 29452 6644 29504
rect 6696 29452 6702 29504
rect 7024 29492 7052 29523
rect 7098 29520 7104 29572
rect 7156 29520 7162 29572
rect 7374 29520 7380 29572
rect 7432 29560 7438 29572
rect 7834 29560 7840 29572
rect 7432 29532 7840 29560
rect 7432 29520 7438 29532
rect 7834 29520 7840 29532
rect 7892 29560 7898 29572
rect 8036 29560 8064 29591
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 10229 29631 10287 29637
rect 10229 29597 10241 29631
rect 10275 29628 10287 29631
rect 11698 29628 11704 29640
rect 10275 29600 11704 29628
rect 10275 29597 10287 29600
rect 10229 29591 10287 29597
rect 11698 29588 11704 29600
rect 11756 29588 11762 29640
rect 12342 29588 12348 29640
rect 12400 29628 12406 29640
rect 12621 29631 12679 29637
rect 12621 29628 12633 29631
rect 12400 29600 12633 29628
rect 12400 29588 12406 29600
rect 12621 29597 12633 29600
rect 12667 29597 12679 29631
rect 12621 29591 12679 29597
rect 12802 29588 12808 29640
rect 12860 29588 12866 29640
rect 17586 29588 17592 29640
rect 17644 29588 17650 29640
rect 17681 29631 17739 29637
rect 17681 29597 17693 29631
rect 17727 29628 17739 29631
rect 17770 29628 17776 29640
rect 17727 29600 17776 29628
rect 17727 29597 17739 29600
rect 17681 29591 17739 29597
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 18800 29637 18828 29668
rect 18966 29656 18972 29708
rect 19024 29696 19030 29708
rect 19429 29699 19487 29705
rect 19429 29696 19441 29699
rect 19024 29668 19441 29696
rect 19024 29656 19030 29668
rect 19429 29665 19441 29668
rect 19475 29665 19487 29699
rect 20254 29696 20260 29708
rect 19429 29659 19487 29665
rect 19720 29668 20260 29696
rect 19720 29637 19748 29668
rect 20254 29656 20260 29668
rect 20312 29656 20318 29708
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18693 29631 18751 29637
rect 18003 29600 18460 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 7892 29532 8064 29560
rect 10496 29563 10554 29569
rect 7892 29520 7898 29532
rect 10496 29529 10508 29563
rect 10542 29560 10554 29563
rect 10686 29560 10692 29572
rect 10542 29532 10692 29560
rect 10542 29529 10554 29532
rect 10496 29523 10554 29529
rect 10686 29520 10692 29532
rect 10744 29520 10750 29572
rect 7745 29495 7803 29501
rect 7745 29492 7757 29495
rect 7024 29464 7757 29492
rect 7745 29461 7757 29464
rect 7791 29492 7803 29495
rect 8386 29492 8392 29504
rect 7791 29464 8392 29492
rect 7791 29461 7803 29464
rect 7745 29455 7803 29461
rect 8386 29452 8392 29464
rect 8444 29452 8450 29504
rect 12713 29495 12771 29501
rect 12713 29461 12725 29495
rect 12759 29492 12771 29495
rect 13354 29492 13360 29504
rect 12759 29464 13360 29492
rect 12759 29461 12771 29464
rect 12713 29455 12771 29461
rect 13354 29452 13360 29464
rect 13412 29452 13418 29504
rect 16206 29452 16212 29504
rect 16264 29452 16270 29504
rect 16574 29452 16580 29504
rect 16632 29452 16638 29504
rect 16669 29495 16727 29501
rect 16669 29461 16681 29495
rect 16715 29492 16727 29495
rect 16850 29492 16856 29504
rect 16715 29464 16856 29492
rect 16715 29461 16727 29464
rect 16669 29455 16727 29461
rect 16850 29452 16856 29464
rect 16908 29452 16914 29504
rect 18230 29452 18236 29504
rect 18288 29492 18294 29504
rect 18432 29501 18460 29600
rect 18693 29597 18705 29631
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 18785 29631 18843 29637
rect 18785 29597 18797 29631
rect 18831 29597 18843 29631
rect 18785 29591 18843 29597
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 18708 29560 18736 29591
rect 19794 29588 19800 29640
rect 19852 29588 19858 29640
rect 19886 29588 19892 29640
rect 19944 29588 19950 29640
rect 20073 29631 20131 29637
rect 20073 29597 20085 29631
rect 20119 29628 20131 29631
rect 20533 29631 20591 29637
rect 20533 29628 20545 29631
rect 20119 29600 20545 29628
rect 20119 29597 20131 29600
rect 20073 29591 20131 29597
rect 20533 29597 20545 29600
rect 20579 29597 20591 29631
rect 20533 29591 20591 29597
rect 20717 29631 20775 29637
rect 20717 29597 20729 29631
rect 20763 29628 20775 29631
rect 20806 29628 20812 29640
rect 20763 29600 20812 29628
rect 20763 29597 20775 29600
rect 20717 29591 20775 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 22848 29628 22876 29736
rect 22940 29736 25688 29764
rect 22940 29708 22968 29736
rect 25682 29724 25688 29736
rect 25740 29724 25746 29776
rect 30006 29764 30012 29776
rect 25792 29736 30012 29764
rect 22922 29656 22928 29708
rect 22980 29656 22986 29708
rect 23109 29699 23167 29705
rect 23109 29665 23121 29699
rect 23155 29696 23167 29699
rect 23198 29696 23204 29708
rect 23155 29668 23204 29696
rect 23155 29665 23167 29668
rect 23109 29659 23167 29665
rect 23198 29656 23204 29668
rect 23256 29656 23262 29708
rect 25792 29696 25820 29736
rect 30006 29724 30012 29736
rect 30064 29724 30070 29776
rect 23308 29668 25820 29696
rect 23308 29628 23336 29668
rect 27246 29656 27252 29708
rect 27304 29696 27310 29708
rect 27525 29699 27583 29705
rect 27525 29696 27537 29699
rect 27304 29668 27537 29696
rect 27304 29656 27310 29668
rect 27525 29665 27537 29668
rect 27571 29665 27583 29699
rect 27525 29659 27583 29665
rect 30098 29656 30104 29708
rect 30156 29656 30162 29708
rect 30374 29656 30380 29708
rect 30432 29656 30438 29708
rect 30561 29699 30619 29705
rect 30561 29665 30573 29699
rect 30607 29696 30619 29699
rect 31294 29696 31300 29708
rect 30607 29668 31300 29696
rect 30607 29665 30619 29668
rect 30561 29659 30619 29665
rect 31294 29656 31300 29668
rect 31352 29656 31358 29708
rect 31570 29656 31576 29708
rect 31628 29656 31634 29708
rect 22848 29600 23336 29628
rect 25314 29588 25320 29640
rect 25372 29628 25378 29640
rect 26605 29631 26663 29637
rect 26605 29628 26617 29631
rect 25372 29600 26617 29628
rect 25372 29588 25378 29600
rect 26605 29597 26617 29600
rect 26651 29597 26663 29631
rect 26605 29591 26663 29597
rect 26970 29588 26976 29640
rect 27028 29588 27034 29640
rect 27982 29588 27988 29640
rect 28040 29588 28046 29640
rect 28074 29588 28080 29640
rect 28132 29628 28138 29640
rect 28629 29631 28687 29637
rect 28629 29628 28641 29631
rect 28132 29600 28641 29628
rect 28132 29588 28138 29600
rect 28629 29597 28641 29600
rect 28675 29597 28687 29631
rect 28629 29591 28687 29597
rect 30653 29631 30711 29637
rect 30653 29597 30665 29631
rect 30699 29628 30711 29631
rect 31386 29628 31392 29640
rect 30699 29600 31392 29628
rect 30699 29597 30711 29600
rect 30653 29591 30711 29597
rect 31386 29588 31392 29600
rect 31444 29588 31450 29640
rect 31481 29631 31539 29637
rect 31481 29597 31493 29631
rect 31527 29597 31539 29631
rect 31588 29628 31616 29656
rect 31665 29631 31723 29637
rect 31665 29628 31677 29631
rect 31588 29600 31677 29628
rect 31481 29591 31539 29597
rect 31665 29597 31677 29600
rect 31711 29597 31723 29631
rect 31665 29591 31723 29597
rect 19334 29560 19340 29572
rect 18708 29532 19340 29560
rect 19334 29520 19340 29532
rect 19392 29520 19398 29572
rect 19587 29563 19645 29569
rect 19587 29529 19599 29563
rect 19633 29560 19645 29563
rect 22370 29560 22376 29572
rect 19633 29532 22376 29560
rect 19633 29529 19645 29532
rect 19587 29523 19645 29529
rect 22370 29520 22376 29532
rect 22428 29520 22434 29572
rect 26421 29563 26479 29569
rect 26421 29529 26433 29563
rect 26467 29560 26479 29563
rect 26510 29560 26516 29572
rect 26467 29532 26516 29560
rect 26467 29529 26479 29532
rect 26421 29523 26479 29529
rect 26510 29520 26516 29532
rect 26568 29520 26574 29572
rect 27522 29520 27528 29572
rect 27580 29560 27586 29572
rect 27617 29563 27675 29569
rect 27617 29560 27629 29563
rect 27580 29532 27629 29560
rect 27580 29520 27586 29532
rect 27617 29529 27629 29532
rect 27663 29529 27675 29563
rect 31110 29560 31116 29572
rect 27617 29523 27675 29529
rect 28000 29532 31116 29560
rect 18417 29495 18475 29501
rect 18417 29492 18429 29495
rect 18288 29464 18429 29492
rect 18288 29452 18294 29464
rect 18417 29461 18429 29464
rect 18463 29461 18475 29495
rect 18417 29455 18475 29461
rect 19426 29452 19432 29504
rect 19484 29492 19490 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 19484 29464 20637 29492
rect 19484 29452 19490 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 20625 29455 20683 29461
rect 23198 29452 23204 29504
rect 23256 29492 23262 29504
rect 28000 29492 28028 29532
rect 31110 29520 31116 29532
rect 31168 29520 31174 29572
rect 31202 29520 31208 29572
rect 31260 29560 31266 29572
rect 31496 29560 31524 29591
rect 31846 29588 31852 29640
rect 31904 29588 31910 29640
rect 32122 29588 32128 29640
rect 32180 29628 32186 29640
rect 32309 29631 32367 29637
rect 32309 29628 32321 29631
rect 32180 29600 32321 29628
rect 32180 29588 32186 29600
rect 32309 29597 32321 29600
rect 32355 29597 32367 29631
rect 32309 29591 32367 29597
rect 32950 29588 32956 29640
rect 33008 29588 33014 29640
rect 33134 29637 33140 29640
rect 33101 29631 33140 29637
rect 33101 29597 33113 29631
rect 33101 29591 33140 29597
rect 33134 29588 33140 29591
rect 33192 29588 33198 29640
rect 33336 29637 33364 29792
rect 35802 29696 35808 29708
rect 34900 29668 35808 29696
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29597 33379 29631
rect 33321 29591 33379 29597
rect 33410 29588 33416 29640
rect 33468 29637 33474 29640
rect 33468 29631 33495 29637
rect 33483 29597 33495 29631
rect 34514 29628 34520 29640
rect 33468 29591 33495 29597
rect 33612 29600 34520 29628
rect 33468 29588 33474 29591
rect 31260 29532 31524 29560
rect 31573 29563 31631 29569
rect 31260 29520 31266 29532
rect 31573 29529 31585 29563
rect 31619 29560 31631 29563
rect 31754 29560 31760 29572
rect 31619 29532 31760 29560
rect 31619 29529 31631 29532
rect 31573 29523 31631 29529
rect 31754 29520 31760 29532
rect 31812 29520 31818 29572
rect 33229 29563 33287 29569
rect 33229 29529 33241 29563
rect 33275 29560 33287 29563
rect 33612 29560 33640 29600
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34900 29637 34928 29668
rect 35802 29656 35808 29668
rect 35860 29656 35866 29708
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 34974 29588 34980 29640
rect 35032 29588 35038 29640
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 33275 29532 33640 29560
rect 33275 29529 33287 29532
rect 33229 29523 33287 29529
rect 34146 29520 34152 29572
rect 34204 29560 34210 29572
rect 35176 29560 35204 29591
rect 35986 29588 35992 29640
rect 36044 29628 36050 29640
rect 36044 29600 37044 29628
rect 36044 29588 36050 29600
rect 34204 29532 35204 29560
rect 35621 29563 35679 29569
rect 34204 29520 34210 29532
rect 35621 29529 35633 29563
rect 35667 29560 35679 29563
rect 36722 29560 36728 29572
rect 35667 29532 36728 29560
rect 35667 29529 35679 29532
rect 35621 29523 35679 29529
rect 36722 29520 36728 29532
rect 36780 29520 36786 29572
rect 23256 29464 28028 29492
rect 23256 29452 23262 29464
rect 28718 29452 28724 29504
rect 28776 29452 28782 29504
rect 30466 29452 30472 29504
rect 30524 29492 30530 29504
rect 31297 29495 31355 29501
rect 31297 29492 31309 29495
rect 30524 29464 31309 29492
rect 30524 29452 30530 29464
rect 31297 29461 31309 29464
rect 31343 29461 31355 29495
rect 37016 29492 37044 29600
rect 37090 29588 37096 29640
rect 37148 29628 37154 29640
rect 37844 29637 37872 29804
rect 41690 29792 41696 29804
rect 41748 29832 41754 29844
rect 41748 29804 42012 29832
rect 41748 29792 41754 29804
rect 41984 29705 42012 29804
rect 41969 29699 42027 29705
rect 41969 29665 41981 29699
rect 42015 29665 42027 29699
rect 41969 29659 42027 29665
rect 37829 29631 37887 29637
rect 37829 29628 37841 29631
rect 37148 29600 37841 29628
rect 37148 29588 37154 29600
rect 37829 29597 37841 29600
rect 37875 29597 37887 29631
rect 37829 29591 37887 29597
rect 41138 29588 41144 29640
rect 41196 29628 41202 29640
rect 41702 29631 41760 29637
rect 41702 29628 41714 29631
rect 41196 29600 41714 29628
rect 41196 29588 41202 29600
rect 41702 29597 41714 29600
rect 41748 29597 41760 29631
rect 41702 29591 41760 29597
rect 42889 29631 42947 29637
rect 42889 29597 42901 29631
rect 42935 29597 42947 29631
rect 42889 29591 42947 29597
rect 37458 29520 37464 29572
rect 37516 29560 37522 29572
rect 37562 29563 37620 29569
rect 37562 29560 37574 29563
rect 37516 29532 37574 29560
rect 37516 29520 37522 29532
rect 37562 29529 37574 29532
rect 37608 29529 37620 29563
rect 37562 29523 37620 29529
rect 37918 29520 37924 29572
rect 37976 29560 37982 29572
rect 42904 29560 42932 29591
rect 37976 29532 42932 29560
rect 37976 29520 37982 29532
rect 43162 29520 43168 29572
rect 43220 29520 43226 29572
rect 39390 29492 39396 29504
rect 37016 29464 39396 29492
rect 31297 29455 31355 29461
rect 39390 29452 39396 29464
rect 39448 29452 39454 29504
rect 40034 29452 40040 29504
rect 40092 29492 40098 29504
rect 40589 29495 40647 29501
rect 40589 29492 40601 29495
rect 40092 29464 40601 29492
rect 40092 29452 40098 29464
rect 40589 29461 40601 29464
rect 40635 29492 40647 29495
rect 41046 29492 41052 29504
rect 40635 29464 41052 29492
rect 40635 29461 40647 29464
rect 40589 29455 40647 29461
rect 41046 29452 41052 29464
rect 41104 29452 41110 29504
rect 1104 29402 43884 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 43884 29402
rect 1104 29328 43884 29350
rect 8294 29248 8300 29300
rect 8352 29288 8358 29300
rect 9033 29291 9091 29297
rect 9033 29288 9045 29291
rect 8352 29260 9045 29288
rect 8352 29248 8358 29260
rect 9033 29257 9045 29260
rect 9079 29288 9091 29291
rect 9214 29288 9220 29300
rect 9079 29260 9220 29288
rect 9079 29257 9091 29260
rect 9033 29251 9091 29257
rect 9214 29248 9220 29260
rect 9272 29248 9278 29300
rect 16850 29248 16856 29300
rect 16908 29248 16914 29300
rect 18046 29248 18052 29300
rect 18104 29248 18110 29300
rect 19334 29288 19340 29300
rect 18156 29260 19340 29288
rect 9122 29220 9128 29232
rect 7668 29192 9128 29220
rect 6914 29112 6920 29164
rect 6972 29152 6978 29164
rect 7668 29161 7696 29192
rect 9122 29180 9128 29192
rect 9180 29180 9186 29232
rect 17218 29180 17224 29232
rect 17276 29180 17282 29232
rect 18156 29220 18184 29260
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 25685 29291 25743 29297
rect 25685 29257 25697 29291
rect 25731 29288 25743 29291
rect 26142 29288 26148 29300
rect 25731 29260 26148 29288
rect 25731 29257 25743 29260
rect 25685 29251 25743 29257
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 27709 29291 27767 29297
rect 27709 29257 27721 29291
rect 27755 29288 27767 29291
rect 28074 29288 28080 29300
rect 27755 29260 28080 29288
rect 27755 29257 27767 29260
rect 27709 29251 27767 29257
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 28445 29291 28503 29297
rect 28445 29257 28457 29291
rect 28491 29288 28503 29291
rect 28626 29288 28632 29300
rect 28491 29260 28632 29288
rect 28491 29257 28503 29260
rect 28445 29251 28503 29257
rect 28626 29248 28632 29260
rect 28684 29248 28690 29300
rect 31110 29288 31116 29300
rect 30024 29260 31116 29288
rect 22922 29220 22928 29232
rect 17328 29192 18184 29220
rect 18800 29192 22928 29220
rect 7926 29161 7932 29164
rect 7653 29155 7711 29161
rect 7653 29152 7665 29155
rect 6972 29124 7665 29152
rect 6972 29112 6978 29124
rect 7653 29121 7665 29124
rect 7699 29121 7711 29155
rect 7653 29115 7711 29121
rect 7920 29115 7932 29161
rect 7926 29112 7932 29115
rect 7984 29112 7990 29164
rect 8202 29112 8208 29164
rect 8260 29152 8266 29164
rect 8260 29124 8800 29152
rect 8260 29112 8266 29124
rect 8772 29084 8800 29124
rect 11698 29112 11704 29164
rect 11756 29152 11762 29164
rect 13630 29161 13636 29164
rect 13357 29155 13415 29161
rect 13357 29152 13369 29155
rect 11756 29124 13369 29152
rect 11756 29112 11762 29124
rect 13357 29121 13369 29124
rect 13403 29121 13415 29155
rect 13357 29115 13415 29121
rect 13624 29115 13636 29161
rect 13630 29112 13636 29115
rect 13688 29112 13694 29164
rect 15930 29112 15936 29164
rect 15988 29152 15994 29164
rect 17328 29152 17356 29192
rect 17862 29152 17868 29164
rect 15988 29124 17356 29152
rect 17420 29124 17868 29152
rect 15988 29112 15994 29124
rect 17420 29096 17448 29124
rect 17862 29112 17868 29124
rect 17920 29112 17926 29164
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29152 18291 29155
rect 18414 29152 18420 29164
rect 18279 29124 18420 29152
rect 18279 29121 18291 29124
rect 18233 29115 18291 29121
rect 18414 29112 18420 29124
rect 18472 29112 18478 29164
rect 18506 29112 18512 29164
rect 18564 29112 18570 29164
rect 13170 29084 13176 29096
rect 8772 29056 13176 29084
rect 13170 29044 13176 29056
rect 13228 29044 13234 29096
rect 17310 29044 17316 29096
rect 17368 29044 17374 29096
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 17586 29044 17592 29096
rect 17644 29084 17650 29096
rect 18325 29087 18383 29093
rect 18325 29084 18337 29087
rect 17644 29056 18337 29084
rect 17644 29044 17650 29056
rect 18325 29053 18337 29056
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 14458 28976 14464 29028
rect 14516 29016 14522 29028
rect 14737 29019 14795 29025
rect 14737 29016 14749 29019
rect 14516 28988 14749 29016
rect 14516 28976 14522 28988
rect 14737 28985 14749 28988
rect 14783 29016 14795 29019
rect 17604 29016 17632 29044
rect 14783 28988 17632 29016
rect 14783 28985 14795 28988
rect 14737 28979 14795 28985
rect 17862 28976 17868 29028
rect 17920 29016 17926 29028
rect 18800 29016 18828 29192
rect 22922 29180 22928 29192
rect 22980 29180 22986 29232
rect 27890 29220 27896 29232
rect 27632 29192 27896 29220
rect 19426 29112 19432 29164
rect 19484 29112 19490 29164
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29152 19671 29155
rect 19978 29152 19984 29164
rect 19659 29124 19984 29152
rect 19659 29121 19671 29124
rect 19613 29115 19671 29121
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 25317 29155 25375 29161
rect 25317 29121 25329 29155
rect 25363 29152 25375 29155
rect 26418 29152 26424 29164
rect 25363 29124 26424 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 27632 29161 27660 29192
rect 27890 29180 27896 29192
rect 27948 29180 27954 29232
rect 28350 29180 28356 29232
rect 28408 29180 28414 29232
rect 28718 29180 28724 29232
rect 28776 29220 28782 29232
rect 29917 29223 29975 29229
rect 29917 29220 29929 29223
rect 28776 29192 29929 29220
rect 28776 29180 28782 29192
rect 29917 29189 29929 29192
rect 29963 29189 29975 29223
rect 29917 29183 29975 29189
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29121 27675 29155
rect 27617 29115 27675 29121
rect 27801 29155 27859 29161
rect 27801 29121 27813 29155
rect 27847 29121 27859 29155
rect 27908 29152 27936 29180
rect 28534 29152 28540 29164
rect 27908 29124 28540 29152
rect 27801 29115 27859 29121
rect 19150 29044 19156 29096
rect 19208 29084 19214 29096
rect 19245 29087 19303 29093
rect 19245 29084 19257 29087
rect 19208 29056 19257 29084
rect 19208 29044 19214 29056
rect 19245 29053 19257 29056
rect 19291 29053 19303 29087
rect 25406 29084 25412 29096
rect 19245 29047 19303 29053
rect 19352 29056 25412 29084
rect 17920 28988 18828 29016
rect 17920 28976 17926 28988
rect 19058 28976 19064 29028
rect 19116 29016 19122 29028
rect 19352 29016 19380 29056
rect 25406 29044 25412 29056
rect 25464 29084 25470 29096
rect 26694 29084 26700 29096
rect 25464 29056 26700 29084
rect 25464 29044 25470 29056
rect 26694 29044 26700 29056
rect 26752 29044 26758 29096
rect 27816 29084 27844 29115
rect 28534 29112 28540 29124
rect 28592 29112 28598 29164
rect 28629 29155 28687 29161
rect 28629 29121 28641 29155
rect 28675 29152 28687 29155
rect 29733 29155 29791 29161
rect 29733 29152 29745 29155
rect 28675 29124 29745 29152
rect 28675 29121 28687 29124
rect 28629 29115 28687 29121
rect 29733 29121 29745 29124
rect 29779 29152 29791 29155
rect 29822 29152 29828 29164
rect 29779 29124 29828 29152
rect 29779 29121 29791 29124
rect 29733 29115 29791 29121
rect 29822 29112 29828 29124
rect 29880 29112 29886 29164
rect 28442 29084 28448 29096
rect 27816 29056 28448 29084
rect 28442 29044 28448 29056
rect 28500 29044 28506 29096
rect 28721 29087 28779 29093
rect 28721 29053 28733 29087
rect 28767 29084 28779 29087
rect 30024 29084 30052 29260
rect 31110 29248 31116 29260
rect 31168 29248 31174 29300
rect 32306 29248 32312 29300
rect 32364 29288 32370 29300
rect 32953 29291 33011 29297
rect 32953 29288 32965 29291
rect 32364 29260 32965 29288
rect 32364 29248 32370 29260
rect 32953 29257 32965 29260
rect 32999 29257 33011 29291
rect 32953 29251 33011 29257
rect 34514 29248 34520 29300
rect 34572 29288 34578 29300
rect 34572 29260 34652 29288
rect 34572 29248 34578 29260
rect 30101 29223 30159 29229
rect 30101 29189 30113 29223
rect 30147 29220 30159 29223
rect 32398 29220 32404 29232
rect 30147 29192 32404 29220
rect 30147 29189 30159 29192
rect 30101 29183 30159 29189
rect 32398 29180 32404 29192
rect 32456 29180 32462 29232
rect 32861 29223 32919 29229
rect 32861 29220 32873 29223
rect 32600 29192 32873 29220
rect 30742 29112 30748 29164
rect 30800 29152 30806 29164
rect 31021 29155 31079 29161
rect 31021 29152 31033 29155
rect 30800 29124 31033 29152
rect 30800 29112 30806 29124
rect 31021 29121 31033 29124
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 31110 29112 31116 29164
rect 31168 29152 31174 29164
rect 31478 29152 31484 29164
rect 31168 29124 31484 29152
rect 31168 29112 31174 29124
rect 31478 29112 31484 29124
rect 31536 29152 31542 29164
rect 32600 29152 32628 29192
rect 32861 29189 32873 29192
rect 32907 29220 32919 29223
rect 33226 29220 33232 29232
rect 32907 29192 33232 29220
rect 32907 29189 32919 29192
rect 32861 29183 32919 29189
rect 33226 29180 33232 29192
rect 33284 29180 33290 29232
rect 34624 29229 34652 29260
rect 36722 29248 36728 29300
rect 36780 29288 36786 29300
rect 37366 29288 37372 29300
rect 36780 29260 37372 29288
rect 36780 29248 36786 29260
rect 37366 29248 37372 29260
rect 37424 29248 37430 29300
rect 38470 29248 38476 29300
rect 38528 29288 38534 29300
rect 39206 29288 39212 29300
rect 38528 29260 39212 29288
rect 38528 29248 38534 29260
rect 39206 29248 39212 29260
rect 39264 29248 39270 29300
rect 39577 29291 39635 29297
rect 39577 29257 39589 29291
rect 39623 29288 39635 29291
rect 39623 29260 40908 29288
rect 39623 29257 39635 29260
rect 39577 29251 39635 29257
rect 34609 29223 34667 29229
rect 34609 29189 34621 29223
rect 34655 29189 34667 29223
rect 34609 29183 34667 29189
rect 35618 29180 35624 29232
rect 35676 29180 35682 29232
rect 38197 29223 38255 29229
rect 38197 29189 38209 29223
rect 38243 29220 38255 29223
rect 38243 29192 39620 29220
rect 38243 29189 38255 29192
rect 38197 29183 38255 29189
rect 31536 29124 32628 29152
rect 31536 29112 31542 29124
rect 33134 29112 33140 29164
rect 33192 29112 33198 29164
rect 34422 29112 34428 29164
rect 34480 29112 34486 29164
rect 34701 29155 34759 29161
rect 34701 29121 34713 29155
rect 34747 29121 34759 29155
rect 34701 29115 34759 29121
rect 28767 29056 30052 29084
rect 30837 29087 30895 29093
rect 28767 29053 28779 29056
rect 28721 29047 28779 29053
rect 30837 29053 30849 29087
rect 30883 29084 30895 29087
rect 31294 29084 31300 29096
rect 30883 29056 31300 29084
rect 30883 29053 30895 29056
rect 30837 29047 30895 29053
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 33321 29087 33379 29093
rect 33321 29053 33333 29087
rect 33367 29084 33379 29087
rect 33962 29084 33968 29096
rect 33367 29056 33968 29084
rect 33367 29053 33379 29056
rect 33321 29047 33379 29053
rect 33962 29044 33968 29056
rect 34020 29044 34026 29096
rect 34716 29084 34744 29115
rect 34790 29112 34796 29164
rect 34848 29112 34854 29164
rect 35986 29112 35992 29164
rect 36044 29152 36050 29164
rect 36357 29155 36415 29161
rect 36357 29152 36369 29155
rect 36044 29124 36369 29152
rect 36044 29112 36050 29124
rect 36357 29121 36369 29124
rect 36403 29121 36415 29155
rect 36357 29115 36415 29121
rect 37274 29112 37280 29164
rect 37332 29152 37338 29164
rect 37461 29155 37519 29161
rect 37461 29152 37473 29155
rect 37332 29124 37473 29152
rect 37332 29112 37338 29124
rect 37461 29121 37473 29124
rect 37507 29152 37519 29155
rect 37550 29152 37556 29164
rect 37507 29124 37556 29152
rect 37507 29121 37519 29124
rect 37461 29115 37519 29121
rect 37550 29112 37556 29124
rect 37608 29112 37614 29164
rect 37642 29112 37648 29164
rect 37700 29161 37706 29164
rect 37700 29155 37749 29161
rect 37700 29121 37703 29155
rect 37737 29152 37749 29155
rect 37737 29124 38240 29152
rect 37737 29121 37749 29124
rect 37700 29115 37749 29121
rect 37700 29112 37706 29115
rect 38212 29096 38240 29124
rect 38286 29112 38292 29164
rect 38344 29152 38350 29164
rect 38654 29152 38660 29164
rect 38344 29124 38660 29152
rect 38344 29112 38350 29124
rect 38654 29112 38660 29124
rect 38712 29152 38718 29164
rect 39114 29161 39120 29164
rect 38933 29155 38991 29161
rect 38933 29152 38945 29155
rect 38712 29124 38945 29152
rect 38712 29112 38718 29124
rect 38933 29121 38945 29124
rect 38979 29121 38991 29155
rect 38933 29115 38991 29121
rect 39081 29155 39120 29161
rect 39081 29121 39093 29155
rect 39081 29115 39120 29121
rect 39114 29112 39120 29115
rect 39172 29112 39178 29164
rect 39206 29112 39212 29164
rect 39264 29112 39270 29164
rect 39301 29155 39359 29161
rect 39301 29121 39313 29155
rect 39347 29121 39359 29155
rect 39301 29115 39359 29121
rect 37829 29087 37887 29093
rect 34716 29056 35112 29084
rect 19116 28988 19380 29016
rect 19444 28988 19656 29016
rect 19116 28976 19122 28988
rect 13998 28908 14004 28960
rect 14056 28948 14062 28960
rect 14642 28948 14648 28960
rect 14056 28920 14648 28948
rect 14056 28908 14062 28920
rect 14642 28908 14648 28920
rect 14700 28908 14706 28960
rect 18509 28951 18567 28957
rect 18509 28917 18521 28951
rect 18555 28948 18567 28951
rect 19444 28948 19472 28988
rect 18555 28920 19472 28948
rect 19628 28948 19656 28988
rect 26050 28976 26056 29028
rect 26108 29016 26114 29028
rect 26108 28988 27384 29016
rect 26108 28976 26114 28988
rect 22554 28948 22560 28960
rect 19628 28920 22560 28948
rect 18555 28917 18567 28920
rect 18509 28911 18567 28917
rect 22554 28908 22560 28920
rect 22612 28908 22618 28960
rect 27356 28948 27384 28988
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 34716 29016 34744 29056
rect 27488 28988 34744 29016
rect 27488 28976 27494 28988
rect 34790 28976 34796 29028
rect 34848 29016 34854 29028
rect 34977 29019 35035 29025
rect 34977 29016 34989 29019
rect 34848 28988 34989 29016
rect 34848 28976 34854 28988
rect 34977 28985 34989 28988
rect 35023 28985 35035 29019
rect 35084 29016 35112 29056
rect 37829 29053 37841 29087
rect 37875 29084 37887 29087
rect 38102 29084 38108 29096
rect 37875 29056 38108 29084
rect 37875 29053 37887 29056
rect 37829 29047 37887 29053
rect 38102 29044 38108 29056
rect 38160 29044 38166 29096
rect 38194 29044 38200 29096
rect 38252 29044 38258 29096
rect 38746 29044 38752 29096
rect 38804 29084 38810 29096
rect 39316 29084 39344 29115
rect 39390 29112 39396 29164
rect 39448 29161 39454 29164
rect 39448 29152 39456 29161
rect 39448 29124 39493 29152
rect 39448 29115 39456 29124
rect 39448 29112 39454 29115
rect 38804 29056 39344 29084
rect 39592 29084 39620 29192
rect 39942 29180 39948 29232
rect 40000 29220 40006 29232
rect 40880 29229 40908 29260
rect 41046 29248 41052 29300
rect 41104 29248 41110 29300
rect 40405 29223 40463 29229
rect 40405 29220 40417 29223
rect 40000 29192 40417 29220
rect 40000 29180 40006 29192
rect 40405 29189 40417 29192
rect 40451 29189 40463 29223
rect 40405 29183 40463 29189
rect 40865 29223 40923 29229
rect 40865 29189 40877 29223
rect 40911 29189 40923 29223
rect 40865 29183 40923 29189
rect 40126 29112 40132 29164
rect 40184 29112 40190 29164
rect 40310 29112 40316 29164
rect 40368 29112 40374 29164
rect 41138 29112 41144 29164
rect 41196 29112 41202 29164
rect 40218 29084 40224 29096
rect 39592 29056 40224 29084
rect 38804 29044 38810 29056
rect 40218 29044 40224 29056
rect 40276 29044 40282 29096
rect 40328 29084 40356 29112
rect 40328 29056 40908 29084
rect 40034 29016 40040 29028
rect 35084 28988 40040 29016
rect 34977 28979 35035 28985
rect 40034 28976 40040 28988
rect 40092 28976 40098 29028
rect 40880 29025 40908 29056
rect 40865 29019 40923 29025
rect 40865 28985 40877 29019
rect 40911 28985 40923 29019
rect 40865 28979 40923 28985
rect 28537 28951 28595 28957
rect 28537 28948 28549 28951
rect 27356 28920 28549 28948
rect 28537 28917 28549 28920
rect 28583 28917 28595 28951
rect 28537 28911 28595 28917
rect 32030 28908 32036 28960
rect 32088 28948 32094 28960
rect 36906 28948 36912 28960
rect 32088 28920 36912 28948
rect 32088 28908 32094 28920
rect 36906 28908 36912 28920
rect 36964 28908 36970 28960
rect 37366 28908 37372 28960
rect 37424 28948 37430 28960
rect 37599 28951 37657 28957
rect 37599 28948 37611 28951
rect 37424 28920 37611 28948
rect 37424 28908 37430 28920
rect 37599 28917 37611 28920
rect 37645 28948 37657 28951
rect 39298 28948 39304 28960
rect 37645 28920 39304 28948
rect 37645 28917 37657 28920
rect 37599 28911 37657 28917
rect 39298 28908 39304 28920
rect 39356 28908 39362 28960
rect 1104 28858 43884 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 43884 28858
rect 1104 28784 43884 28806
rect 7926 28704 7932 28756
rect 7984 28744 7990 28756
rect 8021 28747 8079 28753
rect 8021 28744 8033 28747
rect 7984 28716 8033 28744
rect 7984 28704 7990 28716
rect 8021 28713 8033 28716
rect 8067 28713 8079 28747
rect 8021 28707 8079 28713
rect 8110 28704 8116 28756
rect 8168 28744 8174 28756
rect 11146 28744 11152 28756
rect 8168 28716 11152 28744
rect 8168 28704 8174 28716
rect 11146 28704 11152 28716
rect 11204 28744 11210 28756
rect 12342 28744 12348 28756
rect 11204 28716 12348 28744
rect 11204 28704 11210 28716
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 13630 28704 13636 28756
rect 13688 28744 13694 28756
rect 13725 28747 13783 28753
rect 13725 28744 13737 28747
rect 13688 28716 13737 28744
rect 13688 28704 13694 28716
rect 13725 28713 13737 28716
rect 13771 28713 13783 28747
rect 18506 28744 18512 28756
rect 13725 28707 13783 28713
rect 14568 28716 18512 28744
rect 6917 28679 6975 28685
rect 6917 28645 6929 28679
rect 6963 28676 6975 28679
rect 7098 28676 7104 28688
rect 6963 28648 7104 28676
rect 6963 28645 6975 28648
rect 6917 28639 6975 28645
rect 7098 28636 7104 28648
rect 7156 28676 7162 28688
rect 8202 28676 8208 28688
rect 7156 28648 8208 28676
rect 7156 28636 7162 28648
rect 8202 28636 8208 28648
rect 8260 28636 8266 28688
rect 14458 28608 14464 28620
rect 13464 28580 14464 28608
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28540 5595 28543
rect 5626 28540 5632 28552
rect 5583 28512 5632 28540
rect 5583 28509 5595 28512
rect 5537 28503 5595 28509
rect 5626 28500 5632 28512
rect 5684 28540 5690 28552
rect 6822 28540 6828 28552
rect 5684 28512 6828 28540
rect 5684 28500 5690 28512
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 8110 28500 8116 28552
rect 8168 28540 8174 28552
rect 8205 28543 8263 28549
rect 8205 28540 8217 28543
rect 8168 28512 8217 28540
rect 8168 28500 8174 28512
rect 8205 28509 8217 28512
rect 8251 28509 8263 28543
rect 8205 28503 8263 28509
rect 8294 28500 8300 28552
rect 8352 28500 8358 28552
rect 8570 28500 8576 28552
rect 8628 28500 8634 28552
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 9398 28549 9404 28552
rect 9392 28540 9404 28549
rect 9359 28512 9404 28540
rect 9392 28503 9404 28512
rect 9398 28500 9404 28503
rect 9456 28500 9462 28552
rect 12710 28500 12716 28552
rect 12768 28540 12774 28552
rect 13464 28549 13492 28580
rect 14458 28568 14464 28580
rect 14516 28568 14522 28620
rect 13173 28543 13231 28549
rect 13173 28540 13185 28543
rect 12768 28512 13185 28540
rect 12768 28500 12774 28512
rect 13173 28509 13185 28512
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13449 28543 13507 28549
rect 13449 28509 13461 28543
rect 13495 28509 13507 28543
rect 13449 28503 13507 28509
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13998 28540 14004 28552
rect 13587 28512 14004 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 14568 28549 14596 28716
rect 18506 28704 18512 28716
rect 18564 28704 18570 28756
rect 20898 28704 20904 28756
rect 20956 28704 20962 28756
rect 22830 28704 22836 28756
rect 22888 28704 22894 28756
rect 27154 28704 27160 28756
rect 27212 28744 27218 28756
rect 32490 28744 32496 28756
rect 27212 28716 32496 28744
rect 27212 28704 27218 28716
rect 32490 28704 32496 28716
rect 32548 28704 32554 28756
rect 32769 28747 32827 28753
rect 32769 28713 32781 28747
rect 32815 28744 32827 28747
rect 32950 28744 32956 28756
rect 32815 28716 32956 28744
rect 32815 28713 32827 28716
rect 32769 28707 32827 28713
rect 32950 28704 32956 28716
rect 33008 28704 33014 28756
rect 36906 28704 36912 28756
rect 36964 28744 36970 28756
rect 38102 28744 38108 28756
rect 36964 28716 38108 28744
rect 36964 28704 36970 28716
rect 38102 28704 38108 28716
rect 38160 28704 38166 28756
rect 39114 28704 39120 28756
rect 39172 28744 39178 28756
rect 42978 28744 42984 28756
rect 39172 28716 42984 28744
rect 39172 28704 39178 28716
rect 16574 28636 16580 28688
rect 16632 28676 16638 28688
rect 16853 28679 16911 28685
rect 16853 28676 16865 28679
rect 16632 28648 16865 28676
rect 16632 28636 16638 28648
rect 16853 28645 16865 28648
rect 16899 28676 16911 28679
rect 19518 28676 19524 28688
rect 16899 28648 19524 28676
rect 16899 28645 16911 28648
rect 16853 28639 16911 28645
rect 19518 28636 19524 28648
rect 19576 28636 19582 28688
rect 27614 28636 27620 28688
rect 27672 28676 27678 28688
rect 28077 28679 28135 28685
rect 28077 28676 28089 28679
rect 27672 28648 28089 28676
rect 27672 28636 27678 28648
rect 28077 28645 28089 28648
rect 28123 28645 28135 28679
rect 28077 28639 28135 28645
rect 28258 28636 28264 28688
rect 28316 28676 28322 28688
rect 28316 28648 28764 28676
rect 28316 28636 28322 28648
rect 18414 28568 18420 28620
rect 18472 28568 18478 28620
rect 24578 28608 24584 28620
rect 18524 28580 19458 28608
rect 22848 28580 24584 28608
rect 14553 28543 14611 28549
rect 14553 28540 14565 28543
rect 14384 28512 14565 28540
rect 5804 28475 5862 28481
rect 5804 28441 5816 28475
rect 5850 28472 5862 28475
rect 6638 28472 6644 28484
rect 5850 28444 6644 28472
rect 5850 28441 5862 28444
rect 5804 28435 5862 28441
rect 6638 28432 6644 28444
rect 6696 28432 6702 28484
rect 8386 28432 8392 28484
rect 8444 28472 8450 28484
rect 12434 28472 12440 28484
rect 8444 28444 12440 28472
rect 8444 28432 8450 28444
rect 12434 28432 12440 28444
rect 12492 28432 12498 28484
rect 13354 28432 13360 28484
rect 13412 28432 13418 28484
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14384 28472 14412 28512
rect 14553 28509 14565 28512
rect 14599 28509 14611 28543
rect 14553 28503 14611 28509
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 14734 28540 14740 28552
rect 14691 28512 14740 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 14734 28500 14740 28512
rect 14792 28500 14798 28552
rect 15194 28500 15200 28552
rect 15252 28540 15258 28552
rect 15473 28543 15531 28549
rect 15473 28540 15485 28543
rect 15252 28512 15485 28540
rect 15252 28500 15258 28512
rect 15473 28509 15485 28512
rect 15519 28540 15531 28543
rect 18138 28540 18144 28552
rect 15519 28512 18144 28540
rect 15519 28509 15531 28512
rect 15473 28503 15531 28509
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 13872 28444 14412 28472
rect 13872 28432 13878 28444
rect 14458 28432 14464 28484
rect 14516 28432 14522 28484
rect 15740 28475 15798 28481
rect 14752 28444 14964 28472
rect 10505 28407 10563 28413
rect 10505 28373 10517 28407
rect 10551 28404 10563 28407
rect 14752 28404 14780 28444
rect 10551 28376 14780 28404
rect 10551 28373 10563 28376
rect 10505 28367 10563 28373
rect 14826 28364 14832 28416
rect 14884 28364 14890 28416
rect 14936 28404 14964 28444
rect 15740 28441 15752 28475
rect 15786 28472 15798 28475
rect 16206 28472 16212 28484
rect 15786 28444 16212 28472
rect 15786 28441 15798 28444
rect 15740 28435 15798 28441
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 18524 28472 18552 28580
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28540 19947 28543
rect 21542 28540 21548 28552
rect 19935 28512 21548 28540
rect 19935 28509 19947 28512
rect 19889 28503 19947 28509
rect 21542 28500 21548 28512
rect 21600 28500 21606 28552
rect 22848 28549 22876 28580
rect 24578 28568 24584 28580
rect 24636 28568 24642 28620
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28540 22983 28543
rect 23014 28540 23020 28552
rect 22971 28512 23020 28540
rect 22971 28509 22983 28512
rect 22925 28503 22983 28509
rect 16316 28444 18552 28472
rect 19981 28475 20039 28481
rect 16316 28404 16344 28444
rect 19981 28441 19993 28475
rect 20027 28472 20039 28475
rect 20070 28472 20076 28484
rect 20027 28444 20076 28472
rect 20027 28441 20039 28444
rect 19981 28435 20039 28441
rect 20070 28432 20076 28444
rect 20128 28432 20134 28484
rect 20349 28475 20407 28481
rect 20349 28441 20361 28475
rect 20395 28472 20407 28475
rect 20438 28472 20444 28484
rect 20395 28444 20444 28472
rect 20395 28441 20407 28444
rect 20349 28435 20407 28441
rect 20438 28432 20444 28444
rect 20496 28432 20502 28484
rect 20806 28472 20812 28484
rect 20640 28444 20812 28472
rect 14936 28376 16344 28404
rect 17678 28364 17684 28416
rect 17736 28404 17742 28416
rect 17773 28407 17831 28413
rect 17773 28404 17785 28407
rect 17736 28376 17785 28404
rect 17736 28364 17742 28376
rect 17773 28373 17785 28376
rect 17819 28373 17831 28407
rect 17773 28367 17831 28373
rect 17954 28364 17960 28416
rect 18012 28404 18018 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 18012 28376 18153 28404
rect 18012 28364 18018 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 18141 28367 18199 28373
rect 18233 28407 18291 28413
rect 18233 28373 18245 28407
rect 18279 28404 18291 28407
rect 18506 28404 18512 28416
rect 18279 28376 18512 28404
rect 18279 28373 18291 28376
rect 18233 28367 18291 28373
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 19518 28364 19524 28416
rect 19576 28404 19582 28416
rect 19613 28407 19671 28413
rect 19613 28404 19625 28407
rect 19576 28376 19625 28404
rect 19576 28364 19582 28376
rect 19613 28373 19625 28376
rect 19659 28404 19671 28407
rect 20640 28404 20668 28444
rect 20806 28432 20812 28444
rect 20864 28432 20870 28484
rect 20898 28432 20904 28484
rect 20956 28472 20962 28484
rect 22848 28472 22876 28503
rect 23014 28500 23020 28512
rect 23072 28500 23078 28552
rect 23198 28500 23204 28552
rect 23256 28540 23262 28552
rect 24857 28543 24915 28549
rect 24857 28540 24869 28543
rect 23256 28512 24869 28540
rect 23256 28500 23262 28512
rect 24857 28509 24869 28512
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 26786 28500 26792 28552
rect 26844 28540 26850 28552
rect 26844 28512 27752 28540
rect 26844 28500 26850 28512
rect 20956 28444 22876 28472
rect 20956 28432 20962 28444
rect 23106 28432 23112 28484
rect 23164 28432 23170 28484
rect 24118 28432 24124 28484
rect 24176 28472 24182 28484
rect 25102 28475 25160 28481
rect 25102 28472 25114 28475
rect 24176 28444 25114 28472
rect 24176 28432 24182 28444
rect 25102 28441 25114 28444
rect 25148 28441 25160 28475
rect 25102 28435 25160 28441
rect 27154 28432 27160 28484
rect 27212 28432 27218 28484
rect 19659 28376 20668 28404
rect 20717 28407 20775 28413
rect 19659 28373 19671 28376
rect 19613 28367 19671 28373
rect 20717 28373 20729 28407
rect 20763 28404 20775 28407
rect 21082 28404 21088 28416
rect 20763 28376 21088 28404
rect 20763 28373 20775 28376
rect 20717 28367 20775 28373
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28404 22707 28407
rect 23014 28404 23020 28416
rect 22695 28376 23020 28404
rect 22695 28373 22707 28376
rect 22649 28367 22707 28373
rect 23014 28364 23020 28376
rect 23072 28364 23078 28416
rect 26237 28407 26295 28413
rect 26237 28373 26249 28407
rect 26283 28404 26295 28407
rect 26418 28404 26424 28416
rect 26283 28376 26424 28404
rect 26283 28373 26295 28376
rect 26237 28367 26295 28373
rect 26418 28364 26424 28376
rect 26476 28364 26482 28416
rect 27724 28404 27752 28512
rect 27982 28500 27988 28552
rect 28040 28500 28046 28552
rect 28736 28549 28764 28648
rect 30374 28636 30380 28688
rect 30432 28676 30438 28688
rect 30469 28679 30527 28685
rect 30469 28676 30481 28679
rect 30432 28648 30481 28676
rect 30432 28636 30438 28648
rect 30469 28645 30481 28648
rect 30515 28645 30527 28679
rect 39022 28676 39028 28688
rect 30469 28639 30527 28645
rect 31349 28648 39028 28676
rect 28902 28568 28908 28620
rect 28960 28608 28966 28620
rect 31349 28608 31377 28648
rect 39022 28636 39028 28648
rect 39080 28636 39086 28688
rect 28960 28580 31377 28608
rect 28960 28568 28966 28580
rect 32490 28568 32496 28620
rect 32548 28608 32554 28620
rect 33137 28611 33195 28617
rect 33137 28608 33149 28611
rect 32548 28580 33149 28608
rect 32548 28568 32554 28580
rect 33137 28577 33149 28580
rect 33183 28608 33195 28611
rect 34146 28608 34152 28620
rect 33183 28580 34152 28608
rect 33183 28577 33195 28580
rect 33137 28571 33195 28577
rect 34146 28568 34152 28580
rect 34204 28568 34210 28620
rect 37642 28608 37648 28620
rect 37200 28580 37648 28608
rect 28537 28543 28595 28549
rect 28537 28509 28549 28543
rect 28583 28509 28595 28543
rect 28537 28503 28595 28509
rect 28721 28543 28779 28549
rect 28721 28509 28733 28543
rect 28767 28509 28779 28543
rect 29454 28540 29460 28552
rect 28721 28503 28779 28509
rect 28828 28512 29460 28540
rect 28552 28472 28580 28503
rect 28828 28472 28856 28512
rect 29454 28500 29460 28512
rect 29512 28500 29518 28552
rect 29822 28500 29828 28552
rect 29880 28540 29886 28552
rect 30193 28543 30251 28549
rect 30193 28540 30205 28543
rect 29880 28512 30205 28540
rect 29880 28500 29886 28512
rect 30193 28509 30205 28512
rect 30239 28540 30251 28543
rect 30282 28540 30288 28552
rect 30239 28512 30288 28540
rect 30239 28509 30251 28512
rect 30193 28503 30251 28509
rect 30282 28500 30288 28512
rect 30340 28500 30346 28552
rect 30466 28500 30472 28552
rect 30524 28500 30530 28552
rect 30834 28500 30840 28552
rect 30892 28540 30898 28552
rect 31202 28540 31208 28552
rect 30892 28512 31208 28540
rect 30892 28500 30898 28512
rect 31202 28500 31208 28512
rect 31260 28540 31266 28552
rect 31297 28543 31355 28549
rect 31297 28540 31309 28543
rect 31260 28512 31309 28540
rect 31260 28500 31266 28512
rect 31297 28509 31309 28512
rect 31343 28509 31355 28543
rect 31297 28503 31355 28509
rect 31481 28543 31539 28549
rect 31481 28509 31493 28543
rect 31527 28540 31539 28543
rect 31570 28540 31576 28552
rect 31527 28512 31576 28540
rect 31527 28509 31539 28512
rect 31481 28503 31539 28509
rect 31570 28500 31576 28512
rect 31628 28500 31634 28552
rect 31665 28543 31723 28549
rect 31665 28509 31677 28543
rect 31711 28540 31723 28543
rect 32030 28540 32036 28552
rect 31711 28512 32036 28540
rect 31711 28509 31723 28512
rect 31665 28503 31723 28509
rect 32030 28500 32036 28512
rect 32088 28500 32094 28552
rect 32214 28500 32220 28552
rect 32272 28540 32278 28552
rect 32582 28540 32588 28552
rect 32272 28512 32588 28540
rect 32272 28500 32278 28512
rect 32582 28500 32588 28512
rect 32640 28540 32646 28552
rect 32953 28543 33011 28549
rect 32953 28540 32965 28543
rect 32640 28512 32965 28540
rect 32640 28500 32646 28512
rect 32953 28509 32965 28512
rect 32999 28509 33011 28543
rect 32953 28503 33011 28509
rect 33226 28500 33232 28552
rect 33284 28500 33290 28552
rect 34330 28500 34336 28552
rect 34388 28540 34394 28552
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34388 28512 34897 28540
rect 34388 28500 34394 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 34977 28543 35035 28549
rect 34977 28509 34989 28543
rect 35023 28540 35035 28543
rect 35066 28540 35072 28552
rect 35023 28512 35072 28540
rect 35023 28509 35035 28512
rect 34977 28503 35035 28509
rect 35066 28500 35072 28512
rect 35124 28500 35130 28552
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28509 35219 28543
rect 35161 28503 35219 28509
rect 31389 28475 31447 28481
rect 28552 28444 28856 28472
rect 28920 28444 31340 28472
rect 28920 28404 28948 28444
rect 27724 28376 28948 28404
rect 29546 28364 29552 28416
rect 29604 28404 29610 28416
rect 30285 28407 30343 28413
rect 30285 28404 30297 28407
rect 29604 28376 30297 28404
rect 29604 28364 29610 28376
rect 30285 28373 30297 28376
rect 30331 28373 30343 28407
rect 30285 28367 30343 28373
rect 31113 28407 31171 28413
rect 31113 28373 31125 28407
rect 31159 28404 31171 28407
rect 31202 28404 31208 28416
rect 31159 28376 31208 28404
rect 31159 28373 31171 28376
rect 31113 28367 31171 28373
rect 31202 28364 31208 28376
rect 31260 28364 31266 28416
rect 31312 28404 31340 28444
rect 31389 28441 31401 28475
rect 31435 28472 31447 28475
rect 31846 28472 31852 28484
rect 31435 28444 31852 28472
rect 31435 28441 31447 28444
rect 31389 28435 31447 28441
rect 31846 28432 31852 28444
rect 31904 28432 31910 28484
rect 32858 28432 32864 28484
rect 32916 28472 32922 28484
rect 33134 28472 33140 28484
rect 32916 28444 33140 28472
rect 32916 28432 32922 28444
rect 33134 28432 33140 28444
rect 33192 28432 33198 28484
rect 33244 28472 33272 28500
rect 34238 28472 34244 28484
rect 33244 28444 34244 28472
rect 34238 28432 34244 28444
rect 34296 28472 34302 28484
rect 34422 28472 34428 28484
rect 34296 28444 34428 28472
rect 34296 28432 34302 28444
rect 34422 28432 34428 28444
rect 34480 28472 34486 28484
rect 35176 28472 35204 28503
rect 35434 28500 35440 28552
rect 35492 28540 35498 28552
rect 35621 28543 35679 28549
rect 35621 28540 35633 28543
rect 35492 28512 35633 28540
rect 35492 28500 35498 28512
rect 35621 28509 35633 28512
rect 35667 28540 35679 28543
rect 36906 28540 36912 28552
rect 35667 28512 36912 28540
rect 35667 28509 35679 28512
rect 35621 28503 35679 28509
rect 36906 28500 36912 28512
rect 36964 28500 36970 28552
rect 37200 28549 37228 28580
rect 37642 28568 37648 28580
rect 37700 28568 37706 28620
rect 38212 28580 39068 28608
rect 37185 28543 37243 28549
rect 37185 28509 37197 28543
rect 37231 28509 37243 28543
rect 37185 28503 37243 28509
rect 37366 28500 37372 28552
rect 37424 28500 37430 28552
rect 37550 28500 37556 28552
rect 37608 28540 37614 28552
rect 38212 28540 38240 28580
rect 37608 28512 38240 28540
rect 37608 28500 37614 28512
rect 38838 28500 38844 28552
rect 38896 28500 38902 28552
rect 38934 28543 38992 28549
rect 38934 28509 38946 28543
rect 38980 28509 38992 28543
rect 38934 28503 38992 28509
rect 34480 28444 35204 28472
rect 34480 28432 34486 28444
rect 35250 28432 35256 28484
rect 35308 28472 35314 28484
rect 38948 28472 38976 28503
rect 39040 28484 39068 28580
rect 39224 28549 39252 28716
rect 42978 28704 42984 28716
rect 43036 28744 43042 28756
rect 43257 28747 43315 28753
rect 43257 28744 43269 28747
rect 43036 28716 43269 28744
rect 43036 28704 43042 28716
rect 43257 28713 43269 28716
rect 43303 28713 43315 28747
rect 43257 28707 43315 28713
rect 39485 28679 39543 28685
rect 39485 28645 39497 28679
rect 39531 28676 39543 28679
rect 39531 28648 40448 28676
rect 39531 28645 39543 28648
rect 39485 28639 39543 28645
rect 40129 28611 40187 28617
rect 40129 28577 40141 28611
rect 40175 28608 40187 28611
rect 40218 28608 40224 28620
rect 40175 28580 40224 28608
rect 40175 28577 40187 28580
rect 40129 28571 40187 28577
rect 40218 28568 40224 28580
rect 40276 28568 40282 28620
rect 39209 28543 39267 28549
rect 39209 28509 39221 28543
rect 39255 28509 39267 28543
rect 39209 28503 39267 28509
rect 39298 28500 39304 28552
rect 39356 28549 39362 28552
rect 39356 28540 39364 28549
rect 39356 28512 39401 28540
rect 39356 28503 39364 28512
rect 39356 28500 39362 28503
rect 40034 28500 40040 28552
rect 40092 28500 40098 28552
rect 40310 28500 40316 28552
rect 40368 28500 40374 28552
rect 40420 28549 40448 28648
rect 40405 28543 40463 28549
rect 40405 28509 40417 28543
rect 40451 28509 40463 28543
rect 40405 28503 40463 28509
rect 41874 28500 41880 28552
rect 41932 28500 41938 28552
rect 35308 28444 38976 28472
rect 35308 28432 35314 28444
rect 39022 28432 39028 28484
rect 39080 28472 39086 28484
rect 39117 28475 39175 28481
rect 39117 28472 39129 28475
rect 39080 28444 39129 28472
rect 39080 28432 39086 28444
rect 39117 28441 39129 28444
rect 39163 28441 39175 28475
rect 39117 28435 39175 28441
rect 42144 28475 42202 28481
rect 42144 28441 42156 28475
rect 42190 28472 42202 28475
rect 42610 28472 42616 28484
rect 42190 28444 42616 28472
rect 42190 28441 42202 28444
rect 42144 28435 42202 28441
rect 42610 28432 42616 28444
rect 42668 28432 42674 28484
rect 34606 28404 34612 28416
rect 31312 28376 34612 28404
rect 34606 28364 34612 28376
rect 34664 28364 34670 28416
rect 36906 28364 36912 28416
rect 36964 28404 36970 28416
rect 37366 28404 37372 28416
rect 36964 28376 37372 28404
rect 36964 28364 36970 28376
rect 37366 28364 37372 28376
rect 37424 28364 37430 28416
rect 37461 28407 37519 28413
rect 37461 28373 37473 28407
rect 37507 28404 37519 28407
rect 39482 28404 39488 28416
rect 37507 28376 39488 28404
rect 37507 28373 37519 28376
rect 37461 28367 37519 28373
rect 39482 28364 39488 28376
rect 39540 28364 39546 28416
rect 40589 28407 40647 28413
rect 40589 28373 40601 28407
rect 40635 28404 40647 28407
rect 43070 28404 43076 28416
rect 40635 28376 43076 28404
rect 40635 28373 40647 28376
rect 40589 28367 40647 28373
rect 43070 28364 43076 28376
rect 43128 28364 43134 28416
rect 1104 28314 43884 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 43884 28314
rect 1104 28240 43884 28262
rect 7006 28160 7012 28212
rect 7064 28160 7070 28212
rect 12066 28160 12072 28212
rect 12124 28200 12130 28212
rect 14274 28200 14280 28212
rect 12124 28172 14280 28200
rect 12124 28160 12130 28172
rect 14274 28160 14280 28172
rect 14332 28160 14338 28212
rect 17310 28160 17316 28212
rect 17368 28160 17374 28212
rect 17678 28160 17684 28212
rect 17736 28160 17742 28212
rect 18414 28160 18420 28212
rect 18472 28200 18478 28212
rect 20898 28200 20904 28212
rect 18472 28172 20904 28200
rect 18472 28160 18478 28172
rect 20898 28160 20904 28172
rect 20956 28160 20962 28212
rect 21177 28203 21235 28209
rect 21177 28169 21189 28203
rect 21223 28200 21235 28203
rect 22833 28203 22891 28209
rect 22833 28200 22845 28203
rect 21223 28172 22845 28200
rect 21223 28169 21235 28172
rect 21177 28163 21235 28169
rect 22833 28169 22845 28172
rect 22879 28169 22891 28203
rect 22833 28163 22891 28169
rect 23201 28203 23259 28209
rect 23201 28169 23213 28203
rect 23247 28200 23259 28203
rect 24118 28200 24124 28212
rect 23247 28172 24124 28200
rect 23247 28169 23259 28172
rect 23201 28163 23259 28169
rect 24118 28160 24124 28172
rect 24176 28160 24182 28212
rect 24213 28203 24271 28209
rect 24213 28169 24225 28203
rect 24259 28200 24271 28203
rect 27982 28200 27988 28212
rect 24259 28172 27988 28200
rect 24259 28169 24271 28172
rect 24213 28163 24271 28169
rect 27982 28160 27988 28172
rect 28040 28160 28046 28212
rect 35250 28200 35256 28212
rect 28644 28172 35256 28200
rect 6914 28024 6920 28076
rect 6972 28024 6978 28076
rect 7834 28064 7840 28076
rect 7208 28036 7840 28064
rect 7208 28005 7236 28036
rect 7834 28024 7840 28036
rect 7892 28064 7898 28076
rect 8113 28067 8171 28073
rect 8113 28064 8125 28067
rect 7892 28036 8125 28064
rect 7892 28024 7898 28036
rect 8113 28033 8125 28036
rect 8159 28033 8171 28067
rect 8113 28027 8171 28033
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28064 8355 28067
rect 8938 28064 8944 28076
rect 8343 28036 8944 28064
rect 8343 28033 8355 28036
rect 8297 28027 8355 28033
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 11977 28067 12035 28073
rect 11977 28033 11989 28067
rect 12023 28064 12035 28067
rect 12084 28064 12112 28160
rect 28644 28144 28672 28172
rect 12253 28135 12311 28141
rect 12253 28101 12265 28135
rect 12299 28132 12311 28135
rect 13446 28132 13452 28144
rect 12299 28104 13452 28132
rect 12299 28101 12311 28104
rect 12253 28095 12311 28101
rect 13446 28092 13452 28104
rect 13504 28092 13510 28144
rect 14826 28092 14832 28144
rect 14884 28132 14890 28144
rect 14930 28135 14988 28141
rect 14930 28132 14942 28135
rect 14884 28104 14942 28132
rect 14884 28092 14890 28104
rect 14930 28101 14942 28104
rect 14976 28101 14988 28135
rect 14930 28095 14988 28101
rect 22922 28092 22928 28144
rect 22980 28132 22986 28144
rect 22980 28104 24532 28132
rect 22980 28092 22986 28104
rect 12023 28036 12112 28064
rect 12161 28067 12219 28073
rect 12023 28033 12035 28036
rect 11977 28027 12035 28033
rect 12161 28033 12173 28067
rect 12207 28033 12219 28067
rect 12161 28027 12219 28033
rect 7193 27999 7251 28005
rect 7193 27965 7205 27999
rect 7239 27965 7251 27999
rect 12176 27996 12204 28027
rect 12342 28024 12348 28076
rect 12400 28024 12406 28076
rect 13354 28024 13360 28076
rect 13412 28064 13418 28076
rect 14458 28064 14464 28076
rect 13412 28036 14464 28064
rect 13412 28024 13418 28036
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 19058 28064 19064 28076
rect 17788 28036 19064 28064
rect 12434 27996 12440 28008
rect 12176 27968 12440 27996
rect 7193 27959 7251 27965
rect 12434 27956 12440 27968
rect 12492 27956 12498 28008
rect 16666 27956 16672 28008
rect 16724 27996 16730 28008
rect 17788 28005 17816 28036
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 21082 28024 21088 28076
rect 21140 28024 21146 28076
rect 23566 28064 23572 28076
rect 23400 28036 23572 28064
rect 17773 27999 17831 28005
rect 17773 27996 17785 27999
rect 16724 27968 17785 27996
rect 16724 27956 16730 27968
rect 17773 27965 17785 27968
rect 17819 27965 17831 27999
rect 17773 27959 17831 27965
rect 17957 27999 18015 28005
rect 17957 27965 17969 27999
rect 18003 27996 18015 27999
rect 18230 27996 18236 28008
rect 18003 27968 18236 27996
rect 18003 27965 18015 27968
rect 17957 27959 18015 27965
rect 18230 27956 18236 27968
rect 18288 27956 18294 28008
rect 21358 27956 21364 28008
rect 21416 27956 21422 28008
rect 23290 27956 23296 28008
rect 23348 27956 23354 28008
rect 23400 28005 23428 28036
rect 23566 28024 23572 28036
rect 23624 28024 23630 28076
rect 23385 27999 23443 28005
rect 23385 27965 23397 27999
rect 23431 27965 23443 27999
rect 23385 27959 23443 27965
rect 24026 27956 24032 28008
rect 24084 27956 24090 28008
rect 24504 28005 24532 28104
rect 24670 28092 24676 28144
rect 24728 28132 24734 28144
rect 26513 28135 26571 28141
rect 26513 28132 26525 28135
rect 24728 28104 26525 28132
rect 24728 28092 24734 28104
rect 26513 28101 26525 28104
rect 26559 28132 26571 28135
rect 26878 28132 26884 28144
rect 26559 28104 26884 28132
rect 26559 28101 26571 28104
rect 26513 28095 26571 28101
rect 26878 28092 26884 28104
rect 26936 28092 26942 28144
rect 27706 28092 27712 28144
rect 27764 28132 27770 28144
rect 28626 28132 28632 28144
rect 27764 28104 28632 28132
rect 27764 28092 27770 28104
rect 28626 28092 28632 28104
rect 28684 28092 28690 28144
rect 29638 28092 29644 28144
rect 29696 28132 29702 28144
rect 31021 28135 31079 28141
rect 31021 28132 31033 28135
rect 29696 28104 31033 28132
rect 29696 28092 29702 28104
rect 31021 28101 31033 28104
rect 31067 28101 31079 28135
rect 31021 28095 31079 28101
rect 24578 28024 24584 28076
rect 24636 28024 24642 28076
rect 24946 28024 24952 28076
rect 25004 28064 25010 28076
rect 25406 28064 25412 28076
rect 25004 28036 25412 28064
rect 25004 28024 25010 28036
rect 25406 28024 25412 28036
rect 25464 28064 25470 28076
rect 26145 28067 26203 28073
rect 26145 28064 26157 28067
rect 25464 28036 26157 28064
rect 25464 28024 25470 28036
rect 26145 28033 26157 28036
rect 26191 28033 26203 28067
rect 26145 28027 26203 28033
rect 26329 28067 26387 28073
rect 26329 28033 26341 28067
rect 26375 28064 26387 28067
rect 27154 28064 27160 28076
rect 26375 28036 27160 28064
rect 26375 28033 26387 28036
rect 26329 28027 26387 28033
rect 24489 27999 24547 28005
rect 24489 27965 24501 27999
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 25038 27956 25044 28008
rect 25096 27996 25102 28008
rect 26344 27996 26372 28027
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 28169 28067 28227 28073
rect 28169 28033 28181 28067
rect 28215 28064 28227 28067
rect 29362 28064 29368 28076
rect 28215 28036 29368 28064
rect 28215 28033 28227 28036
rect 28169 28027 28227 28033
rect 29362 28024 29368 28036
rect 29420 28024 29426 28076
rect 29730 28024 29736 28076
rect 29788 28064 29794 28076
rect 30834 28064 30840 28076
rect 29788 28036 30840 28064
rect 29788 28024 29794 28036
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 30929 28067 30987 28073
rect 30929 28033 30941 28067
rect 30975 28064 30987 28067
rect 31128 28064 31156 28172
rect 35250 28160 35256 28172
rect 35308 28160 35314 28212
rect 38105 28203 38163 28209
rect 38105 28169 38117 28203
rect 38151 28200 38163 28203
rect 40310 28200 40316 28212
rect 38151 28172 40316 28200
rect 38151 28169 38163 28172
rect 38105 28163 38163 28169
rect 40310 28160 40316 28172
rect 40368 28160 40374 28212
rect 42610 28160 42616 28212
rect 42668 28160 42674 28212
rect 42978 28160 42984 28212
rect 43036 28160 43042 28212
rect 43070 28160 43076 28212
rect 43128 28160 43134 28212
rect 31754 28092 31760 28144
rect 31812 28132 31818 28144
rect 32677 28135 32735 28141
rect 32677 28132 32689 28135
rect 31812 28104 32689 28132
rect 31812 28092 31818 28104
rect 32677 28101 32689 28104
rect 32723 28101 32735 28135
rect 32677 28095 32735 28101
rect 33502 28092 33508 28144
rect 33560 28092 33566 28144
rect 36078 28132 36084 28144
rect 33888 28104 36084 28132
rect 30975 28036 31156 28064
rect 31205 28067 31263 28073
rect 30975 28033 30987 28036
rect 30929 28027 30987 28033
rect 31205 28033 31217 28067
rect 31251 28064 31263 28067
rect 31662 28064 31668 28076
rect 31251 28036 31668 28064
rect 31251 28033 31263 28036
rect 31205 28027 31263 28033
rect 31662 28024 31668 28036
rect 31720 28024 31726 28076
rect 32447 28067 32505 28073
rect 32447 28064 32459 28067
rect 32048 28036 32459 28064
rect 25096 27968 26372 27996
rect 25096 27956 25102 27968
rect 28350 27956 28356 28008
rect 28408 27956 28414 28008
rect 28442 27956 28448 28008
rect 28500 27956 28506 28008
rect 28534 27956 28540 28008
rect 28592 27956 28598 28008
rect 28626 27956 28632 28008
rect 28684 27956 28690 28008
rect 30852 27996 30880 28024
rect 32048 28008 32076 28036
rect 32447 28033 32459 28036
rect 32493 28033 32505 28067
rect 32447 28027 32505 28033
rect 32582 28024 32588 28076
rect 32640 28024 32646 28076
rect 32766 28024 32772 28076
rect 32824 28064 32830 28076
rect 32861 28067 32919 28073
rect 32861 28064 32873 28067
rect 32824 28036 32873 28064
rect 32824 28024 32830 28036
rect 32861 28033 32873 28036
rect 32907 28033 32919 28067
rect 33321 28067 33379 28073
rect 33321 28064 33333 28067
rect 32861 28027 32919 28033
rect 32968 28036 33333 28064
rect 32968 28008 32996 28036
rect 33321 28033 33333 28036
rect 33367 28033 33379 28067
rect 33321 28027 33379 28033
rect 33597 28067 33655 28073
rect 33597 28033 33609 28067
rect 33643 28033 33655 28067
rect 33597 28027 33655 28033
rect 32030 27996 32036 28008
rect 30852 27968 32036 27996
rect 32030 27956 32036 27968
rect 32088 27956 32094 28008
rect 32950 27956 32956 28008
rect 33008 27956 33014 28008
rect 33226 27956 33232 28008
rect 33284 27996 33290 28008
rect 33612 27996 33640 28027
rect 33284 27968 33640 27996
rect 33284 27956 33290 27968
rect 13814 27888 13820 27940
rect 13872 27888 13878 27940
rect 20806 27888 20812 27940
rect 20864 27928 20870 27940
rect 33888 27928 33916 28104
rect 36078 28092 36084 28104
rect 36136 28092 36142 28144
rect 36817 28135 36875 28141
rect 36817 28101 36829 28135
rect 36863 28132 36875 28135
rect 37090 28132 37096 28144
rect 36863 28104 37096 28132
rect 36863 28101 36875 28104
rect 36817 28095 36875 28101
rect 37090 28092 37096 28104
rect 37148 28092 37154 28144
rect 37461 28135 37519 28141
rect 37461 28101 37473 28135
rect 37507 28132 37519 28135
rect 37642 28132 37648 28144
rect 37507 28104 37648 28132
rect 37507 28101 37519 28104
rect 37461 28095 37519 28101
rect 37642 28092 37648 28104
rect 37700 28092 37706 28144
rect 38838 28092 38844 28144
rect 38896 28132 38902 28144
rect 39209 28135 39267 28141
rect 39209 28132 39221 28135
rect 38896 28104 39221 28132
rect 38896 28092 38902 28104
rect 39209 28101 39221 28104
rect 39255 28101 39267 28135
rect 39209 28095 39267 28101
rect 34241 28067 34299 28073
rect 34241 28033 34253 28067
rect 34287 28033 34299 28067
rect 34241 28027 34299 28033
rect 34256 27996 34284 28027
rect 34330 28024 34336 28076
rect 34388 28064 34394 28076
rect 34977 28067 35035 28073
rect 34977 28064 34989 28067
rect 34388 28036 34989 28064
rect 34388 28024 34394 28036
rect 34977 28033 34989 28036
rect 35023 28033 35035 28067
rect 34977 28027 35035 28033
rect 35066 28024 35072 28076
rect 35124 28064 35130 28076
rect 35161 28067 35219 28073
rect 35161 28064 35173 28067
rect 35124 28036 35173 28064
rect 35124 28024 35130 28036
rect 35161 28033 35173 28036
rect 35207 28064 35219 28067
rect 35618 28064 35624 28076
rect 35207 28036 35624 28064
rect 35207 28033 35219 28036
rect 35161 28027 35219 28033
rect 35618 28024 35624 28036
rect 35676 28024 35682 28076
rect 35986 28024 35992 28076
rect 36044 28024 36050 28076
rect 37826 28064 37832 28076
rect 37384 28036 37832 28064
rect 34422 27996 34428 28008
rect 34256 27968 34428 27996
rect 34422 27956 34428 27968
rect 34480 27956 34486 28008
rect 35253 27999 35311 28005
rect 35253 27965 35265 27999
rect 35299 27996 35311 27999
rect 37384 27996 37412 28036
rect 37826 28024 37832 28036
rect 37884 28024 37890 28076
rect 39482 28024 39488 28076
rect 39540 28024 39546 28076
rect 35299 27968 37412 27996
rect 37553 27999 37611 28005
rect 35299 27965 35311 27968
rect 35253 27959 35311 27965
rect 37553 27965 37565 27999
rect 37599 27965 37611 27999
rect 37553 27959 37611 27965
rect 20864 27900 33916 27928
rect 20864 27888 20870 27900
rect 36906 27888 36912 27940
rect 36964 27928 36970 27940
rect 37568 27928 37596 27959
rect 37918 27956 37924 28008
rect 37976 27956 37982 28008
rect 43254 27956 43260 28008
rect 43312 27956 43318 28008
rect 38746 27928 38752 27940
rect 36964 27900 38752 27928
rect 36964 27888 36970 27900
rect 38746 27888 38752 27900
rect 38804 27888 38810 27940
rect 5534 27820 5540 27872
rect 5592 27860 5598 27872
rect 6549 27863 6607 27869
rect 6549 27860 6561 27863
rect 5592 27832 6561 27860
rect 5592 27820 5598 27832
rect 6549 27829 6561 27832
rect 6595 27829 6607 27863
rect 6549 27823 6607 27829
rect 8202 27820 8208 27872
rect 8260 27820 8266 27872
rect 12526 27820 12532 27872
rect 12584 27820 12590 27872
rect 20714 27820 20720 27872
rect 20772 27820 20778 27872
rect 24118 27820 24124 27872
rect 24176 27860 24182 27872
rect 27706 27860 27712 27872
rect 24176 27832 27712 27860
rect 24176 27820 24182 27832
rect 27706 27820 27712 27832
rect 27764 27820 27770 27872
rect 27798 27820 27804 27872
rect 27856 27860 27862 27872
rect 28813 27863 28871 27869
rect 28813 27860 28825 27863
rect 27856 27832 28825 27860
rect 27856 27820 27862 27832
rect 28813 27829 28825 27832
rect 28859 27829 28871 27863
rect 28813 27823 28871 27829
rect 30653 27863 30711 27869
rect 30653 27829 30665 27863
rect 30699 27860 30711 27863
rect 30834 27860 30840 27872
rect 30699 27832 30840 27860
rect 30699 27829 30711 27832
rect 30653 27823 30711 27829
rect 30834 27820 30840 27832
rect 30892 27820 30898 27872
rect 32306 27820 32312 27872
rect 32364 27820 32370 27872
rect 32398 27820 32404 27872
rect 32456 27860 32462 27872
rect 33321 27863 33379 27869
rect 33321 27860 33333 27863
rect 32456 27832 33333 27860
rect 32456 27820 32462 27832
rect 33321 27829 33333 27832
rect 33367 27829 33379 27863
rect 33321 27823 33379 27829
rect 1104 27770 43884 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 43884 27770
rect 1104 27696 43884 27718
rect 22554 27656 22560 27668
rect 20640 27628 22560 27656
rect 17681 27591 17739 27597
rect 17681 27557 17693 27591
rect 17727 27588 17739 27591
rect 17954 27588 17960 27600
rect 17727 27560 17960 27588
rect 17727 27557 17739 27560
rect 17681 27551 17739 27557
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 7929 27523 7987 27529
rect 7929 27489 7941 27523
rect 7975 27520 7987 27523
rect 8202 27520 8208 27532
rect 7975 27492 8208 27520
rect 7975 27489 7987 27492
rect 7929 27483 7987 27489
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 11698 27480 11704 27532
rect 11756 27480 11762 27532
rect 20640 27464 20668 27628
rect 22554 27616 22560 27628
rect 22612 27656 22618 27668
rect 23198 27656 23204 27668
rect 22612 27628 23204 27656
rect 22612 27616 22618 27628
rect 23198 27616 23204 27628
rect 23256 27616 23262 27668
rect 25774 27616 25780 27668
rect 25832 27656 25838 27668
rect 25832 27628 25912 27656
rect 25832 27616 25838 27628
rect 23477 27591 23535 27597
rect 23477 27557 23489 27591
rect 23523 27588 23535 27591
rect 23566 27588 23572 27600
rect 23523 27560 23572 27588
rect 23523 27557 23535 27560
rect 23477 27551 23535 27557
rect 23566 27548 23572 27560
rect 23624 27588 23630 27600
rect 24670 27588 24676 27600
rect 23624 27560 24676 27588
rect 23624 27548 23630 27560
rect 24670 27548 24676 27560
rect 24728 27548 24734 27600
rect 25884 27588 25912 27628
rect 25958 27616 25964 27668
rect 26016 27616 26022 27668
rect 26068 27628 28994 27656
rect 26068 27588 26096 27628
rect 25884 27560 26096 27588
rect 21634 27480 21640 27532
rect 21692 27520 21698 27532
rect 24854 27520 24860 27532
rect 21692 27492 24860 27520
rect 21692 27480 21698 27492
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27452 5319 27455
rect 5307 27424 5672 27452
rect 5307 27421 5319 27424
rect 5261 27415 5319 27421
rect 5644 27396 5672 27424
rect 8018 27412 8024 27464
rect 8076 27412 8082 27464
rect 8110 27412 8116 27464
rect 8168 27452 8174 27464
rect 8297 27455 8355 27461
rect 8297 27452 8309 27455
rect 8168 27424 8309 27452
rect 8168 27412 8174 27424
rect 8297 27421 8309 27424
rect 8343 27421 8355 27455
rect 8297 27415 8355 27421
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9180 27424 9781 27452
rect 9180 27412 9186 27424
rect 9769 27421 9781 27424
rect 9815 27452 9827 27455
rect 10962 27452 10968 27464
rect 9815 27424 10968 27452
rect 9815 27421 9827 27424
rect 9769 27415 9827 27421
rect 10962 27412 10968 27424
rect 11020 27412 11026 27464
rect 16482 27452 16488 27464
rect 11063 27424 16488 27452
rect 5534 27393 5540 27396
rect 5528 27384 5540 27393
rect 5495 27356 5540 27384
rect 5528 27347 5540 27356
rect 5534 27344 5540 27347
rect 5592 27344 5598 27396
rect 5626 27344 5632 27396
rect 5684 27344 5690 27396
rect 6914 27384 6920 27396
rect 6656 27356 6920 27384
rect 6656 27325 6684 27356
rect 6914 27344 6920 27356
rect 6972 27384 6978 27396
rect 6972 27356 8248 27384
rect 6972 27344 6978 27356
rect 6641 27319 6699 27325
rect 6641 27285 6653 27319
rect 6687 27285 6699 27319
rect 6641 27279 6699 27285
rect 7742 27276 7748 27328
rect 7800 27276 7806 27328
rect 8220 27316 8248 27356
rect 8386 27344 8392 27396
rect 8444 27344 8450 27396
rect 10036 27387 10094 27393
rect 10036 27353 10048 27387
rect 10082 27384 10094 27387
rect 10318 27384 10324 27396
rect 10082 27356 10324 27384
rect 10082 27353 10094 27356
rect 10036 27347 10094 27353
rect 10318 27344 10324 27356
rect 10376 27344 10382 27396
rect 11063 27384 11091 27424
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 18782 27412 18788 27464
rect 18840 27452 18846 27464
rect 20346 27452 20352 27464
rect 18840 27424 20352 27452
rect 18840 27412 18846 27424
rect 20346 27412 20352 27424
rect 20404 27412 20410 27464
rect 20622 27412 20628 27464
rect 20680 27412 20686 27464
rect 20714 27412 20720 27464
rect 20772 27452 20778 27464
rect 20892 27455 20950 27461
rect 20772 27446 20852 27452
rect 20892 27446 20904 27455
rect 20772 27424 20904 27446
rect 20772 27412 20778 27424
rect 20824 27421 20904 27424
rect 20938 27421 20950 27455
rect 20824 27418 20950 27421
rect 20892 27415 20950 27418
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 23584 27461 23612 27492
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 23072 27424 23213 27452
rect 23072 27412 23078 27424
rect 23201 27421 23213 27424
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27421 23627 27455
rect 23569 27415 23627 27421
rect 10428 27356 11091 27384
rect 11968 27387 12026 27393
rect 10428 27316 10456 27356
rect 11968 27353 11980 27387
rect 12014 27384 12026 27387
rect 12158 27384 12164 27396
rect 12014 27356 12164 27384
rect 12014 27353 12026 27356
rect 11968 27347 12026 27353
rect 12158 27344 12164 27356
rect 12216 27344 12222 27396
rect 21174 27384 21180 27396
rect 12406 27356 21180 27384
rect 8220 27288 10456 27316
rect 10686 27276 10692 27328
rect 10744 27316 10750 27328
rect 11149 27319 11207 27325
rect 11149 27316 11161 27319
rect 10744 27288 11161 27316
rect 10744 27276 10750 27288
rect 11149 27285 11161 27288
rect 11195 27316 11207 27319
rect 12406 27316 12434 27356
rect 21174 27344 21180 27356
rect 21232 27384 21238 27396
rect 23308 27384 23336 27415
rect 24578 27412 24584 27464
rect 24636 27412 24642 27464
rect 24780 27461 24808 27492
rect 24854 27480 24860 27492
rect 24912 27480 24918 27532
rect 25884 27529 25912 27560
rect 26602 27548 26608 27600
rect 26660 27588 26666 27600
rect 27157 27591 27215 27597
rect 27157 27588 27169 27591
rect 26660 27560 27169 27588
rect 26660 27548 26666 27560
rect 27157 27557 27169 27560
rect 27203 27557 27215 27591
rect 28966 27588 28994 27628
rect 32766 27616 32772 27668
rect 32824 27656 32830 27668
rect 34514 27656 34520 27668
rect 32824 27628 34520 27656
rect 32824 27616 32830 27628
rect 34514 27616 34520 27628
rect 34572 27616 34578 27668
rect 35986 27616 35992 27668
rect 36044 27656 36050 27668
rect 37090 27656 37096 27668
rect 36044 27628 37096 27656
rect 36044 27616 36050 27628
rect 37090 27616 37096 27628
rect 37148 27616 37154 27668
rect 29546 27588 29552 27600
rect 28966 27560 29552 27588
rect 27157 27551 27215 27557
rect 29546 27548 29552 27560
rect 29604 27548 29610 27600
rect 30558 27548 30564 27600
rect 30616 27588 30622 27600
rect 31018 27588 31024 27600
rect 30616 27560 31024 27588
rect 30616 27548 30622 27560
rect 31018 27548 31024 27560
rect 31076 27588 31082 27600
rect 31570 27588 31576 27600
rect 31076 27560 31576 27588
rect 31076 27548 31082 27560
rect 31570 27548 31576 27560
rect 31628 27548 31634 27600
rect 32493 27591 32551 27597
rect 32493 27557 32505 27591
rect 32539 27588 32551 27591
rect 32950 27588 32956 27600
rect 32539 27560 32956 27588
rect 32539 27557 32551 27560
rect 32493 27551 32551 27557
rect 32950 27548 32956 27560
rect 33008 27548 33014 27600
rect 33962 27548 33968 27600
rect 34020 27588 34026 27600
rect 34020 27560 35388 27588
rect 34020 27548 34026 27560
rect 25869 27523 25927 27529
rect 25869 27489 25881 27523
rect 25915 27489 25927 27523
rect 25869 27483 25927 27489
rect 26970 27480 26976 27532
rect 27028 27520 27034 27532
rect 31938 27520 31944 27532
rect 27028 27492 28994 27520
rect 27028 27480 27034 27492
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27421 24823 27455
rect 25038 27452 25044 27464
rect 24765 27415 24823 27421
rect 24964 27424 25044 27452
rect 21232 27356 23336 27384
rect 21232 27344 21238 27356
rect 11195 27288 12434 27316
rect 11195 27285 11207 27288
rect 11149 27279 11207 27285
rect 13078 27276 13084 27328
rect 13136 27276 13142 27328
rect 16669 27319 16727 27325
rect 16669 27285 16681 27319
rect 16715 27316 16727 27319
rect 17126 27316 17132 27328
rect 16715 27288 17132 27316
rect 16715 27285 16727 27288
rect 16669 27279 16727 27285
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 18690 27276 18696 27328
rect 18748 27316 18754 27328
rect 20806 27316 20812 27328
rect 18748 27288 20812 27316
rect 18748 27276 18754 27288
rect 20806 27276 20812 27288
rect 20864 27276 20870 27328
rect 21082 27276 21088 27328
rect 21140 27316 21146 27328
rect 22005 27319 22063 27325
rect 22005 27316 22017 27319
rect 21140 27288 22017 27316
rect 21140 27276 21146 27288
rect 22005 27285 22017 27288
rect 22051 27316 22063 27319
rect 22738 27316 22744 27328
rect 22051 27288 22744 27316
rect 22051 27285 22063 27288
rect 22005 27279 22063 27285
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 23014 27276 23020 27328
rect 23072 27276 23078 27328
rect 23198 27276 23204 27328
rect 23256 27316 23262 27328
rect 24964 27316 24992 27424
rect 25038 27412 25044 27424
rect 25096 27412 25102 27464
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27421 26019 27455
rect 25961 27415 26019 27421
rect 25682 27344 25688 27396
rect 25740 27344 25746 27396
rect 25976 27384 26004 27415
rect 26510 27412 26516 27464
rect 26568 27452 26574 27464
rect 27062 27452 27068 27464
rect 26568 27424 27068 27452
rect 26568 27412 26574 27424
rect 27062 27412 27068 27424
rect 27120 27452 27126 27464
rect 27289 27455 27347 27461
rect 27289 27452 27301 27455
rect 27120 27424 27301 27452
rect 27120 27412 27126 27424
rect 27289 27421 27301 27424
rect 27335 27421 27347 27455
rect 27289 27415 27347 27421
rect 27430 27412 27436 27464
rect 27488 27412 27494 27464
rect 27522 27412 27528 27464
rect 27580 27412 27586 27464
rect 27706 27412 27712 27464
rect 27764 27412 27770 27464
rect 28966 27452 28994 27492
rect 30300 27492 31944 27520
rect 29730 27452 29736 27464
rect 28966 27424 29736 27452
rect 29730 27412 29736 27424
rect 29788 27452 29794 27464
rect 29871 27455 29929 27461
rect 29871 27452 29883 27455
rect 29788 27424 29883 27452
rect 29788 27412 29794 27424
rect 29871 27421 29883 27424
rect 29917 27421 29929 27455
rect 29871 27415 29929 27421
rect 30006 27412 30012 27464
rect 30064 27412 30070 27464
rect 30300 27461 30328 27492
rect 31938 27480 31944 27492
rect 31996 27480 32002 27532
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 32088 27492 32536 27520
rect 32088 27480 32094 27492
rect 30285 27455 30343 27461
rect 30285 27421 30297 27455
rect 30331 27421 30343 27455
rect 30285 27415 30343 27421
rect 30926 27412 30932 27464
rect 30984 27412 30990 27464
rect 31113 27455 31171 27461
rect 31113 27421 31125 27455
rect 31159 27452 31171 27455
rect 31662 27452 31668 27464
rect 31159 27424 31668 27452
rect 31159 27421 31171 27424
rect 31113 27415 31171 27421
rect 31662 27412 31668 27424
rect 31720 27412 31726 27464
rect 32508 27452 32536 27492
rect 32582 27480 32588 27532
rect 32640 27520 32646 27532
rect 33870 27520 33876 27532
rect 32640 27492 33876 27520
rect 32640 27480 32646 27492
rect 32784 27461 32812 27492
rect 33870 27480 33876 27492
rect 33928 27480 33934 27532
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 34848 27492 35112 27520
rect 34848 27480 34854 27492
rect 32677 27455 32735 27461
rect 32677 27452 32689 27455
rect 32508 27424 32689 27452
rect 32677 27421 32689 27424
rect 32723 27421 32735 27455
rect 32677 27415 32735 27421
rect 32769 27455 32827 27461
rect 32769 27421 32781 27455
rect 32815 27421 32827 27455
rect 32769 27415 32827 27421
rect 33045 27455 33103 27461
rect 33045 27421 33057 27455
rect 33091 27452 33103 27455
rect 33134 27452 33140 27464
rect 33091 27424 33140 27452
rect 33091 27421 33103 27424
rect 33045 27415 33103 27421
rect 33134 27412 33140 27424
rect 33192 27412 33198 27464
rect 34974 27412 34980 27464
rect 35032 27412 35038 27464
rect 35084 27461 35112 27492
rect 35360 27461 35388 27560
rect 35618 27548 35624 27600
rect 35676 27588 35682 27600
rect 35676 27560 37228 27588
rect 35676 27548 35682 27560
rect 35069 27455 35127 27461
rect 35069 27421 35081 27455
rect 35115 27421 35127 27455
rect 35069 27415 35127 27421
rect 35253 27455 35311 27461
rect 35253 27421 35265 27455
rect 35299 27421 35311 27455
rect 35253 27415 35311 27421
rect 35345 27455 35403 27461
rect 35345 27421 35357 27455
rect 35391 27421 35403 27455
rect 35345 27415 35403 27421
rect 29270 27384 29276 27396
rect 25976 27356 29276 27384
rect 29270 27344 29276 27356
rect 29328 27344 29334 27396
rect 30101 27387 30159 27393
rect 30101 27384 30113 27387
rect 29380 27356 30113 27384
rect 23256 27288 24992 27316
rect 23256 27276 23262 27288
rect 25222 27276 25228 27328
rect 25280 27276 25286 27328
rect 26145 27319 26203 27325
rect 26145 27285 26157 27319
rect 26191 27316 26203 27319
rect 26510 27316 26516 27328
rect 26191 27288 26516 27316
rect 26191 27285 26203 27288
rect 26145 27279 26203 27285
rect 26510 27276 26516 27288
rect 26568 27276 26574 27328
rect 27338 27276 27344 27328
rect 27396 27316 27402 27328
rect 29380 27316 29408 27356
rect 30101 27353 30113 27356
rect 30147 27384 30159 27387
rect 31754 27384 31760 27396
rect 30147 27356 31760 27384
rect 30147 27353 30159 27356
rect 30101 27347 30159 27353
rect 31754 27344 31760 27356
rect 31812 27384 31818 27396
rect 32861 27387 32919 27393
rect 32861 27384 32873 27387
rect 31812 27356 32873 27384
rect 31812 27344 31818 27356
rect 32784 27328 32812 27356
rect 32861 27353 32873 27356
rect 32907 27353 32919 27387
rect 32861 27347 32919 27353
rect 32950 27344 32956 27396
rect 33008 27384 33014 27396
rect 35268 27384 35296 27415
rect 33008 27356 35296 27384
rect 35360 27384 35388 27415
rect 36078 27412 36084 27464
rect 36136 27412 36142 27464
rect 36354 27412 36360 27464
rect 36412 27412 36418 27464
rect 36464 27461 36492 27560
rect 36449 27455 36507 27461
rect 36449 27421 36461 27455
rect 36495 27421 36507 27455
rect 36449 27415 36507 27421
rect 37090 27412 37096 27464
rect 37148 27412 37154 27464
rect 37200 27452 37228 27560
rect 38378 27548 38384 27600
rect 38436 27588 38442 27600
rect 39022 27588 39028 27600
rect 38436 27560 39028 27588
rect 38436 27548 38442 27560
rect 39022 27548 39028 27560
rect 39080 27548 39086 27600
rect 40126 27548 40132 27600
rect 40184 27588 40190 27600
rect 40221 27591 40279 27597
rect 40221 27588 40233 27591
rect 40184 27560 40233 27588
rect 40184 27548 40190 27560
rect 40221 27557 40233 27560
rect 40267 27557 40279 27591
rect 40221 27551 40279 27557
rect 37921 27523 37979 27529
rect 37921 27489 37933 27523
rect 37967 27520 37979 27523
rect 43165 27523 43223 27529
rect 37967 27492 41414 27520
rect 37967 27489 37979 27492
rect 37921 27483 37979 27489
rect 38657 27455 38715 27461
rect 38657 27452 38669 27455
rect 37200 27424 38669 27452
rect 38657 27421 38669 27424
rect 38703 27421 38715 27455
rect 38657 27415 38715 27421
rect 38749 27455 38807 27461
rect 38749 27421 38761 27455
rect 38795 27452 38807 27455
rect 38795 27424 38976 27452
rect 38795 27421 38807 27424
rect 38749 27415 38807 27421
rect 35434 27384 35440 27396
rect 35360 27356 35440 27384
rect 33008 27344 33014 27356
rect 35434 27344 35440 27356
rect 35492 27384 35498 27396
rect 36265 27387 36323 27393
rect 36265 27384 36277 27387
rect 35492 27356 36277 27384
rect 35492 27344 35498 27356
rect 36265 27353 36277 27356
rect 36311 27353 36323 27387
rect 36265 27347 36323 27353
rect 36722 27344 36728 27396
rect 36780 27384 36786 27396
rect 38841 27387 38899 27393
rect 38841 27384 38853 27387
rect 36780 27356 38853 27384
rect 36780 27344 36786 27356
rect 38841 27353 38853 27356
rect 38887 27353 38899 27387
rect 38948 27384 38976 27424
rect 39022 27412 39028 27464
rect 39080 27412 39086 27464
rect 40405 27455 40463 27461
rect 40405 27421 40417 27455
rect 40451 27452 40463 27455
rect 40678 27452 40684 27464
rect 40451 27424 40684 27452
rect 40451 27421 40463 27424
rect 40405 27415 40463 27421
rect 40678 27412 40684 27424
rect 40736 27412 40742 27464
rect 41386 27452 41414 27492
rect 43165 27489 43177 27523
rect 43211 27520 43223 27523
rect 43990 27520 43996 27532
rect 43211 27492 43996 27520
rect 43211 27489 43223 27492
rect 43165 27483 43223 27489
rect 43990 27480 43996 27492
rect 44048 27480 44054 27532
rect 41874 27452 41880 27464
rect 41386 27424 41880 27452
rect 41874 27412 41880 27424
rect 41932 27412 41938 27464
rect 42889 27455 42947 27461
rect 42889 27421 42901 27455
rect 42935 27452 42947 27455
rect 43070 27452 43076 27464
rect 42935 27424 43076 27452
rect 42935 27421 42947 27424
rect 42889 27415 42947 27421
rect 43070 27412 43076 27424
rect 43128 27412 43134 27464
rect 38948 27356 39712 27384
rect 38841 27347 38899 27353
rect 27396 27288 29408 27316
rect 27396 27276 27402 27288
rect 29730 27276 29736 27328
rect 29788 27276 29794 27328
rect 30926 27276 30932 27328
rect 30984 27316 30990 27328
rect 31021 27319 31079 27325
rect 31021 27316 31033 27319
rect 30984 27288 31033 27316
rect 30984 27276 30990 27288
rect 31021 27285 31033 27288
rect 31067 27285 31079 27319
rect 31021 27279 31079 27285
rect 32766 27276 32772 27328
rect 32824 27276 32830 27328
rect 34698 27276 34704 27328
rect 34756 27316 34762 27328
rect 35529 27319 35587 27325
rect 35529 27316 35541 27319
rect 34756 27288 35541 27316
rect 34756 27276 34762 27288
rect 35529 27285 35541 27288
rect 35575 27285 35587 27319
rect 35529 27279 35587 27285
rect 36078 27276 36084 27328
rect 36136 27316 36142 27328
rect 36633 27319 36691 27325
rect 36633 27316 36645 27319
rect 36136 27288 36645 27316
rect 36136 27276 36142 27288
rect 36633 27285 36645 27288
rect 36679 27285 36691 27319
rect 36633 27279 36691 27285
rect 38470 27276 38476 27328
rect 38528 27276 38534 27328
rect 39684 27316 39712 27356
rect 40310 27344 40316 27396
rect 40368 27384 40374 27396
rect 40589 27387 40647 27393
rect 40589 27384 40601 27387
rect 40368 27356 40601 27384
rect 40368 27344 40374 27356
rect 40589 27353 40601 27356
rect 40635 27353 40647 27387
rect 40589 27347 40647 27353
rect 40770 27316 40776 27328
rect 39684 27288 40776 27316
rect 40770 27276 40776 27288
rect 40828 27276 40834 27328
rect 1104 27226 43884 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 43884 27226
rect 1104 27152 43884 27174
rect 8110 27072 8116 27124
rect 8168 27112 8174 27124
rect 8168 27084 9260 27112
rect 8168 27072 8174 27084
rect 9122 27044 9128 27056
rect 7208 27016 9128 27044
rect 7208 26985 7236 27016
rect 9122 27004 9128 27016
rect 9180 27004 9186 27056
rect 7193 26979 7251 26985
rect 7193 26945 7205 26979
rect 7239 26945 7251 26979
rect 7193 26939 7251 26945
rect 7460 26979 7518 26985
rect 7460 26945 7472 26979
rect 7506 26976 7518 26979
rect 7742 26976 7748 26988
rect 7506 26948 7748 26976
rect 7506 26945 7518 26948
rect 7460 26939 7518 26945
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 9030 26936 9036 26988
rect 9088 26936 9094 26988
rect 9232 26985 9260 27084
rect 10318 27072 10324 27124
rect 10376 27072 10382 27124
rect 10686 27072 10692 27124
rect 10744 27072 10750 27124
rect 10781 27115 10839 27121
rect 10781 27081 10793 27115
rect 10827 27112 10839 27115
rect 10870 27112 10876 27124
rect 10827 27084 10876 27112
rect 10827 27081 10839 27084
rect 10781 27075 10839 27081
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 13446 27072 13452 27124
rect 13504 27072 13510 27124
rect 14918 27072 14924 27124
rect 14976 27112 14982 27124
rect 17218 27112 17224 27124
rect 14976 27084 17224 27112
rect 14976 27072 14982 27084
rect 17218 27072 17224 27084
rect 17276 27072 17282 27124
rect 18046 27072 18052 27124
rect 18104 27112 18110 27124
rect 18322 27112 18328 27124
rect 18104 27084 18328 27112
rect 18104 27072 18110 27084
rect 18322 27072 18328 27084
rect 18380 27112 18386 27124
rect 21266 27112 21272 27124
rect 18380 27084 21272 27112
rect 18380 27072 18386 27084
rect 21266 27072 21272 27084
rect 21324 27072 21330 27124
rect 21358 27072 21364 27124
rect 21416 27112 21422 27124
rect 22005 27115 22063 27121
rect 22005 27112 22017 27115
rect 21416 27084 22017 27112
rect 21416 27072 21422 27084
rect 22005 27081 22017 27084
rect 22051 27081 22063 27115
rect 22005 27075 22063 27081
rect 23106 27072 23112 27124
rect 23164 27112 23170 27124
rect 23201 27115 23259 27121
rect 23201 27112 23213 27115
rect 23164 27084 23213 27112
rect 23164 27072 23170 27084
rect 23201 27081 23213 27084
rect 23247 27081 23259 27115
rect 23201 27075 23259 27081
rect 25041 27115 25099 27121
rect 25041 27081 25053 27115
rect 25087 27112 25099 27115
rect 25777 27115 25835 27121
rect 25777 27112 25789 27115
rect 25087 27084 25789 27112
rect 25087 27081 25099 27084
rect 25041 27075 25099 27081
rect 25777 27081 25789 27084
rect 25823 27081 25835 27115
rect 25777 27075 25835 27081
rect 26234 27072 26240 27124
rect 26292 27112 26298 27124
rect 27982 27112 27988 27124
rect 26292 27084 27988 27112
rect 26292 27072 26298 27084
rect 27982 27072 27988 27084
rect 28040 27112 28046 27124
rect 28258 27112 28264 27124
rect 28040 27084 28264 27112
rect 28040 27072 28046 27084
rect 28258 27072 28264 27084
rect 28316 27072 28322 27124
rect 28350 27072 28356 27124
rect 28408 27072 28414 27124
rect 30558 27112 30564 27124
rect 28644 27084 30564 27112
rect 12336 27047 12394 27053
rect 12336 27013 12348 27047
rect 12382 27044 12394 27047
rect 12526 27044 12532 27056
rect 12382 27016 12532 27044
rect 12382 27013 12394 27016
rect 12336 27007 12394 27013
rect 12526 27004 12532 27016
rect 12584 27004 12590 27056
rect 16482 27004 16488 27056
rect 16540 27044 16546 27056
rect 24026 27044 24032 27056
rect 16540 27016 24032 27044
rect 16540 27004 16546 27016
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11698 26976 11704 26988
rect 11020 26948 11704 26976
rect 11020 26936 11026 26948
rect 11698 26936 11704 26948
rect 11756 26976 11762 26988
rect 12069 26979 12127 26985
rect 12069 26976 12081 26979
rect 11756 26948 12081 26976
rect 11756 26936 11762 26948
rect 12069 26945 12081 26948
rect 12115 26945 12127 26979
rect 12069 26939 12127 26945
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 15841 26979 15899 26985
rect 15841 26976 15853 26979
rect 14792 26948 15853 26976
rect 14792 26936 14798 26948
rect 15841 26945 15853 26948
rect 15887 26976 15899 26979
rect 16117 26979 16175 26985
rect 15887 26948 16068 26976
rect 15887 26945 15899 26948
rect 15841 26939 15899 26945
rect 10226 26868 10232 26920
rect 10284 26908 10290 26920
rect 10870 26908 10876 26920
rect 10284 26880 10876 26908
rect 10284 26868 10290 26880
rect 10870 26868 10876 26880
rect 10928 26868 10934 26920
rect 13446 26868 13452 26920
rect 13504 26908 13510 26920
rect 15933 26911 15991 26917
rect 15933 26908 15945 26911
rect 13504 26880 15945 26908
rect 13504 26868 13510 26880
rect 15933 26877 15945 26880
rect 15979 26877 15991 26911
rect 16040 26908 16068 26948
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16942 26976 16948 26988
rect 16163 26948 16948 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 18049 26979 18107 26985
rect 18049 26976 18061 26979
rect 17788 26948 18061 26976
rect 17034 26908 17040 26920
rect 16040 26880 17040 26908
rect 15933 26871 15991 26877
rect 17034 26868 17040 26880
rect 17092 26868 17098 26920
rect 17310 26868 17316 26920
rect 17368 26868 17374 26920
rect 17402 26868 17408 26920
rect 17460 26868 17466 26920
rect 8386 26800 8392 26852
rect 8444 26840 8450 26852
rect 8573 26843 8631 26849
rect 8573 26840 8585 26843
rect 8444 26812 8585 26840
rect 8444 26800 8450 26812
rect 8573 26809 8585 26812
rect 8619 26840 8631 26843
rect 16301 26843 16359 26849
rect 8619 26812 9812 26840
rect 8619 26809 8631 26812
rect 8573 26803 8631 26809
rect 9217 26775 9275 26781
rect 9217 26741 9229 26775
rect 9263 26772 9275 26775
rect 9674 26772 9680 26784
rect 9263 26744 9680 26772
rect 9263 26741 9275 26744
rect 9217 26735 9275 26741
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 9784 26772 9812 26812
rect 16301 26809 16313 26843
rect 16347 26840 16359 26843
rect 17678 26840 17684 26852
rect 16347 26812 17684 26840
rect 16347 26809 16359 26812
rect 16301 26803 16359 26809
rect 17678 26800 17684 26812
rect 17736 26800 17742 26852
rect 17788 26840 17816 26948
rect 18049 26945 18061 26948
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18414 26976 18420 26988
rect 18279 26948 18420 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18414 26936 18420 26948
rect 18472 26936 18478 26988
rect 19337 26979 19395 26985
rect 19337 26945 19349 26979
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26976 19855 26979
rect 20806 26976 20812 26988
rect 19843 26948 20812 26976
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 19352 26908 19380 26939
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 21082 26936 21088 26988
rect 21140 26936 21146 26988
rect 21174 26936 21180 26988
rect 21232 26936 21238 26988
rect 21266 26936 21272 26988
rect 21324 26982 21330 26988
rect 21361 26982 21419 26985
rect 21324 26979 21419 26982
rect 21324 26954 21373 26979
rect 21324 26936 21330 26954
rect 21361 26945 21373 26954
rect 21407 26945 21419 26979
rect 21361 26939 21419 26945
rect 21453 26982 21511 26985
rect 21453 26979 21588 26982
rect 21453 26945 21465 26979
rect 21499 26976 21588 26979
rect 21634 26976 21640 26988
rect 21499 26954 21640 26976
rect 21499 26945 21511 26954
rect 21560 26948 21640 26954
rect 21453 26939 21511 26945
rect 21634 26936 21640 26948
rect 21692 26936 21698 26988
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26976 22247 26979
rect 22922 26976 22928 26988
rect 22235 26948 22928 26976
rect 22235 26945 22247 26948
rect 22189 26939 22247 26945
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 23400 26985 23428 27016
rect 24026 27004 24032 27016
rect 24084 27004 24090 27056
rect 24949 27047 25007 27053
rect 24949 27013 24961 27047
rect 24995 27044 25007 27047
rect 27246 27044 27252 27056
rect 24995 27016 27252 27044
rect 24995 27013 25007 27016
rect 24949 27007 25007 27013
rect 27246 27004 27252 27016
rect 27304 27004 27310 27056
rect 28644 27044 28672 27084
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 31018 27072 31024 27124
rect 31076 27112 31082 27124
rect 31076 27084 31616 27112
rect 31076 27072 31082 27084
rect 28460 27016 28672 27044
rect 28721 27047 28779 27053
rect 23385 26979 23443 26985
rect 23385 26945 23397 26979
rect 23431 26945 23443 26979
rect 23385 26939 23443 26945
rect 23566 26936 23572 26988
rect 23624 26976 23630 26988
rect 23750 26976 23756 26988
rect 23624 26948 23756 26976
rect 23624 26936 23630 26948
rect 23750 26936 23756 26948
rect 23808 26936 23814 26988
rect 24854 26936 24860 26988
rect 24912 26976 24918 26988
rect 24912 26948 25360 26976
rect 24912 26936 24918 26948
rect 20901 26911 20959 26917
rect 20901 26908 20913 26911
rect 19352 26880 20913 26908
rect 20901 26877 20913 26880
rect 20947 26877 20959 26911
rect 20901 26871 20959 26877
rect 22373 26911 22431 26917
rect 22373 26877 22385 26911
rect 22419 26877 22431 26911
rect 22373 26871 22431 26877
rect 22465 26911 22523 26917
rect 22465 26877 22477 26911
rect 22511 26908 22523 26911
rect 23198 26908 23204 26920
rect 22511 26880 23204 26908
rect 22511 26877 22523 26880
rect 22465 26871 22523 26877
rect 19521 26843 19579 26849
rect 19521 26840 19533 26843
rect 17788 26812 19533 26840
rect 12250 26772 12256 26784
rect 9784 26744 12256 26772
rect 12250 26732 12256 26744
rect 12308 26732 12314 26784
rect 13078 26732 13084 26784
rect 13136 26772 13142 26784
rect 15841 26775 15899 26781
rect 15841 26772 15853 26775
rect 13136 26744 15853 26772
rect 13136 26732 13142 26744
rect 15841 26741 15853 26744
rect 15887 26772 15899 26775
rect 16574 26772 16580 26784
rect 15887 26744 16580 26772
rect 15887 26741 15899 26744
rect 15841 26735 15899 26741
rect 16574 26732 16580 26744
rect 16632 26732 16638 26784
rect 16850 26732 16856 26784
rect 16908 26732 16914 26784
rect 17402 26732 17408 26784
rect 17460 26772 17466 26784
rect 17788 26772 17816 26812
rect 19521 26809 19533 26812
rect 19567 26809 19579 26843
rect 20916 26840 20944 26871
rect 21174 26840 21180 26852
rect 20916 26812 21180 26840
rect 19521 26803 19579 26809
rect 21174 26800 21180 26812
rect 21232 26800 21238 26852
rect 21450 26800 21456 26852
rect 21508 26840 21514 26852
rect 22388 26840 22416 26871
rect 21508 26812 22416 26840
rect 21508 26800 21514 26812
rect 17460 26744 17816 26772
rect 17460 26732 17466 26744
rect 18046 26732 18052 26784
rect 18104 26732 18110 26784
rect 18966 26732 18972 26784
rect 19024 26772 19030 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 19024 26744 19073 26772
rect 19024 26732 19030 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 19061 26735 19119 26741
rect 19334 26732 19340 26784
rect 19392 26772 19398 26784
rect 19429 26775 19487 26781
rect 19429 26772 19441 26775
rect 19392 26744 19441 26772
rect 19392 26732 19398 26744
rect 19429 26741 19441 26744
rect 19475 26741 19487 26775
rect 19429 26735 19487 26741
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 20070 26772 20076 26784
rect 19668 26744 20076 26772
rect 19668 26732 19674 26744
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 20162 26732 20168 26784
rect 20220 26772 20226 26784
rect 22480 26772 22508 26871
rect 23198 26868 23204 26880
rect 23256 26868 23262 26920
rect 23661 26911 23719 26917
rect 23661 26877 23673 26911
rect 23707 26908 23719 26911
rect 24210 26908 24216 26920
rect 23707 26880 24216 26908
rect 23707 26877 23719 26880
rect 23661 26871 23719 26877
rect 24210 26868 24216 26880
rect 24268 26868 24274 26920
rect 25222 26868 25228 26920
rect 25280 26868 25286 26920
rect 25332 26908 25360 26948
rect 25958 26936 25964 26988
rect 26016 26976 26022 26988
rect 26145 26979 26203 26985
rect 26145 26976 26157 26979
rect 26016 26948 26157 26976
rect 26016 26936 26022 26948
rect 26145 26945 26157 26948
rect 26191 26976 26203 26979
rect 28460 26976 28488 27016
rect 28721 27013 28733 27047
rect 28767 27044 28779 27047
rect 30193 27047 30251 27053
rect 28767 27016 29500 27044
rect 28767 27013 28779 27016
rect 28721 27007 28779 27013
rect 29472 26988 29500 27016
rect 30193 27013 30205 27047
rect 30239 27044 30251 27047
rect 30466 27044 30472 27056
rect 30239 27016 30472 27044
rect 30239 27013 30251 27016
rect 30193 27007 30251 27013
rect 30466 27004 30472 27016
rect 30524 27004 30530 27056
rect 30650 27004 30656 27056
rect 30708 27044 30714 27056
rect 31588 27044 31616 27084
rect 31662 27072 31668 27124
rect 31720 27112 31726 27124
rect 31720 27084 34928 27112
rect 31720 27072 31726 27084
rect 30708 27016 31064 27044
rect 31588 27016 31984 27044
rect 30708 27004 30714 27016
rect 26191 26948 28488 26976
rect 26191 26945 26203 26948
rect 26145 26939 26203 26945
rect 28534 26936 28540 26988
rect 28592 26936 28598 26988
rect 28810 26936 28816 26988
rect 28868 26976 28874 26988
rect 29273 26979 29331 26985
rect 29273 26976 29285 26979
rect 28868 26948 29285 26976
rect 28868 26936 28874 26948
rect 29273 26945 29285 26948
rect 29319 26945 29331 26979
rect 29273 26939 29331 26945
rect 29362 26936 29368 26988
rect 29420 26936 29426 26988
rect 29454 26936 29460 26988
rect 29512 26936 29518 26988
rect 29822 26936 29828 26988
rect 29880 26976 29886 26988
rect 29880 26948 30788 26976
rect 29880 26936 29886 26948
rect 26329 26911 26387 26917
rect 26329 26908 26341 26911
rect 25332 26880 26341 26908
rect 26329 26877 26341 26880
rect 26375 26877 26387 26911
rect 26329 26871 26387 26877
rect 26786 26868 26792 26920
rect 26844 26908 26850 26920
rect 28902 26908 28908 26920
rect 26844 26880 28908 26908
rect 26844 26868 26850 26880
rect 28902 26868 28908 26880
rect 28960 26868 28966 26920
rect 30760 26908 30788 26948
rect 30834 26936 30840 26988
rect 30892 26936 30898 26988
rect 30926 26936 30932 26988
rect 30984 26936 30990 26988
rect 31036 26976 31064 27016
rect 31205 26979 31263 26985
rect 31205 26976 31217 26979
rect 31036 26948 31217 26976
rect 31205 26945 31217 26948
rect 31251 26976 31263 26979
rect 31846 26976 31852 26988
rect 31251 26948 31852 26976
rect 31251 26945 31263 26948
rect 31205 26939 31263 26945
rect 31846 26936 31852 26948
rect 31904 26936 31910 26988
rect 31956 26976 31984 27016
rect 32490 26976 32496 26988
rect 31956 26948 32496 26976
rect 32490 26936 32496 26948
rect 32548 26976 32554 26988
rect 32861 26979 32919 26985
rect 32861 26976 32873 26979
rect 32548 26948 32873 26976
rect 32548 26936 32554 26948
rect 32861 26945 32873 26948
rect 32907 26945 32919 26979
rect 32861 26939 32919 26945
rect 33045 26979 33103 26985
rect 33045 26945 33057 26979
rect 33091 26976 33103 26979
rect 33134 26976 33140 26988
rect 33091 26948 33140 26976
rect 33091 26945 33103 26948
rect 33045 26939 33103 26945
rect 33134 26936 33140 26948
rect 33192 26936 33198 26988
rect 33796 26948 34100 26976
rect 31297 26911 31355 26917
rect 31297 26908 31309 26911
rect 30760 26880 31309 26908
rect 31297 26877 31309 26880
rect 31343 26908 31355 26911
rect 31478 26908 31484 26920
rect 31343 26880 31484 26908
rect 31343 26877 31355 26880
rect 31297 26871 31355 26877
rect 31478 26868 31484 26880
rect 31536 26868 31542 26920
rect 31938 26868 31944 26920
rect 31996 26908 32002 26920
rect 33796 26908 33824 26948
rect 31996 26880 33824 26908
rect 34072 26908 34100 26948
rect 34146 26936 34152 26988
rect 34204 26936 34210 26988
rect 34238 26936 34244 26988
rect 34296 26976 34302 26988
rect 34333 26979 34391 26985
rect 34333 26976 34345 26979
rect 34296 26948 34345 26976
rect 34296 26936 34302 26948
rect 34333 26945 34345 26948
rect 34379 26976 34391 26979
rect 34790 26976 34796 26988
rect 34379 26948 34796 26976
rect 34379 26945 34391 26948
rect 34333 26939 34391 26945
rect 34790 26936 34796 26948
rect 34848 26936 34854 26988
rect 34900 26976 34928 27084
rect 34974 27072 34980 27124
rect 35032 27112 35038 27124
rect 36081 27115 36139 27121
rect 36081 27112 36093 27115
rect 35032 27084 36093 27112
rect 35032 27072 35038 27084
rect 36081 27081 36093 27084
rect 36127 27081 36139 27115
rect 36081 27075 36139 27081
rect 35894 27004 35900 27056
rect 35952 27044 35958 27056
rect 36722 27044 36728 27056
rect 35952 27016 36728 27044
rect 35952 27004 35958 27016
rect 36722 27004 36728 27016
rect 36780 27004 36786 27056
rect 37090 27004 37096 27056
rect 37148 27044 37154 27056
rect 37461 27047 37519 27053
rect 37461 27044 37473 27047
rect 37148 27016 37473 27044
rect 37148 27004 37154 27016
rect 37461 27013 37473 27016
rect 37507 27013 37519 27047
rect 37461 27007 37519 27013
rect 37734 27004 37740 27056
rect 37792 27044 37798 27056
rect 37792 27016 39344 27044
rect 37792 27004 37798 27016
rect 36357 26979 36415 26985
rect 36357 26976 36369 26979
rect 34900 26948 36369 26976
rect 36357 26945 36369 26948
rect 36403 26976 36415 26979
rect 37918 26976 37924 26988
rect 36403 26948 37924 26976
rect 36403 26945 36415 26948
rect 36357 26939 36415 26945
rect 37918 26936 37924 26948
rect 37976 26936 37982 26988
rect 38654 26936 38660 26988
rect 38712 26976 38718 26988
rect 39022 26985 39028 26988
rect 38841 26979 38899 26985
rect 38841 26976 38853 26979
rect 38712 26948 38853 26976
rect 38712 26936 38718 26948
rect 38841 26945 38853 26948
rect 38887 26945 38899 26979
rect 38841 26939 38899 26945
rect 38989 26979 39028 26985
rect 38989 26945 39001 26979
rect 38989 26939 39028 26945
rect 39022 26936 39028 26939
rect 39080 26936 39086 26988
rect 39114 26936 39120 26988
rect 39172 26936 39178 26988
rect 39316 26985 39344 27016
rect 39209 26979 39267 26985
rect 39209 26945 39221 26979
rect 39255 26945 39267 26979
rect 39209 26939 39267 26945
rect 39306 26979 39364 26985
rect 39306 26945 39318 26979
rect 39352 26945 39364 26979
rect 39306 26939 39364 26945
rect 36170 26908 36176 26920
rect 34072 26880 36176 26908
rect 31996 26868 32002 26880
rect 36170 26868 36176 26880
rect 36228 26868 36234 26920
rect 36265 26911 36323 26917
rect 36265 26877 36277 26911
rect 36311 26877 36323 26911
rect 36265 26871 36323 26877
rect 36633 26911 36691 26917
rect 36633 26877 36645 26911
rect 36679 26908 36691 26911
rect 36906 26908 36912 26920
rect 36679 26880 36912 26908
rect 36679 26877 36691 26880
rect 36633 26871 36691 26877
rect 22738 26800 22744 26852
rect 22796 26840 22802 26852
rect 22796 26812 26372 26840
rect 22796 26800 22802 26812
rect 20220 26744 22508 26772
rect 20220 26732 20226 26744
rect 23382 26732 23388 26784
rect 23440 26772 23446 26784
rect 24581 26775 24639 26781
rect 24581 26772 24593 26775
rect 23440 26744 24593 26772
rect 23440 26732 23446 26744
rect 24581 26741 24593 26744
rect 24627 26741 24639 26775
rect 24581 26735 24639 26741
rect 24670 26732 24676 26784
rect 24728 26772 24734 26784
rect 26234 26772 26240 26784
rect 24728 26744 26240 26772
rect 24728 26732 24734 26744
rect 26234 26732 26240 26744
rect 26292 26732 26298 26784
rect 26344 26772 26372 26812
rect 26878 26800 26884 26852
rect 26936 26840 26942 26852
rect 33778 26840 33784 26852
rect 26936 26812 33784 26840
rect 26936 26800 26942 26812
rect 33778 26800 33784 26812
rect 33836 26800 33842 26852
rect 36280 26840 36308 26871
rect 36906 26868 36912 26880
rect 36964 26868 36970 26920
rect 38194 26868 38200 26920
rect 38252 26868 38258 26920
rect 36814 26840 36820 26852
rect 34072 26812 36820 26840
rect 32950 26772 32956 26784
rect 26344 26744 32956 26772
rect 32950 26732 32956 26744
rect 33008 26732 33014 26784
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33410 26772 33416 26784
rect 33091 26744 33416 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33410 26732 33416 26744
rect 33468 26732 33474 26784
rect 34072 26781 34100 26812
rect 36814 26800 36820 26812
rect 36872 26800 36878 26852
rect 36998 26800 37004 26852
rect 37056 26840 37062 26852
rect 37734 26840 37740 26852
rect 37056 26812 37740 26840
rect 37056 26800 37062 26812
rect 37734 26800 37740 26812
rect 37792 26840 37798 26852
rect 39224 26840 39252 26939
rect 40770 26936 40776 26988
rect 40828 26976 40834 26988
rect 41794 26979 41852 26985
rect 41794 26976 41806 26979
rect 40828 26948 41806 26976
rect 40828 26936 40834 26948
rect 41794 26945 41806 26948
rect 41840 26945 41852 26979
rect 41794 26939 41852 26945
rect 41966 26936 41972 26988
rect 42024 26976 42030 26988
rect 42061 26979 42119 26985
rect 42061 26976 42073 26979
rect 42024 26948 42073 26976
rect 42024 26936 42030 26948
rect 42061 26945 42073 26948
rect 42107 26945 42119 26979
rect 42061 26939 42119 26945
rect 42978 26936 42984 26988
rect 43036 26936 43042 26988
rect 43070 26868 43076 26920
rect 43128 26868 43134 26920
rect 43254 26868 43260 26920
rect 43312 26868 43318 26920
rect 37792 26812 39252 26840
rect 37792 26800 37798 26812
rect 34057 26775 34115 26781
rect 34057 26741 34069 26775
rect 34103 26741 34115 26775
rect 34057 26735 34115 26741
rect 39482 26732 39488 26784
rect 39540 26732 39546 26784
rect 40034 26732 40040 26784
rect 40092 26772 40098 26784
rect 40681 26775 40739 26781
rect 40681 26772 40693 26775
rect 40092 26744 40693 26772
rect 40092 26732 40098 26744
rect 40681 26741 40693 26744
rect 40727 26741 40739 26775
rect 40681 26735 40739 26741
rect 42610 26732 42616 26784
rect 42668 26732 42674 26784
rect 1104 26682 43884 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 43884 26682
rect 1104 26608 43884 26630
rect 12158 26528 12164 26580
rect 12216 26528 12222 26580
rect 12250 26528 12256 26580
rect 12308 26568 12314 26580
rect 17402 26568 17408 26580
rect 12308 26540 17408 26568
rect 12308 26528 12314 26540
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 17494 26528 17500 26580
rect 17552 26568 17558 26580
rect 24857 26571 24915 26577
rect 24857 26568 24869 26571
rect 17552 26540 24869 26568
rect 17552 26528 17558 26540
rect 24857 26537 24869 26540
rect 24903 26568 24915 26571
rect 24903 26540 27752 26568
rect 24903 26537 24915 26540
rect 24857 26531 24915 26537
rect 9030 26460 9036 26512
rect 9088 26500 9094 26512
rect 9125 26503 9183 26509
rect 9125 26500 9137 26503
rect 9088 26472 9137 26500
rect 9088 26460 9094 26472
rect 9125 26469 9137 26472
rect 9171 26469 9183 26503
rect 13262 26500 13268 26512
rect 9125 26463 9183 26469
rect 12360 26472 13268 26500
rect 10962 26392 10968 26444
rect 11020 26392 11026 26444
rect 8110 26324 8116 26376
rect 8168 26364 8174 26376
rect 9309 26367 9367 26373
rect 9309 26364 9321 26367
rect 8168 26336 9321 26364
rect 8168 26324 8174 26336
rect 9309 26333 9321 26336
rect 9355 26333 9367 26367
rect 9309 26327 9367 26333
rect 9490 26324 9496 26376
rect 9548 26324 9554 26376
rect 9674 26324 9680 26376
rect 9732 26324 9738 26376
rect 12360 26373 12388 26472
rect 13262 26460 13268 26472
rect 13320 26460 13326 26512
rect 14369 26503 14427 26509
rect 14369 26469 14381 26503
rect 14415 26500 14427 26503
rect 14415 26472 14780 26500
rect 14415 26469 14427 26472
rect 14369 26463 14427 26469
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 12492 26404 12572 26432
rect 12492 26392 12498 26404
rect 12544 26373 12572 26404
rect 12345 26367 12403 26373
rect 12345 26333 12357 26367
rect 12391 26333 12403 26367
rect 12345 26327 12403 26333
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 12710 26324 12716 26376
rect 12768 26324 12774 26376
rect 14752 26364 14780 26472
rect 18322 26460 18328 26512
rect 18380 26460 18386 26512
rect 20824 26472 25544 26500
rect 16942 26392 16948 26444
rect 17000 26392 17006 26444
rect 17034 26392 17040 26444
rect 17092 26432 17098 26444
rect 19334 26432 19340 26444
rect 17092 26404 19340 26432
rect 17092 26392 17098 26404
rect 19334 26392 19340 26404
rect 19392 26392 19398 26444
rect 15194 26364 15200 26376
rect 14752 26336 15200 26364
rect 15194 26324 15200 26336
rect 15252 26324 15258 26376
rect 15746 26324 15752 26376
rect 15804 26324 15810 26376
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 17236 26336 17632 26364
rect 9398 26256 9404 26308
rect 9456 26256 9462 26308
rect 11701 26299 11759 26305
rect 11701 26265 11713 26299
rect 11747 26296 11759 26299
rect 12437 26299 12495 26305
rect 11747 26268 12388 26296
rect 11747 26265 11759 26268
rect 11701 26259 11759 26265
rect 12360 26228 12388 26268
rect 12437 26265 12449 26299
rect 12483 26296 12495 26299
rect 13078 26296 13084 26308
rect 12483 26268 13084 26296
rect 12483 26265 12495 26268
rect 12437 26259 12495 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 15504 26299 15562 26305
rect 15504 26265 15516 26299
rect 15550 26296 15562 26299
rect 15838 26296 15844 26308
rect 15550 26268 15844 26296
rect 15550 26265 15562 26268
rect 15504 26259 15562 26265
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 17037 26299 17095 26305
rect 17037 26265 17049 26299
rect 17083 26296 17095 26299
rect 17236 26296 17264 26336
rect 17083 26268 17264 26296
rect 17083 26265 17095 26268
rect 17037 26259 17095 26265
rect 17310 26256 17316 26308
rect 17368 26296 17374 26308
rect 17604 26296 17632 26336
rect 17678 26324 17684 26376
rect 17736 26364 17742 26376
rect 18141 26367 18199 26373
rect 18141 26364 18153 26367
rect 17736 26336 18153 26364
rect 17736 26324 17742 26336
rect 18141 26333 18153 26336
rect 18187 26333 18199 26367
rect 18141 26327 18199 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18782 26364 18788 26376
rect 18463 26336 18788 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 18782 26324 18788 26336
rect 18840 26324 18846 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 20622 26364 20628 26376
rect 19475 26336 20628 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 17368 26268 17540 26296
rect 17604 26268 17816 26296
rect 17368 26256 17374 26268
rect 12618 26228 12624 26240
rect 12360 26200 12624 26228
rect 12618 26188 12624 26200
rect 12676 26188 12682 26240
rect 17512 26237 17540 26268
rect 17497 26231 17555 26237
rect 17497 26197 17509 26231
rect 17543 26197 17555 26231
rect 17788 26228 17816 26268
rect 17862 26256 17868 26308
rect 17920 26296 17926 26308
rect 17957 26299 18015 26305
rect 17957 26296 17969 26299
rect 17920 26268 17969 26296
rect 17920 26256 17926 26268
rect 17957 26265 17969 26268
rect 18003 26265 18015 26299
rect 18322 26296 18328 26308
rect 17957 26259 18015 26265
rect 18064 26268 18328 26296
rect 18064 26228 18092 26268
rect 18322 26256 18328 26268
rect 18380 26296 18386 26308
rect 18690 26296 18696 26308
rect 18380 26268 18696 26296
rect 18380 26256 18386 26268
rect 18690 26256 18696 26268
rect 18748 26256 18754 26308
rect 17788 26200 18092 26228
rect 17497 26191 17555 26197
rect 18138 26188 18144 26240
rect 18196 26228 18202 26240
rect 19444 26228 19472 26327
rect 20622 26324 20628 26336
rect 20680 26324 20686 26376
rect 19518 26256 19524 26308
rect 19576 26296 19582 26308
rect 19674 26299 19732 26305
rect 19674 26296 19686 26299
rect 19576 26268 19686 26296
rect 19576 26256 19582 26268
rect 19674 26265 19686 26268
rect 19720 26265 19732 26299
rect 19674 26259 19732 26265
rect 18196 26200 19472 26228
rect 18196 26188 18202 26200
rect 20070 26188 20076 26240
rect 20128 26228 20134 26240
rect 20438 26228 20444 26240
rect 20128 26200 20444 26228
rect 20128 26188 20134 26200
rect 20438 26188 20444 26200
rect 20496 26228 20502 26240
rect 20824 26237 20852 26472
rect 23014 26392 23020 26444
rect 23072 26432 23078 26444
rect 23477 26435 23535 26441
rect 23477 26432 23489 26435
rect 23072 26404 23489 26432
rect 23072 26392 23078 26404
rect 23477 26401 23489 26404
rect 23523 26401 23535 26435
rect 25516 26432 25544 26472
rect 25590 26460 25596 26512
rect 25648 26500 25654 26512
rect 27617 26503 27675 26509
rect 27617 26500 27629 26503
rect 25648 26472 27629 26500
rect 25648 26460 25654 26472
rect 27617 26469 27629 26472
rect 27663 26469 27675 26503
rect 27724 26500 27752 26540
rect 28074 26528 28080 26580
rect 28132 26568 28138 26580
rect 32585 26571 32643 26577
rect 32585 26568 32597 26571
rect 28132 26540 32597 26568
rect 28132 26528 28138 26540
rect 32585 26537 32597 26540
rect 32631 26537 32643 26571
rect 32585 26531 32643 26537
rect 34606 26528 34612 26580
rect 34664 26568 34670 26580
rect 34977 26571 35035 26577
rect 34977 26568 34989 26571
rect 34664 26540 34989 26568
rect 34664 26528 34670 26540
rect 34977 26537 34989 26540
rect 35023 26537 35035 26571
rect 34977 26531 35035 26537
rect 35526 26528 35532 26580
rect 35584 26568 35590 26580
rect 37182 26568 37188 26580
rect 35584 26540 37188 26568
rect 35584 26528 35590 26540
rect 37182 26528 37188 26540
rect 37240 26528 37246 26580
rect 40770 26528 40776 26580
rect 40828 26528 40834 26580
rect 42978 26528 42984 26580
rect 43036 26568 43042 26580
rect 43349 26571 43407 26577
rect 43349 26568 43361 26571
rect 43036 26540 43361 26568
rect 43036 26528 43042 26540
rect 43349 26537 43361 26540
rect 43395 26537 43407 26571
rect 43349 26531 43407 26537
rect 29733 26503 29791 26509
rect 27724 26472 28212 26500
rect 27617 26463 27675 26469
rect 26878 26432 26884 26444
rect 25516 26404 26884 26432
rect 23477 26395 23535 26401
rect 26878 26392 26884 26404
rect 26936 26392 26942 26444
rect 27709 26435 27767 26441
rect 27709 26401 27721 26435
rect 27755 26432 27767 26435
rect 28074 26432 28080 26444
rect 27755 26404 28080 26432
rect 27755 26401 27767 26404
rect 27709 26395 27767 26401
rect 28074 26392 28080 26404
rect 28132 26392 28138 26444
rect 28184 26432 28212 26472
rect 29733 26469 29745 26503
rect 29779 26500 29791 26503
rect 30006 26500 30012 26512
rect 29779 26472 30012 26500
rect 29779 26469 29791 26472
rect 29733 26463 29791 26469
rect 30006 26460 30012 26472
rect 30064 26460 30070 26512
rect 31294 26460 31300 26512
rect 31352 26500 31358 26512
rect 34238 26500 34244 26512
rect 31352 26472 34244 26500
rect 31352 26460 31358 26472
rect 34238 26460 34244 26472
rect 34296 26460 34302 26512
rect 34333 26503 34391 26509
rect 34333 26469 34345 26503
rect 34379 26500 34391 26503
rect 35802 26500 35808 26512
rect 34379 26472 35808 26500
rect 34379 26469 34391 26472
rect 34333 26463 34391 26469
rect 35802 26460 35808 26472
rect 35860 26460 35866 26512
rect 38194 26460 38200 26512
rect 38252 26500 38258 26512
rect 38252 26472 42012 26500
rect 38252 26460 38258 26472
rect 41984 26444 42012 26472
rect 30190 26432 30196 26444
rect 28184 26404 30196 26432
rect 30190 26392 30196 26404
rect 30248 26432 30254 26444
rect 35986 26432 35992 26444
rect 30248 26404 35992 26432
rect 30248 26392 30254 26404
rect 35986 26392 35992 26404
rect 36044 26392 36050 26444
rect 39666 26432 39672 26444
rect 39040 26404 39672 26432
rect 21542 26324 21548 26376
rect 21600 26364 21606 26376
rect 23198 26364 23204 26376
rect 21600 26336 23204 26364
rect 21600 26324 21606 26336
rect 23198 26324 23204 26336
rect 23256 26364 23262 26376
rect 23293 26367 23351 26373
rect 23293 26364 23305 26367
rect 23256 26336 23305 26364
rect 23256 26324 23262 26336
rect 23293 26333 23305 26336
rect 23339 26333 23351 26367
rect 23293 26327 23351 26333
rect 23382 26324 23388 26376
rect 23440 26324 23446 26376
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26364 26387 26367
rect 26786 26364 26792 26376
rect 26375 26336 26792 26364
rect 26375 26333 26387 26336
rect 26329 26327 26387 26333
rect 26786 26324 26792 26336
rect 26844 26324 26850 26376
rect 26970 26324 26976 26376
rect 27028 26364 27034 26376
rect 27157 26367 27215 26373
rect 27157 26364 27169 26367
rect 27028 26336 27169 26364
rect 27028 26324 27034 26336
rect 27157 26333 27169 26336
rect 27203 26364 27215 26367
rect 27341 26367 27399 26373
rect 27203 26336 27292 26364
rect 27203 26333 27215 26336
rect 27157 26327 27215 26333
rect 20809 26231 20867 26237
rect 20809 26228 20821 26231
rect 20496 26200 20821 26228
rect 20496 26188 20502 26200
rect 20809 26197 20821 26200
rect 20855 26197 20867 26231
rect 20809 26191 20867 26197
rect 22922 26188 22928 26240
rect 22980 26188 22986 26240
rect 27264 26228 27292 26336
rect 27341 26333 27353 26367
rect 27387 26364 27399 26367
rect 27430 26364 27436 26376
rect 27387 26336 27436 26364
rect 27387 26333 27399 26336
rect 27341 26327 27399 26333
rect 27430 26324 27436 26336
rect 27488 26324 27494 26376
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 28721 26367 28779 26373
rect 28721 26333 28733 26367
rect 28767 26364 28779 26367
rect 28902 26364 28908 26376
rect 28767 26336 28908 26364
rect 28767 26333 28779 26336
rect 28721 26327 28779 26333
rect 28184 26296 28212 26327
rect 27724 26268 28212 26296
rect 27724 26228 27752 26268
rect 27264 26200 27752 26228
rect 27890 26188 27896 26240
rect 27948 26228 27954 26240
rect 28368 26228 28396 26327
rect 28902 26324 28908 26336
rect 28960 26324 28966 26376
rect 29730 26324 29736 26376
rect 29788 26324 29794 26376
rect 29822 26324 29828 26376
rect 29880 26364 29886 26376
rect 30009 26367 30067 26373
rect 30009 26364 30021 26367
rect 29880 26336 30021 26364
rect 29880 26324 29886 26336
rect 30009 26333 30021 26336
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 31202 26324 31208 26376
rect 31260 26324 31266 26376
rect 31478 26324 31484 26376
rect 31536 26364 31542 26376
rect 32766 26373 32772 26376
rect 32764 26364 32772 26373
rect 31536 26336 31754 26364
rect 32727 26336 32772 26364
rect 31536 26324 31542 26336
rect 28534 26256 28540 26308
rect 28592 26296 28598 26308
rect 29917 26299 29975 26305
rect 28592 26268 29868 26296
rect 28592 26256 28598 26268
rect 27948 26200 28396 26228
rect 27948 26188 27954 26200
rect 28626 26188 28632 26240
rect 28684 26188 28690 26240
rect 29840 26228 29868 26268
rect 29917 26265 29929 26299
rect 29963 26296 29975 26299
rect 30282 26296 30288 26308
rect 29963 26268 30288 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 30282 26256 30288 26268
rect 30340 26256 30346 26308
rect 31021 26299 31079 26305
rect 31021 26265 31033 26299
rect 31067 26296 31079 26299
rect 31110 26296 31116 26308
rect 31067 26268 31116 26296
rect 31067 26265 31079 26268
rect 31021 26259 31079 26265
rect 31110 26256 31116 26268
rect 31168 26256 31174 26308
rect 31389 26299 31447 26305
rect 31389 26265 31401 26299
rect 31435 26296 31447 26299
rect 31570 26296 31576 26308
rect 31435 26268 31576 26296
rect 31435 26265 31447 26268
rect 31389 26259 31447 26265
rect 31570 26256 31576 26268
rect 31628 26256 31634 26308
rect 31726 26296 31754 26336
rect 32764 26327 32772 26336
rect 32766 26324 32772 26327
rect 32824 26324 32830 26376
rect 32858 26324 32864 26376
rect 32916 26324 32922 26376
rect 33136 26367 33194 26373
rect 33136 26333 33148 26367
rect 33182 26333 33194 26367
rect 33136 26327 33194 26333
rect 32953 26299 33011 26305
rect 32953 26296 32965 26299
rect 31726 26268 32965 26296
rect 32953 26265 32965 26268
rect 32999 26296 33011 26299
rect 33151 26296 33179 26327
rect 33226 26324 33232 26376
rect 33284 26324 33290 26376
rect 33778 26324 33784 26376
rect 33836 26324 33842 26376
rect 33962 26324 33968 26376
rect 34020 26324 34026 26376
rect 34149 26367 34207 26373
rect 34149 26333 34161 26367
rect 34195 26364 34207 26367
rect 34238 26364 34244 26376
rect 34195 26336 34244 26364
rect 34195 26333 34207 26336
rect 34149 26327 34207 26333
rect 34238 26324 34244 26336
rect 34296 26324 34302 26376
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34480 26336 34897 26364
rect 34480 26324 34486 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 35158 26324 35164 26376
rect 35216 26324 35222 26376
rect 36446 26324 36452 26376
rect 36504 26373 36510 26376
rect 36504 26367 36553 26373
rect 36504 26333 36507 26367
rect 36541 26333 36553 26367
rect 36504 26327 36553 26333
rect 36504 26324 36510 26327
rect 36630 26324 36636 26376
rect 36688 26324 36694 26376
rect 36722 26324 36728 26376
rect 36780 26324 36786 26376
rect 36853 26367 36911 26373
rect 36853 26333 36865 26367
rect 36899 26333 36911 26367
rect 36853 26327 36911 26333
rect 33502 26296 33508 26308
rect 32999 26268 33088 26296
rect 33151 26268 33508 26296
rect 32999 26265 33011 26268
rect 32953 26259 33011 26265
rect 30926 26228 30932 26240
rect 29840 26200 30932 26228
rect 30926 26188 30932 26200
rect 30984 26188 30990 26240
rect 33060 26228 33088 26268
rect 33502 26256 33508 26268
rect 33560 26256 33566 26308
rect 34054 26256 34060 26308
rect 34112 26256 34118 26308
rect 35345 26299 35403 26305
rect 35345 26265 35357 26299
rect 35391 26296 35403 26299
rect 36170 26296 36176 26308
rect 35391 26268 36176 26296
rect 35391 26265 35403 26268
rect 35345 26259 35403 26265
rect 36170 26256 36176 26268
rect 36228 26256 36234 26308
rect 36868 26296 36896 26327
rect 36998 26324 37004 26376
rect 37056 26324 37062 26376
rect 37550 26324 37556 26376
rect 37608 26324 37614 26376
rect 37734 26364 37740 26376
rect 37660 26336 37740 26364
rect 37660 26305 37688 26336
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 37826 26324 37832 26376
rect 37884 26364 37890 26376
rect 37921 26367 37979 26373
rect 37921 26364 37933 26367
rect 37884 26336 37933 26364
rect 37884 26324 37890 26336
rect 37921 26333 37933 26336
rect 37967 26333 37979 26367
rect 37921 26327 37979 26333
rect 38013 26367 38071 26373
rect 38013 26333 38025 26367
rect 38059 26333 38071 26367
rect 38013 26327 38071 26333
rect 37645 26299 37703 26305
rect 37645 26296 37657 26299
rect 36464 26268 37657 26296
rect 33134 26228 33140 26240
rect 33060 26200 33140 26228
rect 33134 26188 33140 26200
rect 33192 26188 33198 26240
rect 33520 26228 33548 26256
rect 36464 26240 36492 26268
rect 37645 26265 37657 26268
rect 37691 26265 37703 26299
rect 38028 26296 38056 26327
rect 38654 26324 38660 26376
rect 38712 26324 38718 26376
rect 38805 26367 38863 26373
rect 38805 26333 38817 26367
rect 38851 26364 38863 26367
rect 39040 26364 39068 26404
rect 39666 26392 39672 26404
rect 39724 26392 39730 26444
rect 40310 26392 40316 26444
rect 40368 26392 40374 26444
rect 41966 26392 41972 26444
rect 42024 26392 42030 26444
rect 38851 26336 39068 26364
rect 39163 26367 39221 26373
rect 38851 26333 38863 26336
rect 38805 26327 38863 26333
rect 39163 26333 39175 26367
rect 39209 26364 39221 26367
rect 39298 26364 39304 26376
rect 39209 26336 39304 26364
rect 39209 26333 39221 26336
rect 39163 26327 39221 26333
rect 39298 26324 39304 26336
rect 39356 26324 39362 26376
rect 40405 26367 40463 26373
rect 40405 26333 40417 26367
rect 40451 26364 40463 26367
rect 40678 26364 40684 26376
rect 40451 26336 40684 26364
rect 40451 26333 40463 26336
rect 40405 26327 40463 26333
rect 40678 26324 40684 26336
rect 40736 26324 40742 26376
rect 42236 26367 42294 26373
rect 42236 26333 42248 26367
rect 42282 26364 42294 26367
rect 42610 26364 42616 26376
rect 42282 26336 42616 26364
rect 42282 26333 42294 26336
rect 42236 26327 42294 26333
rect 42610 26324 42616 26336
rect 42668 26324 42674 26376
rect 37645 26259 37703 26265
rect 37752 26268 38056 26296
rect 35158 26228 35164 26240
rect 33520 26200 35164 26228
rect 35158 26188 35164 26200
rect 35216 26228 35222 26240
rect 35526 26228 35532 26240
rect 35216 26200 35532 26228
rect 35216 26188 35222 26200
rect 35526 26188 35532 26200
rect 35584 26188 35590 26240
rect 36262 26188 36268 26240
rect 36320 26228 36326 26240
rect 36357 26231 36415 26237
rect 36357 26228 36369 26231
rect 36320 26200 36369 26228
rect 36320 26188 36326 26200
rect 36357 26197 36369 26200
rect 36403 26197 36415 26231
rect 36357 26191 36415 26197
rect 36446 26188 36452 26240
rect 36504 26188 36510 26240
rect 36538 26188 36544 26240
rect 36596 26228 36602 26240
rect 37752 26228 37780 26268
rect 38930 26256 38936 26308
rect 38988 26256 38994 26308
rect 39022 26256 39028 26308
rect 39080 26296 39086 26308
rect 42996 26296 43024 26528
rect 39080 26268 43024 26296
rect 39080 26256 39086 26268
rect 36596 26200 37780 26228
rect 38197 26231 38255 26237
rect 36596 26188 36602 26200
rect 38197 26197 38209 26231
rect 38243 26228 38255 26231
rect 38838 26228 38844 26240
rect 38243 26200 38844 26228
rect 38243 26197 38255 26200
rect 38197 26191 38255 26197
rect 38838 26188 38844 26200
rect 38896 26188 38902 26240
rect 39114 26188 39120 26240
rect 39172 26228 39178 26240
rect 39301 26231 39359 26237
rect 39301 26228 39313 26231
rect 39172 26200 39313 26228
rect 39172 26188 39178 26200
rect 39301 26197 39313 26200
rect 39347 26197 39359 26231
rect 39301 26191 39359 26197
rect 1104 26138 43884 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 43884 26138
rect 1104 26064 43884 26086
rect 15838 25984 15844 26036
rect 15896 25984 15902 26036
rect 19426 25984 19432 26036
rect 19484 26024 19490 26036
rect 19521 26027 19579 26033
rect 19521 26024 19533 26027
rect 19484 25996 19533 26024
rect 19484 25984 19490 25996
rect 19521 25993 19533 25996
rect 19567 25993 19579 26027
rect 19521 25987 19579 25993
rect 21266 25984 21272 26036
rect 21324 26024 21330 26036
rect 25225 26027 25283 26033
rect 25225 26024 25237 26027
rect 21324 25996 25237 26024
rect 21324 25984 21330 25996
rect 25225 25993 25237 25996
rect 25271 25993 25283 26027
rect 25225 25987 25283 25993
rect 25976 25996 27148 26024
rect 12618 25916 12624 25968
rect 12676 25956 12682 25968
rect 17405 25959 17463 25965
rect 17405 25956 17417 25959
rect 12676 25928 17417 25956
rect 12676 25916 12682 25928
rect 17405 25925 17417 25928
rect 17451 25956 17463 25959
rect 17494 25956 17500 25968
rect 17451 25928 17500 25956
rect 17451 25925 17463 25928
rect 17405 25919 17463 25925
rect 17494 25916 17500 25928
rect 17552 25916 17558 25968
rect 18138 25916 18144 25968
rect 18196 25916 18202 25968
rect 19153 25959 19211 25965
rect 19153 25925 19165 25959
rect 19199 25956 19211 25959
rect 20070 25956 20076 25968
rect 19199 25928 20076 25956
rect 19199 25925 19211 25928
rect 19153 25919 19211 25925
rect 20070 25916 20076 25928
rect 20128 25916 20134 25968
rect 22824 25959 22882 25965
rect 22824 25925 22836 25959
rect 22870 25956 22882 25959
rect 22922 25956 22928 25968
rect 22870 25928 22928 25956
rect 22870 25925 22882 25928
rect 22824 25919 22882 25925
rect 22922 25916 22928 25928
rect 22980 25916 22986 25968
rect 23198 25916 23204 25968
rect 23256 25956 23262 25968
rect 23934 25956 23940 25968
rect 23256 25928 23940 25956
rect 23256 25916 23262 25928
rect 23934 25916 23940 25928
rect 23992 25916 23998 25968
rect 15194 25848 15200 25900
rect 15252 25888 15258 25900
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15252 25860 15485 25888
rect 15252 25848 15258 25860
rect 15473 25857 15485 25860
rect 15519 25888 15531 25891
rect 19978 25888 19984 25900
rect 15519 25860 19984 25888
rect 15519 25857 15531 25860
rect 15473 25851 15531 25857
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 20162 25848 20168 25900
rect 20220 25848 20226 25900
rect 22554 25848 22560 25900
rect 22612 25848 22618 25900
rect 22664 25860 23612 25888
rect 11882 25780 11888 25832
rect 11940 25780 11946 25832
rect 15289 25823 15347 25829
rect 15289 25789 15301 25823
rect 15335 25789 15347 25823
rect 15289 25783 15347 25789
rect 15381 25823 15439 25829
rect 15381 25789 15393 25823
rect 15427 25820 15439 25823
rect 16850 25820 16856 25832
rect 15427 25792 16856 25820
rect 15427 25789 15439 25792
rect 15381 25783 15439 25789
rect 15304 25752 15332 25783
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 18966 25780 18972 25832
rect 19024 25780 19030 25832
rect 19058 25780 19064 25832
rect 19116 25780 19122 25832
rect 20070 25780 20076 25832
rect 20128 25820 20134 25832
rect 22664 25820 22692 25860
rect 20128 25792 22692 25820
rect 23584 25820 23612 25860
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25976 25897 26004 25996
rect 27120 25956 27148 25996
rect 27246 25984 27252 26036
rect 27304 25984 27310 26036
rect 28353 26027 28411 26033
rect 28353 25993 28365 26027
rect 28399 26024 28411 26027
rect 28810 26024 28816 26036
rect 28399 25996 28816 26024
rect 28399 25993 28411 25996
rect 28353 25987 28411 25993
rect 28810 25984 28816 25996
rect 28868 25984 28874 26036
rect 28902 25984 28908 26036
rect 28960 26024 28966 26036
rect 32769 26027 32827 26033
rect 32769 26024 32781 26027
rect 28960 25996 32781 26024
rect 28960 25984 28966 25996
rect 32769 25993 32781 25996
rect 32815 25993 32827 26027
rect 32769 25987 32827 25993
rect 32950 25984 32956 26036
rect 33008 26024 33014 26036
rect 36446 26024 36452 26036
rect 33008 25996 36452 26024
rect 33008 25984 33014 25996
rect 30742 25956 30748 25968
rect 27120 25928 30748 25956
rect 30742 25916 30748 25928
rect 30800 25916 30806 25968
rect 31294 25956 31300 25968
rect 31128 25928 31300 25956
rect 25593 25891 25651 25897
rect 25593 25888 25605 25891
rect 25004 25860 25605 25888
rect 25004 25848 25010 25860
rect 25593 25857 25605 25860
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25857 25743 25891
rect 25685 25851 25743 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 25700 25820 25728 25851
rect 23584 25792 25728 25820
rect 26252 25820 26280 25851
rect 26418 25848 26424 25900
rect 26476 25848 26482 25900
rect 26510 25848 26516 25900
rect 26568 25888 26574 25900
rect 27163 25891 27221 25897
rect 26568 25886 27016 25888
rect 27163 25886 27175 25891
rect 26568 25860 27175 25886
rect 26568 25848 26574 25860
rect 26988 25858 27175 25860
rect 27163 25857 27175 25858
rect 27209 25857 27221 25891
rect 27163 25851 27221 25857
rect 27353 25891 27411 25897
rect 27353 25857 27365 25891
rect 27399 25888 27411 25891
rect 27706 25888 27712 25900
rect 27399 25860 27712 25888
rect 27399 25857 27411 25860
rect 27353 25851 27411 25857
rect 27706 25848 27712 25860
rect 27764 25848 27770 25900
rect 27985 25891 28043 25897
rect 27985 25857 27997 25891
rect 28031 25888 28043 25891
rect 30650 25888 30656 25900
rect 28031 25860 30656 25888
rect 28031 25857 28043 25860
rect 27985 25851 28043 25857
rect 27246 25820 27252 25832
rect 26252 25792 27252 25820
rect 20128 25780 20134 25792
rect 27246 25780 27252 25792
rect 27304 25780 27310 25832
rect 17862 25752 17868 25764
rect 15304 25724 17868 25752
rect 17862 25712 17868 25724
rect 17920 25712 17926 25764
rect 18230 25712 18236 25764
rect 18288 25752 18294 25764
rect 18288 25724 22094 25752
rect 18288 25712 18294 25724
rect 20346 25644 20352 25696
rect 20404 25644 20410 25696
rect 22066 25684 22094 25724
rect 23492 25724 26832 25752
rect 23492 25684 23520 25724
rect 22066 25656 23520 25684
rect 23934 25644 23940 25696
rect 23992 25684 23998 25696
rect 24762 25684 24768 25696
rect 23992 25656 24768 25684
rect 23992 25644 23998 25656
rect 24762 25644 24768 25656
rect 24820 25644 24826 25696
rect 26804 25684 26832 25724
rect 26878 25712 26884 25764
rect 26936 25752 26942 25764
rect 28000 25752 28028 25851
rect 30650 25848 30656 25860
rect 30708 25848 30714 25900
rect 28074 25780 28080 25832
rect 28132 25780 28138 25832
rect 31128 25829 31156 25928
rect 31294 25916 31300 25928
rect 31352 25916 31358 25968
rect 31481 25959 31539 25965
rect 31481 25925 31493 25959
rect 31527 25956 31539 25959
rect 32674 25956 32680 25968
rect 31527 25928 32680 25956
rect 31527 25925 31539 25928
rect 31481 25919 31539 25925
rect 32674 25916 32680 25928
rect 32732 25916 32738 25968
rect 33042 25916 33048 25968
rect 33100 25916 33106 25968
rect 33134 25916 33140 25968
rect 33192 25916 33198 25968
rect 31202 25848 31208 25900
rect 31260 25888 31266 25900
rect 31386 25888 31392 25900
rect 31260 25860 31392 25888
rect 31260 25848 31266 25860
rect 31386 25848 31392 25860
rect 31444 25848 31450 25900
rect 32766 25848 32772 25900
rect 32824 25888 32830 25900
rect 33244 25897 33272 25996
rect 36446 25984 36452 25996
rect 36504 25984 36510 26036
rect 36538 25984 36544 26036
rect 36596 26024 36602 26036
rect 36633 26027 36691 26033
rect 36633 26024 36645 26027
rect 36596 25996 36645 26024
rect 36596 25984 36602 25996
rect 36633 25993 36645 25996
rect 36679 25993 36691 26027
rect 40034 26024 40040 26036
rect 36633 25987 36691 25993
rect 38764 25996 40040 26024
rect 35253 25959 35311 25965
rect 35253 25925 35265 25959
rect 35299 25956 35311 25959
rect 35986 25956 35992 25968
rect 35299 25928 35992 25956
rect 35299 25925 35311 25928
rect 35253 25919 35311 25925
rect 35986 25916 35992 25928
rect 36044 25956 36050 25968
rect 36044 25928 36492 25956
rect 36044 25916 36050 25928
rect 32907 25891 32965 25897
rect 32907 25888 32919 25891
rect 32824 25860 32919 25888
rect 32824 25848 32830 25860
rect 32907 25857 32919 25860
rect 32953 25857 32965 25891
rect 33244 25891 33323 25897
rect 33244 25860 33277 25891
rect 32907 25851 32965 25857
rect 33265 25857 33277 25860
rect 33311 25857 33323 25891
rect 33265 25851 33323 25857
rect 33410 25848 33416 25900
rect 33468 25848 33474 25900
rect 34422 25848 34428 25900
rect 34480 25888 34486 25900
rect 34517 25891 34575 25897
rect 34517 25888 34529 25891
rect 34480 25860 34529 25888
rect 34480 25848 34486 25860
rect 34517 25857 34529 25860
rect 34563 25857 34575 25891
rect 34517 25851 34575 25857
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 34977 25891 35035 25897
rect 34977 25888 34989 25891
rect 34848 25860 34989 25888
rect 34848 25848 34854 25860
rect 34977 25857 34989 25860
rect 35023 25857 35035 25891
rect 34977 25851 35035 25857
rect 35802 25848 35808 25900
rect 35860 25888 35866 25900
rect 36173 25891 36231 25897
rect 36173 25888 36185 25891
rect 35860 25860 36185 25888
rect 35860 25848 35866 25860
rect 36173 25857 36185 25860
rect 36219 25857 36231 25891
rect 36464 25888 36492 25928
rect 36635 25891 36693 25897
rect 36635 25888 36647 25891
rect 36464 25860 36647 25888
rect 36173 25851 36231 25857
rect 36635 25857 36647 25860
rect 36681 25888 36693 25891
rect 36998 25888 37004 25900
rect 36681 25860 37004 25888
rect 36681 25857 36693 25860
rect 36635 25851 36693 25857
rect 36998 25848 37004 25860
rect 37056 25848 37062 25900
rect 38654 25848 38660 25900
rect 38712 25888 38718 25900
rect 38764 25897 38792 25996
rect 40034 25984 40040 25996
rect 40092 25984 40098 26036
rect 39482 25916 39488 25968
rect 39540 25956 39546 25968
rect 39853 25959 39911 25965
rect 39853 25956 39865 25959
rect 39540 25928 39865 25956
rect 39540 25916 39546 25928
rect 39853 25925 39865 25928
rect 39899 25925 39911 25959
rect 39853 25919 39911 25925
rect 43162 25916 43168 25968
rect 43220 25916 43226 25968
rect 38749 25891 38807 25897
rect 38749 25888 38761 25891
rect 38712 25860 38761 25888
rect 38712 25848 38718 25860
rect 38749 25857 38761 25860
rect 38795 25857 38807 25891
rect 38749 25851 38807 25857
rect 38838 25848 38844 25900
rect 38896 25888 38902 25900
rect 39025 25891 39083 25897
rect 39025 25888 39037 25891
rect 38896 25860 39037 25888
rect 38896 25848 38902 25860
rect 39025 25857 39037 25860
rect 39071 25857 39083 25891
rect 39025 25851 39083 25857
rect 39114 25848 39120 25900
rect 39172 25848 39178 25900
rect 40126 25848 40132 25900
rect 40184 25888 40190 25900
rect 41138 25888 41144 25900
rect 40184 25860 41144 25888
rect 40184 25848 40190 25860
rect 41138 25848 41144 25860
rect 41196 25848 41202 25900
rect 42889 25891 42947 25897
rect 42889 25857 42901 25891
rect 42935 25888 42947 25891
rect 43070 25888 43076 25900
rect 42935 25860 43076 25888
rect 42935 25857 42947 25860
rect 42889 25851 42947 25857
rect 31113 25823 31171 25829
rect 31113 25789 31125 25823
rect 31159 25789 31171 25823
rect 31113 25783 31171 25789
rect 31220 25761 31248 25848
rect 35618 25780 35624 25832
rect 35676 25820 35682 25832
rect 37458 25820 37464 25832
rect 35676 25792 37464 25820
rect 35676 25780 35682 25792
rect 37458 25780 37464 25792
rect 37516 25780 37522 25832
rect 39301 25823 39359 25829
rect 39301 25789 39313 25823
rect 39347 25820 39359 25823
rect 42904 25820 42932 25851
rect 43070 25848 43076 25860
rect 43128 25848 43134 25900
rect 39347 25792 42932 25820
rect 39347 25789 39359 25792
rect 39301 25783 39359 25789
rect 26936 25724 28028 25752
rect 31205 25755 31263 25761
rect 26936 25712 26942 25724
rect 31205 25721 31217 25755
rect 31251 25721 31263 25755
rect 31205 25715 31263 25721
rect 36262 25712 36268 25764
rect 36320 25712 36326 25764
rect 38562 25752 38568 25764
rect 36745 25724 38568 25752
rect 27890 25684 27896 25696
rect 26804 25656 27896 25684
rect 27890 25644 27896 25656
rect 27948 25644 27954 25696
rect 31018 25644 31024 25696
rect 31076 25684 31082 25696
rect 31316 25687 31374 25693
rect 31316 25684 31328 25687
rect 31076 25656 31328 25684
rect 31076 25644 31082 25656
rect 31316 25653 31328 25656
rect 31362 25653 31374 25687
rect 31316 25647 31374 25653
rect 31938 25644 31944 25696
rect 31996 25684 32002 25696
rect 34054 25684 34060 25696
rect 31996 25656 34060 25684
rect 31996 25644 32002 25656
rect 34054 25644 34060 25656
rect 34112 25684 34118 25696
rect 36745 25684 36773 25724
rect 38562 25712 38568 25724
rect 38620 25712 38626 25764
rect 39853 25755 39911 25761
rect 39853 25721 39865 25755
rect 39899 25752 39911 25755
rect 40310 25752 40316 25764
rect 39899 25724 40316 25752
rect 39899 25721 39911 25724
rect 39853 25715 39911 25721
rect 40310 25712 40316 25724
rect 40368 25712 40374 25764
rect 34112 25656 36773 25684
rect 34112 25644 34118 25656
rect 36814 25644 36820 25696
rect 36872 25644 36878 25696
rect 38841 25687 38899 25693
rect 38841 25653 38853 25687
rect 38887 25684 38899 25687
rect 39022 25684 39028 25696
rect 38887 25656 39028 25684
rect 38887 25653 38899 25656
rect 38841 25647 38899 25653
rect 39022 25644 39028 25656
rect 39080 25644 39086 25696
rect 1104 25594 43884 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 43884 25594
rect 1104 25520 43884 25542
rect 10594 25440 10600 25492
rect 10652 25480 10658 25492
rect 11057 25483 11115 25489
rect 11057 25480 11069 25483
rect 10652 25452 11069 25480
rect 10652 25440 10658 25452
rect 11057 25449 11069 25452
rect 11103 25480 11115 25483
rect 18325 25483 18383 25489
rect 11103 25452 17908 25480
rect 11103 25449 11115 25452
rect 11057 25443 11115 25449
rect 10870 25372 10876 25424
rect 10928 25412 10934 25424
rect 12253 25415 12311 25421
rect 12253 25412 12265 25415
rect 10928 25384 12265 25412
rect 10928 25372 10934 25384
rect 12253 25381 12265 25384
rect 12299 25381 12311 25415
rect 12253 25375 12311 25381
rect 17773 25415 17831 25421
rect 17773 25381 17785 25415
rect 17819 25381 17831 25415
rect 17880 25412 17908 25452
rect 18325 25449 18337 25483
rect 18371 25480 18383 25483
rect 18598 25480 18604 25492
rect 18371 25452 18604 25480
rect 18371 25449 18383 25452
rect 18325 25443 18383 25449
rect 18598 25440 18604 25452
rect 18656 25440 18662 25492
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 19058 25480 19064 25492
rect 18739 25452 19064 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 19058 25440 19064 25452
rect 19116 25440 19122 25492
rect 19978 25440 19984 25492
rect 20036 25480 20042 25492
rect 21542 25480 21548 25492
rect 20036 25452 21548 25480
rect 20036 25440 20042 25452
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 24486 25440 24492 25492
rect 24544 25480 24550 25492
rect 25501 25483 25559 25489
rect 25501 25480 25513 25483
rect 24544 25452 25513 25480
rect 24544 25440 24550 25452
rect 25501 25449 25513 25452
rect 25547 25449 25559 25483
rect 25501 25443 25559 25449
rect 25961 25483 26019 25489
rect 25961 25449 25973 25483
rect 26007 25480 26019 25483
rect 27706 25480 27712 25492
rect 26007 25452 27712 25480
rect 26007 25449 26019 25452
rect 25961 25443 26019 25449
rect 27706 25440 27712 25452
rect 27764 25440 27770 25492
rect 31386 25440 31392 25492
rect 31444 25480 31450 25492
rect 32214 25480 32220 25492
rect 31444 25452 32220 25480
rect 31444 25440 31450 25452
rect 32214 25440 32220 25452
rect 32272 25440 32278 25492
rect 32861 25483 32919 25489
rect 32861 25449 32873 25483
rect 32907 25480 32919 25483
rect 33226 25480 33232 25492
rect 32907 25452 33232 25480
rect 32907 25449 32919 25452
rect 32861 25443 32919 25449
rect 33226 25440 33232 25452
rect 33284 25440 33290 25492
rect 36170 25440 36176 25492
rect 36228 25480 36234 25492
rect 36541 25483 36599 25489
rect 36541 25480 36553 25483
rect 36228 25452 36553 25480
rect 36228 25440 36234 25452
rect 36541 25449 36553 25452
rect 36587 25449 36599 25483
rect 36541 25443 36599 25449
rect 40678 25440 40684 25492
rect 40736 25440 40742 25492
rect 20070 25412 20076 25424
rect 17880 25384 20076 25412
rect 17773 25375 17831 25381
rect 13173 25347 13231 25353
rect 13173 25313 13185 25347
rect 13219 25344 13231 25347
rect 17788 25344 17816 25375
rect 20070 25372 20076 25384
rect 20128 25372 20134 25424
rect 22186 25372 22192 25424
rect 22244 25412 22250 25424
rect 26973 25415 27031 25421
rect 26973 25412 26985 25415
rect 22244 25384 26985 25412
rect 22244 25372 22250 25384
rect 26973 25381 26985 25384
rect 27019 25381 27031 25415
rect 26973 25375 27031 25381
rect 30009 25415 30067 25421
rect 30009 25381 30021 25415
rect 30055 25412 30067 25415
rect 30834 25412 30840 25424
rect 30055 25384 30840 25412
rect 30055 25381 30067 25384
rect 30009 25375 30067 25381
rect 30834 25372 30840 25384
rect 30892 25372 30898 25424
rect 31294 25372 31300 25424
rect 31352 25412 31358 25424
rect 31754 25412 31760 25424
rect 31352 25384 31760 25412
rect 31352 25372 31358 25384
rect 31754 25372 31760 25384
rect 31812 25372 31818 25424
rect 31846 25372 31852 25424
rect 31904 25372 31910 25424
rect 32876 25384 37688 25412
rect 13219 25316 17724 25344
rect 17788 25316 18552 25344
rect 13219 25313 13231 25316
rect 13173 25307 13231 25313
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 10962 25276 10968 25288
rect 9723 25248 10968 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 11826 25279 11884 25285
rect 11826 25276 11838 25279
rect 11063 25248 11838 25276
rect 9944 25211 10002 25217
rect 9944 25177 9956 25211
rect 9990 25208 10002 25211
rect 10226 25208 10232 25220
rect 9990 25180 10232 25208
rect 9990 25177 10002 25180
rect 9944 25171 10002 25177
rect 10226 25168 10232 25180
rect 10284 25168 10290 25220
rect 10686 25168 10692 25220
rect 10744 25208 10750 25220
rect 11063 25208 11091 25248
rect 11826 25245 11838 25248
rect 11872 25245 11884 25279
rect 11826 25239 11884 25245
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 12710 25276 12716 25288
rect 12391 25248 12716 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 12986 25236 12992 25288
rect 13044 25236 13050 25288
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 13906 25276 13912 25288
rect 13311 25248 13912 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 13906 25236 13912 25248
rect 13964 25236 13970 25288
rect 14366 25236 14372 25288
rect 14424 25276 14430 25288
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 14424 25248 14841 25276
rect 14424 25236 14430 25248
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15194 25236 15200 25288
rect 15252 25236 15258 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17129 25279 17187 25285
rect 17129 25276 17141 25279
rect 17092 25248 17141 25276
rect 17092 25236 17098 25248
rect 17129 25245 17141 25248
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17222 25279 17280 25285
rect 17222 25245 17234 25279
rect 17268 25245 17280 25279
rect 17222 25239 17280 25245
rect 13354 25208 13360 25220
rect 10744 25180 11091 25208
rect 11900 25180 13360 25208
rect 10744 25168 10750 25180
rect 11698 25100 11704 25152
rect 11756 25100 11762 25152
rect 11900 25149 11928 25180
rect 13354 25168 13360 25180
rect 13412 25168 13418 25220
rect 14921 25211 14979 25217
rect 14921 25177 14933 25211
rect 14967 25177 14979 25211
rect 14921 25171 14979 25177
rect 11885 25143 11943 25149
rect 11885 25109 11897 25143
rect 11931 25109 11943 25143
rect 11885 25103 11943 25109
rect 12802 25100 12808 25152
rect 12860 25100 12866 25152
rect 14645 25143 14703 25149
rect 14645 25109 14657 25143
rect 14691 25140 14703 25143
rect 14734 25140 14740 25152
rect 14691 25112 14740 25140
rect 14691 25109 14703 25112
rect 14645 25103 14703 25109
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 14936 25140 14964 25171
rect 15102 25168 15108 25220
rect 15160 25208 15166 25220
rect 17236 25208 17264 25239
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 17594 25279 17652 25285
rect 17594 25276 17606 25279
rect 17368 25248 17606 25276
rect 17368 25236 17374 25248
rect 17594 25245 17606 25248
rect 17640 25245 17652 25279
rect 17696 25276 17724 25316
rect 17696 25248 17908 25276
rect 17594 25239 17652 25245
rect 15160 25180 17264 25208
rect 17405 25211 17463 25217
rect 15160 25168 15166 25180
rect 17405 25177 17417 25211
rect 17451 25177 17463 25211
rect 17405 25171 17463 25177
rect 17497 25211 17555 25217
rect 17497 25177 17509 25211
rect 17543 25208 17555 25211
rect 17770 25208 17776 25220
rect 17543 25180 17776 25208
rect 17543 25177 17555 25180
rect 17497 25171 17555 25177
rect 15838 25140 15844 25152
rect 14936 25112 15844 25140
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 17420 25140 17448 25171
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 17880 25208 17908 25248
rect 18230 25236 18236 25288
rect 18288 25236 18294 25288
rect 18524 25285 18552 25316
rect 20622 25304 20628 25356
rect 20680 25304 20686 25356
rect 28166 25304 28172 25356
rect 28224 25344 28230 25356
rect 31938 25344 31944 25356
rect 28224 25316 31944 25344
rect 28224 25304 28230 25316
rect 31938 25304 31944 25316
rect 31996 25304 32002 25356
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 20346 25236 20352 25288
rect 20404 25276 20410 25288
rect 20881 25279 20939 25285
rect 20881 25276 20893 25279
rect 20404 25248 20893 25276
rect 20404 25236 20410 25248
rect 20881 25245 20893 25248
rect 20927 25245 20939 25279
rect 20881 25239 20939 25245
rect 25682 25236 25688 25288
rect 25740 25236 25746 25288
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25276 25835 25279
rect 25866 25276 25872 25288
rect 25823 25248 25872 25276
rect 25823 25245 25835 25248
rect 25777 25239 25835 25245
rect 25866 25236 25872 25248
rect 25924 25236 25930 25288
rect 27062 25236 27068 25288
rect 27120 25285 27126 25288
rect 27120 25279 27163 25285
rect 27151 25245 27163 25279
rect 27120 25239 27163 25245
rect 27120 25236 27126 25239
rect 27338 25236 27344 25288
rect 27396 25236 27402 25288
rect 27525 25279 27583 25285
rect 27525 25245 27537 25279
rect 27571 25276 27583 25279
rect 27890 25276 27896 25288
rect 27571 25248 27896 25276
rect 27571 25245 27583 25248
rect 27525 25239 27583 25245
rect 27890 25236 27896 25248
rect 27948 25276 27954 25288
rect 27948 25248 29684 25276
rect 27948 25236 27954 25248
rect 18782 25208 18788 25220
rect 17880 25180 18788 25208
rect 18782 25168 18788 25180
rect 18840 25168 18846 25220
rect 23290 25168 23296 25220
rect 23348 25208 23354 25220
rect 25501 25211 25559 25217
rect 25501 25208 25513 25211
rect 23348 25180 25513 25208
rect 23348 25168 23354 25180
rect 25501 25177 25513 25180
rect 25547 25208 25559 25211
rect 26878 25208 26884 25220
rect 25547 25180 26884 25208
rect 25547 25177 25559 25180
rect 25501 25171 25559 25177
rect 26878 25168 26884 25180
rect 26936 25168 26942 25220
rect 27249 25211 27307 25217
rect 27249 25177 27261 25211
rect 27295 25208 27307 25211
rect 28166 25208 28172 25220
rect 27295 25180 28172 25208
rect 27295 25177 27307 25180
rect 27249 25171 27307 25177
rect 28166 25168 28172 25180
rect 28224 25168 28230 25220
rect 29656 25208 29684 25248
rect 29730 25236 29736 25288
rect 29788 25236 29794 25288
rect 30558 25276 30564 25288
rect 29932 25248 30564 25276
rect 29932 25208 29960 25248
rect 30558 25236 30564 25248
rect 30616 25236 30622 25288
rect 30926 25236 30932 25288
rect 30984 25276 30990 25288
rect 31294 25276 31300 25288
rect 30984 25248 31300 25276
rect 30984 25236 30990 25248
rect 31294 25236 31300 25248
rect 31352 25236 31358 25288
rect 31478 25236 31484 25288
rect 31536 25276 31542 25288
rect 31573 25279 31631 25285
rect 31573 25276 31585 25279
rect 31536 25248 31585 25276
rect 31536 25236 31542 25248
rect 31573 25245 31585 25248
rect 31619 25245 31631 25279
rect 31573 25239 31631 25245
rect 31849 25279 31907 25285
rect 31849 25245 31861 25279
rect 31895 25276 31907 25279
rect 32306 25276 32312 25288
rect 31895 25248 32312 25276
rect 31895 25245 31907 25248
rect 31849 25239 31907 25245
rect 32306 25236 32312 25248
rect 32364 25236 32370 25288
rect 32490 25236 32496 25288
rect 32548 25276 32554 25288
rect 32876 25285 32904 25384
rect 34238 25304 34244 25356
rect 34296 25344 34302 25356
rect 36633 25347 36691 25353
rect 34296 25316 35945 25344
rect 34296 25304 34302 25316
rect 32677 25279 32735 25285
rect 32677 25276 32689 25279
rect 32548 25248 32689 25276
rect 32548 25236 32554 25248
rect 32677 25245 32689 25248
rect 32723 25245 32735 25279
rect 32677 25239 32735 25245
rect 32861 25279 32919 25285
rect 32861 25245 32873 25279
rect 32907 25245 32919 25279
rect 32861 25239 32919 25245
rect 35434 25236 35440 25288
rect 35492 25236 35498 25288
rect 35618 25285 35624 25288
rect 35585 25279 35624 25285
rect 35585 25245 35597 25279
rect 35585 25239 35624 25245
rect 35618 25236 35624 25239
rect 35676 25236 35682 25288
rect 35917 25285 35945 25316
rect 36633 25313 36645 25347
rect 36679 25344 36691 25347
rect 37553 25347 37611 25353
rect 37553 25344 37565 25347
rect 36679 25316 37565 25344
rect 36679 25313 36691 25316
rect 36633 25307 36691 25313
rect 37553 25313 37565 25316
rect 37599 25313 37611 25347
rect 37553 25307 37611 25313
rect 37660 25288 37688 25384
rect 39022 25304 39028 25356
rect 39080 25344 39086 25356
rect 40218 25344 40224 25356
rect 39080 25316 40224 25344
rect 39080 25304 39086 25316
rect 40218 25304 40224 25316
rect 40276 25304 40282 25356
rect 35902 25279 35960 25285
rect 35902 25245 35914 25279
rect 35948 25245 35960 25279
rect 36541 25279 36599 25285
rect 36541 25276 36553 25279
rect 35902 25239 35960 25245
rect 36096 25248 36553 25276
rect 29656 25180 29960 25208
rect 30009 25211 30067 25217
rect 30009 25177 30021 25211
rect 30055 25208 30067 25211
rect 30098 25208 30104 25220
rect 30055 25180 30104 25208
rect 30055 25177 30067 25180
rect 30009 25171 30067 25177
rect 30098 25168 30104 25180
rect 30156 25168 30162 25220
rect 30466 25168 30472 25220
rect 30524 25208 30530 25220
rect 30653 25211 30711 25217
rect 30653 25208 30665 25211
rect 30524 25180 30665 25208
rect 30524 25168 30530 25180
rect 30653 25177 30665 25180
rect 30699 25177 30711 25211
rect 30653 25171 30711 25177
rect 32766 25168 32772 25220
rect 32824 25208 32830 25220
rect 35710 25208 35716 25220
rect 32824 25180 35716 25208
rect 32824 25168 32830 25180
rect 35710 25168 35716 25180
rect 35768 25168 35774 25220
rect 35802 25168 35808 25220
rect 35860 25168 35866 25220
rect 18046 25140 18052 25152
rect 17420 25112 18052 25140
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 22005 25143 22063 25149
rect 22005 25109 22017 25143
rect 22051 25140 22063 25143
rect 26970 25140 26976 25152
rect 22051 25112 26976 25140
rect 22051 25109 22063 25112
rect 22005 25103 22063 25109
rect 26970 25100 26976 25112
rect 27028 25100 27034 25152
rect 29270 25100 29276 25152
rect 29328 25140 29334 25152
rect 29825 25143 29883 25149
rect 29825 25140 29837 25143
rect 29328 25112 29837 25140
rect 29328 25100 29334 25112
rect 29825 25109 29837 25112
rect 29871 25140 29883 25143
rect 30282 25140 30288 25152
rect 29871 25112 30288 25140
rect 29871 25109 29883 25112
rect 29825 25103 29883 25109
rect 30282 25100 30288 25112
rect 30340 25100 30346 25152
rect 31386 25100 31392 25152
rect 31444 25140 31450 25152
rect 36096 25149 36124 25248
rect 36541 25245 36553 25248
rect 36587 25245 36599 25279
rect 36541 25239 36599 25245
rect 36722 25236 36728 25288
rect 36780 25276 36786 25288
rect 36906 25276 36912 25288
rect 36780 25248 36912 25276
rect 36780 25236 36786 25248
rect 36906 25236 36912 25248
rect 36964 25276 36970 25288
rect 37461 25279 37519 25285
rect 37461 25276 37473 25279
rect 36964 25248 37473 25276
rect 36964 25236 36970 25248
rect 37461 25245 37473 25248
rect 37507 25245 37519 25279
rect 37461 25239 37519 25245
rect 37642 25236 37648 25288
rect 37700 25236 37706 25288
rect 38930 25236 38936 25288
rect 38988 25236 38994 25288
rect 39206 25236 39212 25288
rect 39264 25236 39270 25288
rect 39298 25236 39304 25288
rect 39356 25236 39362 25288
rect 39485 25279 39543 25285
rect 39485 25245 39497 25279
rect 39531 25276 39543 25279
rect 42889 25279 42947 25285
rect 42889 25276 42901 25279
rect 39531 25248 42901 25276
rect 39531 25245 39543 25248
rect 39485 25239 39543 25245
rect 42889 25245 42901 25248
rect 42935 25276 42947 25279
rect 43070 25276 43076 25288
rect 42935 25248 43076 25276
rect 42935 25245 42947 25248
rect 42889 25239 42947 25245
rect 43070 25236 43076 25248
rect 43128 25236 43134 25288
rect 40310 25168 40316 25220
rect 40368 25168 40374 25220
rect 40402 25168 40408 25220
rect 40460 25208 40466 25220
rect 40497 25211 40555 25217
rect 40497 25208 40509 25211
rect 40460 25180 40509 25208
rect 40460 25168 40466 25180
rect 40497 25177 40509 25180
rect 40543 25177 40555 25211
rect 40497 25171 40555 25177
rect 43165 25211 43223 25217
rect 43165 25177 43177 25211
rect 43211 25208 43223 25211
rect 43990 25208 43996 25220
rect 43211 25180 43996 25208
rect 43211 25177 43223 25180
rect 43165 25171 43223 25177
rect 43990 25168 43996 25180
rect 44048 25168 44054 25220
rect 31665 25143 31723 25149
rect 31665 25140 31677 25143
rect 31444 25112 31677 25140
rect 31444 25100 31450 25112
rect 31665 25109 31677 25112
rect 31711 25109 31723 25143
rect 31665 25103 31723 25109
rect 36081 25143 36139 25149
rect 36081 25109 36093 25143
rect 36127 25109 36139 25143
rect 36081 25103 36139 25109
rect 36906 25100 36912 25152
rect 36964 25100 36970 25152
rect 1104 25050 43884 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 43884 25050
rect 1104 24976 43884 24998
rect 10226 24896 10232 24948
rect 10284 24896 10290 24948
rect 10594 24896 10600 24948
rect 10652 24896 10658 24948
rect 17310 24896 17316 24948
rect 17368 24936 17374 24948
rect 25682 24936 25688 24948
rect 17368 24908 25688 24936
rect 17368 24896 17374 24908
rect 25682 24896 25688 24908
rect 25740 24896 25746 24948
rect 25866 24896 25872 24948
rect 25924 24936 25930 24948
rect 25924 24908 28488 24936
rect 25924 24896 25930 24908
rect 12802 24877 12808 24880
rect 12796 24868 12808 24877
rect 12763 24840 12808 24868
rect 12796 24831 12808 24840
rect 12802 24828 12808 24831
rect 12860 24828 12866 24880
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 17773 24871 17831 24877
rect 17773 24868 17785 24871
rect 17552 24840 17785 24868
rect 17552 24828 17558 24840
rect 17773 24837 17785 24840
rect 17819 24837 17831 24871
rect 24946 24868 24952 24880
rect 17773 24831 17831 24837
rect 23124 24840 23336 24868
rect 9030 24760 9036 24812
rect 9088 24809 9094 24812
rect 9088 24800 9100 24809
rect 9088 24772 9133 24800
rect 9088 24763 9100 24772
rect 9088 24760 9094 24763
rect 10686 24760 10692 24812
rect 10744 24760 10750 24812
rect 14734 24809 14740 24812
rect 14728 24800 14740 24809
rect 14695 24772 14740 24800
rect 14728 24763 14740 24772
rect 14734 24760 14740 24763
rect 14792 24760 14798 24812
rect 19705 24803 19763 24809
rect 19705 24769 19717 24803
rect 19751 24800 19763 24803
rect 21082 24800 21088 24812
rect 19751 24772 21088 24800
rect 19751 24769 19763 24772
rect 19705 24763 19763 24769
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 22370 24760 22376 24812
rect 22428 24760 22434 24812
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 23124 24800 23152 24840
rect 22756 24772 23152 24800
rect 23201 24803 23259 24809
rect 9309 24735 9367 24741
rect 9309 24701 9321 24735
rect 9355 24701 9367 24735
rect 9309 24695 9367 24701
rect 9324 24664 9352 24695
rect 10870 24692 10876 24744
rect 10928 24692 10934 24744
rect 11882 24692 11888 24744
rect 11940 24732 11946 24744
rect 12529 24735 12587 24741
rect 12529 24732 12541 24735
rect 11940 24704 12541 24732
rect 11940 24692 11946 24704
rect 12529 24701 12541 24704
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 14461 24735 14519 24741
rect 14461 24701 14473 24735
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 11054 24664 11060 24676
rect 9324 24636 11060 24664
rect 11054 24624 11060 24636
rect 11112 24624 11118 24676
rect 7929 24599 7987 24605
rect 7929 24565 7941 24599
rect 7975 24596 7987 24599
rect 8294 24596 8300 24608
rect 7975 24568 8300 24596
rect 7975 24565 7987 24568
rect 7929 24559 7987 24565
rect 8294 24556 8300 24568
rect 8352 24556 8358 24608
rect 13906 24556 13912 24608
rect 13964 24556 13970 24608
rect 14476 24596 14504 24695
rect 16850 24692 16856 24744
rect 16908 24732 16914 24744
rect 16945 24735 17003 24741
rect 16945 24732 16957 24735
rect 16908 24704 16957 24732
rect 16908 24692 16914 24704
rect 16945 24701 16957 24704
rect 16991 24701 17003 24735
rect 16945 24695 17003 24701
rect 19889 24735 19947 24741
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 22388 24732 22416 24760
rect 22756 24744 22784 24772
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23308 24800 23336 24840
rect 23676 24840 24952 24868
rect 23676 24809 23704 24840
rect 24946 24828 24952 24840
rect 25004 24828 25010 24880
rect 25700 24868 25728 24896
rect 28460 24868 28488 24908
rect 28534 24896 28540 24948
rect 28592 24936 28598 24948
rect 33502 24936 33508 24948
rect 28592 24908 33508 24936
rect 28592 24896 28598 24908
rect 33502 24896 33508 24908
rect 33560 24896 33566 24948
rect 35802 24896 35808 24948
rect 35860 24936 35866 24948
rect 38930 24936 38936 24948
rect 35860 24908 38936 24936
rect 35860 24896 35866 24908
rect 38930 24896 38936 24908
rect 38988 24896 38994 24948
rect 39209 24939 39267 24945
rect 39209 24905 39221 24939
rect 39255 24936 39267 24939
rect 39298 24936 39304 24948
rect 39255 24908 39304 24936
rect 39255 24905 39267 24908
rect 39209 24899 39267 24905
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 43070 24896 43076 24948
rect 43128 24896 43134 24948
rect 31386 24868 31392 24880
rect 25700 24840 27568 24868
rect 28460 24840 31392 24868
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23308 24772 23673 24800
rect 23201 24763 23259 24769
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 22738 24732 22744 24744
rect 22388 24704 22744 24732
rect 19889 24695 19947 24701
rect 15746 24664 15752 24676
rect 15396 24636 15752 24664
rect 15396 24596 15424 24636
rect 15746 24624 15752 24636
rect 15804 24664 15810 24676
rect 16868 24664 16896 24692
rect 19904 24664 19932 24695
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 23216 24732 23244 24763
rect 23750 24760 23756 24812
rect 23808 24760 23814 24812
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24765 24803 24823 24809
rect 24765 24800 24777 24803
rect 23983 24772 24777 24800
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 24765 24769 24777 24772
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 23474 24732 23480 24744
rect 23216 24704 23480 24732
rect 23474 24692 23480 24704
rect 23532 24732 23538 24744
rect 23952 24732 23980 24763
rect 24854 24732 24860 24744
rect 23532 24704 23980 24732
rect 24136 24704 24860 24732
rect 23532 24692 23538 24704
rect 22830 24664 22836 24676
rect 15804 24636 16896 24664
rect 18156 24636 22836 24664
rect 15804 24624 15810 24636
rect 14476 24568 15424 24596
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 18156 24596 18184 24636
rect 22830 24624 22836 24636
rect 22888 24624 22894 24676
rect 23109 24667 23167 24673
rect 23109 24633 23121 24667
rect 23155 24664 23167 24667
rect 24136 24664 24164 24704
rect 24854 24692 24860 24704
rect 24912 24692 24918 24744
rect 24964 24741 24992 24828
rect 25041 24803 25099 24809
rect 25041 24769 25053 24803
rect 25087 24800 25099 24803
rect 25406 24800 25412 24812
rect 25087 24772 25412 24800
rect 25087 24769 25099 24772
rect 25041 24763 25099 24769
rect 25406 24760 25412 24772
rect 25464 24760 25470 24812
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24800 25927 24803
rect 25915 24772 27476 24800
rect 25915 24769 25927 24772
rect 25869 24763 25927 24769
rect 24949 24735 25007 24741
rect 24949 24701 24961 24735
rect 24995 24701 25007 24735
rect 24949 24695 25007 24701
rect 23155 24636 24164 24664
rect 27448 24664 27476 24772
rect 27540 24732 27568 24840
rect 31386 24828 31392 24840
rect 31444 24828 31450 24880
rect 32674 24828 32680 24880
rect 32732 24828 32738 24880
rect 35710 24828 35716 24880
rect 35768 24868 35774 24880
rect 38948 24868 38976 24896
rect 35768 24840 36773 24868
rect 38948 24840 39896 24868
rect 35768 24828 35774 24840
rect 28350 24760 28356 24812
rect 28408 24800 28414 24812
rect 28445 24803 28503 24809
rect 28445 24800 28457 24803
rect 28408 24772 28457 24800
rect 28408 24760 28414 24772
rect 28445 24769 28457 24772
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 28629 24803 28687 24809
rect 28629 24769 28641 24803
rect 28675 24769 28687 24803
rect 28629 24763 28687 24769
rect 29089 24803 29147 24809
rect 29089 24769 29101 24803
rect 29135 24800 29147 24803
rect 29454 24800 29460 24812
rect 29135 24772 29460 24800
rect 29135 24769 29147 24772
rect 29089 24763 29147 24769
rect 28644 24732 28672 24763
rect 29454 24760 29460 24772
rect 29512 24760 29518 24812
rect 30098 24800 30104 24812
rect 29656 24772 30104 24800
rect 27540 24704 28672 24732
rect 27706 24664 27712 24676
rect 27448 24636 27712 24664
rect 23155 24633 23167 24636
rect 23109 24627 23167 24633
rect 15896 24568 18184 24596
rect 15896 24556 15902 24568
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 19521 24599 19579 24605
rect 19521 24596 19533 24599
rect 19392 24568 19533 24596
rect 19392 24556 19398 24568
rect 19521 24565 19533 24568
rect 19567 24565 19579 24599
rect 19521 24559 19579 24565
rect 22370 24556 22376 24608
rect 22428 24596 22434 24608
rect 23124 24596 23152 24627
rect 27706 24624 27712 24636
rect 27764 24624 27770 24676
rect 22428 24568 23152 24596
rect 22428 24556 22434 24568
rect 23842 24556 23848 24608
rect 23900 24596 23906 24608
rect 24121 24599 24179 24605
rect 24121 24596 24133 24599
rect 23900 24568 24133 24596
rect 23900 24556 23906 24568
rect 24121 24565 24133 24568
rect 24167 24565 24179 24599
rect 28460 24596 28488 24704
rect 29270 24692 29276 24744
rect 29328 24692 29334 24744
rect 29365 24735 29423 24741
rect 29365 24701 29377 24735
rect 29411 24732 29423 24735
rect 29656 24732 29684 24772
rect 30098 24760 30104 24772
rect 30156 24760 30162 24812
rect 30377 24803 30435 24809
rect 30377 24769 30389 24803
rect 30423 24800 30435 24803
rect 30558 24800 30564 24812
rect 30423 24772 30564 24800
rect 30423 24769 30435 24772
rect 30377 24763 30435 24769
rect 30558 24760 30564 24772
rect 30616 24760 30622 24812
rect 30742 24760 30748 24812
rect 30800 24760 30806 24812
rect 30834 24760 30840 24812
rect 30892 24809 30898 24812
rect 30892 24803 30915 24809
rect 30903 24769 30915 24803
rect 30892 24763 30915 24769
rect 30892 24760 30898 24763
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32493 24803 32551 24809
rect 32493 24800 32505 24803
rect 31812 24772 32505 24800
rect 31812 24760 31818 24772
rect 32493 24769 32505 24772
rect 32539 24769 32551 24803
rect 32493 24763 32551 24769
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 29411 24704 29684 24732
rect 29411 24701 29423 24704
rect 29365 24695 29423 24701
rect 29730 24692 29736 24744
rect 29788 24692 29794 24744
rect 30466 24692 30472 24744
rect 30524 24692 30530 24744
rect 32214 24692 32220 24744
rect 32272 24732 32278 24744
rect 32600 24732 32628 24763
rect 32858 24760 32864 24812
rect 32916 24760 32922 24812
rect 35986 24760 35992 24812
rect 36044 24800 36050 24812
rect 36745 24809 36773 24840
rect 36265 24803 36323 24809
rect 36265 24800 36277 24803
rect 36044 24772 36277 24800
rect 36044 24760 36050 24772
rect 36265 24769 36277 24772
rect 36311 24769 36323 24803
rect 36265 24763 36323 24769
rect 36358 24803 36416 24809
rect 36358 24769 36370 24803
rect 36404 24769 36416 24803
rect 36541 24803 36599 24809
rect 36541 24800 36553 24803
rect 36358 24763 36416 24769
rect 36464 24772 36553 24800
rect 32272 24704 32628 24732
rect 32272 24692 32278 24704
rect 28537 24667 28595 24673
rect 28537 24633 28549 24667
rect 28583 24664 28595 24667
rect 29748 24664 29776 24692
rect 28583 24636 29776 24664
rect 28583 24633 28595 24636
rect 28537 24627 28595 24633
rect 30650 24624 30656 24676
rect 30708 24664 30714 24676
rect 31570 24664 31576 24676
rect 30708 24636 31576 24664
rect 30708 24624 30714 24636
rect 31570 24624 31576 24636
rect 31628 24664 31634 24676
rect 36262 24664 36268 24676
rect 31628 24636 36268 24664
rect 31628 24624 31634 24636
rect 36262 24624 36268 24636
rect 36320 24664 36326 24676
rect 36372 24664 36400 24763
rect 36320 24636 36400 24664
rect 36320 24624 36326 24636
rect 30834 24596 30840 24608
rect 28460 24568 30840 24596
rect 24121 24559 24179 24565
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31018 24556 31024 24608
rect 31076 24556 31082 24608
rect 32309 24599 32367 24605
rect 32309 24565 32321 24599
rect 32355 24596 32367 24599
rect 32582 24596 32588 24608
rect 32355 24568 32588 24596
rect 32355 24565 32367 24568
rect 32309 24559 32367 24565
rect 32582 24556 32588 24568
rect 32640 24556 32646 24608
rect 35894 24556 35900 24608
rect 35952 24596 35958 24608
rect 36464 24596 36492 24772
rect 36541 24769 36553 24772
rect 36587 24769 36599 24803
rect 36541 24763 36599 24769
rect 36633 24803 36691 24809
rect 36633 24769 36645 24803
rect 36679 24769 36691 24803
rect 36633 24763 36691 24769
rect 36730 24803 36788 24809
rect 36730 24769 36742 24803
rect 36776 24769 36788 24803
rect 36730 24763 36788 24769
rect 36648 24732 36676 24763
rect 38562 24760 38568 24812
rect 38620 24760 38626 24812
rect 38713 24803 38771 24809
rect 38713 24769 38725 24803
rect 38759 24800 38771 24803
rect 38759 24769 38792 24800
rect 38713 24763 38792 24769
rect 38010 24732 38016 24744
rect 36648 24704 38016 24732
rect 38010 24692 38016 24704
rect 38068 24692 38074 24744
rect 35952 24568 36492 24596
rect 35952 24556 35958 24568
rect 36722 24556 36728 24608
rect 36780 24596 36786 24608
rect 36909 24599 36967 24605
rect 36909 24596 36921 24599
rect 36780 24568 36921 24596
rect 36780 24556 36786 24568
rect 36909 24565 36921 24568
rect 36955 24565 36967 24599
rect 36909 24559 36967 24565
rect 38654 24556 38660 24608
rect 38712 24596 38718 24608
rect 38764 24596 38792 24763
rect 38838 24760 38844 24812
rect 38896 24760 38902 24812
rect 38930 24760 38936 24812
rect 38988 24760 38994 24812
rect 39071 24803 39129 24809
rect 39071 24769 39083 24803
rect 39117 24800 39129 24803
rect 39390 24800 39396 24812
rect 39117 24772 39396 24800
rect 39117 24769 39129 24772
rect 39071 24763 39129 24769
rect 39390 24760 39396 24772
rect 39448 24760 39454 24812
rect 39482 24760 39488 24812
rect 39540 24800 39546 24812
rect 39868 24809 39896 24840
rect 39669 24803 39727 24809
rect 39669 24800 39681 24803
rect 39540 24772 39681 24800
rect 39540 24760 39546 24772
rect 39669 24769 39681 24772
rect 39715 24769 39727 24803
rect 39669 24763 39727 24769
rect 39853 24803 39911 24809
rect 39853 24769 39865 24803
rect 39899 24769 39911 24803
rect 39853 24763 39911 24769
rect 38856 24732 38884 24760
rect 39868 24732 39896 24763
rect 39942 24760 39948 24812
rect 40000 24800 40006 24812
rect 40126 24800 40132 24812
rect 40000 24772 40132 24800
rect 40000 24760 40006 24772
rect 40126 24760 40132 24772
rect 40184 24760 40190 24812
rect 40770 24760 40776 24812
rect 40828 24800 40834 24812
rect 41794 24803 41852 24809
rect 41794 24800 41806 24803
rect 40828 24772 41806 24800
rect 40828 24760 40834 24772
rect 41794 24769 41806 24772
rect 41840 24769 41852 24803
rect 41794 24763 41852 24769
rect 41966 24760 41972 24812
rect 42024 24800 42030 24812
rect 42061 24803 42119 24809
rect 42061 24800 42073 24803
rect 42024 24772 42073 24800
rect 42024 24760 42030 24772
rect 42061 24769 42073 24772
rect 42107 24769 42119 24803
rect 42061 24763 42119 24769
rect 42978 24760 42984 24812
rect 43036 24760 43042 24812
rect 38856 24704 39160 24732
rect 39868 24704 40448 24732
rect 39132 24676 39160 24704
rect 39114 24624 39120 24676
rect 39172 24624 39178 24676
rect 39669 24667 39727 24673
rect 39669 24633 39681 24667
rect 39715 24664 39727 24667
rect 40310 24664 40316 24676
rect 39715 24636 40316 24664
rect 39715 24633 39727 24636
rect 39669 24627 39727 24633
rect 40310 24624 40316 24636
rect 40368 24624 40374 24676
rect 39758 24596 39764 24608
rect 38712 24568 39764 24596
rect 38712 24556 38718 24568
rect 39758 24556 39764 24568
rect 39816 24556 39822 24608
rect 40420 24596 40448 24704
rect 43254 24692 43260 24744
rect 43312 24692 43318 24744
rect 40681 24599 40739 24605
rect 40681 24596 40693 24599
rect 40420 24568 40693 24596
rect 40681 24565 40693 24568
rect 40727 24565 40739 24599
rect 40681 24559 40739 24565
rect 42610 24556 42616 24608
rect 42668 24556 42674 24608
rect 1104 24506 43884 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 43884 24506
rect 1104 24432 43884 24454
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 9398 24392 9404 24404
rect 8352 24364 9404 24392
rect 8352 24352 8358 24364
rect 9398 24352 9404 24364
rect 9456 24392 9462 24404
rect 9456 24364 12434 24392
rect 9456 24352 9462 24364
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10321 24259 10379 24265
rect 10321 24256 10333 24259
rect 10192 24228 10333 24256
rect 10192 24216 10198 24228
rect 10321 24225 10333 24228
rect 10367 24225 10379 24259
rect 10321 24219 10379 24225
rect 10505 24259 10563 24265
rect 10505 24225 10517 24259
rect 10551 24256 10563 24259
rect 10870 24256 10876 24268
rect 10551 24228 10876 24256
rect 10551 24225 10563 24228
rect 10505 24219 10563 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 12406 24256 12434 24364
rect 14550 24352 14556 24404
rect 14608 24392 14614 24404
rect 14921 24395 14979 24401
rect 14921 24392 14933 24395
rect 14608 24364 14933 24392
rect 14608 24352 14614 24364
rect 14921 24361 14933 24364
rect 14967 24361 14979 24395
rect 22462 24392 22468 24404
rect 14921 24355 14979 24361
rect 15028 24364 22468 24392
rect 13906 24284 13912 24336
rect 13964 24324 13970 24336
rect 15028 24324 15056 24364
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 27246 24392 27252 24404
rect 22888 24364 27252 24392
rect 22888 24352 22894 24364
rect 27246 24352 27252 24364
rect 27304 24352 27310 24404
rect 28074 24352 28080 24404
rect 28132 24392 28138 24404
rect 28445 24395 28503 24401
rect 28445 24392 28457 24395
rect 28132 24364 28457 24392
rect 28132 24352 28138 24364
rect 28445 24361 28457 24364
rect 28491 24361 28503 24395
rect 28445 24355 28503 24361
rect 28813 24395 28871 24401
rect 28813 24361 28825 24395
rect 28859 24392 28871 24395
rect 30098 24392 30104 24404
rect 28859 24364 30104 24392
rect 28859 24361 28871 24364
rect 28813 24355 28871 24361
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 30469 24395 30527 24401
rect 30469 24361 30481 24395
rect 30515 24392 30527 24395
rect 30742 24392 30748 24404
rect 30515 24364 30748 24392
rect 30515 24361 30527 24364
rect 30469 24355 30527 24361
rect 30742 24352 30748 24364
rect 30800 24352 30806 24404
rect 38197 24395 38255 24401
rect 38197 24361 38209 24395
rect 38243 24392 38255 24395
rect 39206 24392 39212 24404
rect 38243 24364 39212 24392
rect 38243 24361 38255 24364
rect 38197 24355 38255 24361
rect 39206 24352 39212 24364
rect 39264 24352 39270 24404
rect 39482 24352 39488 24404
rect 39540 24352 39546 24404
rect 40770 24352 40776 24404
rect 40828 24352 40834 24404
rect 42978 24392 42984 24404
rect 41156 24364 42984 24392
rect 21082 24324 21088 24336
rect 13964 24296 15056 24324
rect 20088 24296 21088 24324
rect 13964 24284 13970 24296
rect 14645 24259 14703 24265
rect 14645 24256 14657 24259
rect 12406 24228 14657 24256
rect 14645 24225 14657 24228
rect 14691 24225 14703 24259
rect 14645 24219 14703 24225
rect 15378 24216 15384 24268
rect 15436 24256 15442 24268
rect 17313 24259 17371 24265
rect 17313 24256 17325 24259
rect 15436 24228 17325 24256
rect 15436 24216 15442 24228
rect 17313 24225 17325 24228
rect 17359 24225 17371 24259
rect 19978 24256 19984 24268
rect 17313 24219 17371 24225
rect 17972 24228 19984 24256
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11333 24191 11391 24197
rect 11333 24188 11345 24191
rect 11112 24160 11345 24188
rect 11112 24148 11118 24160
rect 11333 24157 11345 24160
rect 11379 24188 11391 24191
rect 11882 24188 11888 24200
rect 11379 24160 11888 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 14734 24148 14740 24200
rect 14792 24148 14798 24200
rect 16850 24148 16856 24200
rect 16908 24188 16914 24200
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16908 24160 17049 24188
rect 16908 24148 16914 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 11600 24123 11658 24129
rect 11600 24089 11612 24123
rect 11646 24120 11658 24123
rect 11698 24120 11704 24132
rect 11646 24092 11704 24120
rect 11646 24089 11658 24092
rect 11600 24083 11658 24089
rect 11698 24080 11704 24092
rect 11756 24080 11762 24132
rect 9858 24012 9864 24064
rect 9916 24012 9922 24064
rect 10226 24012 10232 24064
rect 10284 24012 10290 24064
rect 12710 24012 12716 24064
rect 12768 24052 12774 24064
rect 17972 24052 18000 24228
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20088 24197 20116 24296
rect 21082 24284 21088 24296
rect 21140 24284 21146 24336
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 23201 24327 23259 24333
rect 23201 24324 23213 24327
rect 22060 24296 23213 24324
rect 22060 24284 22066 24296
rect 23201 24293 23213 24296
rect 23247 24293 23259 24327
rect 23201 24287 23259 24293
rect 25314 24284 25320 24336
rect 25372 24324 25378 24336
rect 26881 24327 26939 24333
rect 26881 24324 26893 24327
rect 25372 24296 26893 24324
rect 25372 24284 25378 24296
rect 26881 24293 26893 24296
rect 26927 24293 26939 24327
rect 35802 24324 35808 24336
rect 26881 24287 26939 24293
rect 27172 24296 35808 24324
rect 20162 24216 20168 24268
rect 20220 24256 20226 24268
rect 23750 24256 23756 24268
rect 20220 24228 23756 24256
rect 20220 24216 20226 24228
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24188 20315 24191
rect 20530 24188 20536 24200
rect 20303 24160 20536 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 21729 24191 21787 24197
rect 21729 24157 21741 24191
rect 21775 24188 21787 24191
rect 22370 24188 22376 24200
rect 21775 24160 22376 24188
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24188 22707 24191
rect 22738 24188 22744 24200
rect 22695 24160 22744 24188
rect 22695 24157 22707 24160
rect 22649 24151 22707 24157
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 22848 24197 22876 24228
rect 23750 24216 23756 24228
rect 23808 24216 23814 24268
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 23474 24148 23480 24200
rect 23532 24148 23538 24200
rect 24578 24148 24584 24200
rect 24636 24148 24642 24200
rect 27062 24197 27068 24200
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 27060 24188 27068 24197
rect 27023 24160 27068 24188
rect 24765 24151 24823 24157
rect 27060 24151 27068 24160
rect 18693 24123 18751 24129
rect 18693 24089 18705 24123
rect 18739 24120 18751 24123
rect 24486 24120 24492 24132
rect 18739 24092 24492 24120
rect 18739 24089 18751 24092
rect 18693 24083 18751 24089
rect 24486 24080 24492 24092
rect 24544 24080 24550 24132
rect 24780 24120 24808 24151
rect 27062 24148 27068 24151
rect 27120 24148 27126 24200
rect 27172 24197 27200 24296
rect 35802 24284 35808 24296
rect 35860 24284 35866 24336
rect 38930 24284 38936 24336
rect 38988 24324 38994 24336
rect 41156 24324 41184 24364
rect 42978 24352 42984 24364
rect 43036 24392 43042 24404
rect 43349 24395 43407 24401
rect 43349 24392 43361 24395
rect 43036 24364 43361 24392
rect 43036 24352 43042 24364
rect 43349 24361 43361 24364
rect 43395 24361 43407 24395
rect 43349 24355 43407 24361
rect 38988 24296 41184 24324
rect 38988 24284 38994 24296
rect 27706 24216 27712 24268
rect 27764 24256 27770 24268
rect 29178 24256 29184 24268
rect 27764 24228 29184 24256
rect 27764 24216 27770 24228
rect 29178 24216 29184 24228
rect 29236 24216 29242 24268
rect 29730 24216 29736 24268
rect 29788 24256 29794 24268
rect 30285 24259 30343 24265
rect 30285 24256 30297 24259
rect 29788 24228 30297 24256
rect 29788 24216 29794 24228
rect 30285 24225 30297 24228
rect 30331 24225 30343 24259
rect 30285 24219 30343 24225
rect 31202 24216 31208 24268
rect 31260 24256 31266 24268
rect 34333 24259 34391 24265
rect 31260 24228 32904 24256
rect 31260 24216 31266 24228
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 27249 24191 27307 24197
rect 27249 24157 27261 24191
rect 27295 24188 27307 24191
rect 27338 24188 27344 24200
rect 27295 24160 27344 24188
rect 27295 24157 27307 24160
rect 27249 24151 27307 24157
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 27433 24191 27491 24197
rect 27433 24157 27445 24191
rect 27479 24188 27491 24191
rect 27522 24188 27528 24200
rect 27479 24160 27528 24188
rect 27479 24157 27491 24160
rect 27433 24151 27491 24157
rect 27522 24148 27528 24160
rect 27580 24188 27586 24200
rect 28258 24188 28264 24200
rect 27580 24160 28264 24188
rect 27580 24148 27586 24160
rect 28258 24148 28264 24160
rect 28316 24148 28322 24200
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 28534 24148 28540 24200
rect 28592 24188 28598 24200
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 28592 24160 28641 24188
rect 28592 24148 28598 24160
rect 28629 24157 28641 24160
rect 28675 24188 28687 24191
rect 28902 24188 28908 24200
rect 28675 24160 28908 24188
rect 28675 24157 28687 24160
rect 28629 24151 28687 24157
rect 28902 24148 28908 24160
rect 28960 24148 28966 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 24596 24092 24808 24120
rect 27356 24120 27384 24148
rect 27706 24120 27712 24132
rect 27356 24092 27712 24120
rect 12768 24024 18000 24052
rect 12768 24012 12774 24024
rect 19426 24012 19432 24064
rect 19484 24052 19490 24064
rect 20165 24055 20223 24061
rect 20165 24052 20177 24055
rect 19484 24024 20177 24052
rect 19484 24012 19490 24024
rect 20165 24021 20177 24024
rect 20211 24021 20223 24055
rect 20165 24015 20223 24021
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 21140 24024 21465 24052
rect 21140 24012 21146 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 24596 24052 24624 24092
rect 22520 24024 24624 24052
rect 22520 24012 22526 24024
rect 24670 24012 24676 24064
rect 24728 24012 24734 24064
rect 24780 24052 24808 24092
rect 27706 24080 27712 24092
rect 27764 24080 27770 24132
rect 28626 24052 28632 24064
rect 24780 24024 28632 24052
rect 28626 24012 28632 24024
rect 28684 24012 28690 24064
rect 30024 24052 30052 24151
rect 30098 24148 30104 24200
rect 30156 24148 30162 24200
rect 32876 24197 32904 24228
rect 34333 24225 34345 24259
rect 34379 24256 34391 24259
rect 34422 24256 34428 24268
rect 34379 24228 34428 24256
rect 34379 24225 34391 24228
rect 34333 24219 34391 24225
rect 34422 24216 34428 24228
rect 34480 24216 34486 24268
rect 37550 24216 37556 24268
rect 37608 24216 37614 24268
rect 37642 24216 37648 24268
rect 37700 24256 37706 24268
rect 38010 24256 38016 24268
rect 37700 24228 38016 24256
rect 37700 24216 37706 24228
rect 38010 24216 38016 24228
rect 38068 24216 38074 24268
rect 30193 24191 30251 24197
rect 30193 24157 30205 24191
rect 30239 24188 30251 24191
rect 31297 24191 31355 24197
rect 31297 24188 31309 24191
rect 30239 24160 31309 24188
rect 30239 24157 30251 24160
rect 30193 24151 30251 24157
rect 30300 24132 30328 24160
rect 31297 24157 31309 24160
rect 31343 24157 31355 24191
rect 31297 24151 31355 24157
rect 32861 24191 32919 24197
rect 32861 24157 32873 24191
rect 32907 24157 32919 24191
rect 32861 24151 32919 24157
rect 33042 24148 33048 24200
rect 33100 24188 33106 24200
rect 33229 24191 33287 24197
rect 33229 24188 33241 24191
rect 33100 24160 33241 24188
rect 33100 24148 33106 24160
rect 33229 24157 33241 24160
rect 33275 24157 33287 24191
rect 33229 24151 33287 24157
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 34241 24191 34299 24197
rect 34241 24157 34253 24191
rect 34287 24188 34299 24191
rect 35342 24188 35348 24200
rect 34287 24160 35348 24188
rect 34287 24157 34299 24160
rect 34241 24151 34299 24157
rect 30282 24080 30288 24132
rect 30340 24080 30346 24132
rect 30926 24080 30932 24132
rect 30984 24080 30990 24132
rect 31113 24123 31171 24129
rect 31113 24089 31125 24123
rect 31159 24120 31171 24123
rect 32950 24120 32956 24132
rect 31159 24092 32956 24120
rect 31159 24089 31171 24092
rect 31113 24083 31171 24089
rect 30466 24052 30472 24064
rect 30024 24024 30472 24052
rect 30466 24012 30472 24024
rect 30524 24012 30530 24064
rect 30834 24012 30840 24064
rect 30892 24052 30898 24064
rect 31128 24052 31156 24083
rect 32950 24080 32956 24092
rect 33008 24080 33014 24132
rect 33980 24120 34008 24151
rect 35342 24148 35348 24160
rect 35400 24148 35406 24200
rect 37826 24148 37832 24200
rect 37884 24188 37890 24200
rect 37921 24191 37979 24197
rect 37921 24188 37933 24191
rect 37884 24160 37933 24188
rect 37884 24148 37890 24160
rect 37921 24157 37933 24160
rect 37967 24157 37979 24191
rect 37921 24151 37979 24157
rect 38838 24148 38844 24200
rect 38896 24148 38902 24200
rect 38948 24197 38976 24284
rect 40310 24216 40316 24268
rect 40368 24216 40374 24268
rect 41966 24216 41972 24268
rect 42024 24216 42030 24268
rect 38934 24191 38992 24197
rect 38934 24157 38946 24191
rect 38980 24157 38992 24191
rect 38934 24151 38992 24157
rect 39022 24148 39028 24200
rect 39080 24197 39086 24200
rect 39080 24191 39129 24197
rect 39080 24157 39083 24191
rect 39117 24157 39129 24191
rect 39080 24151 39129 24157
rect 39347 24191 39405 24197
rect 39347 24157 39359 24191
rect 39393 24188 39405 24191
rect 39574 24188 39580 24200
rect 39393 24160 39580 24188
rect 39393 24157 39405 24160
rect 39347 24151 39405 24157
rect 39080 24148 39086 24151
rect 39574 24148 39580 24160
rect 39632 24148 39638 24200
rect 40402 24148 40408 24200
rect 40460 24148 40466 24200
rect 42236 24191 42294 24197
rect 42236 24157 42248 24191
rect 42282 24188 42294 24191
rect 42610 24188 42616 24200
rect 42282 24160 42616 24188
rect 42282 24157 42294 24160
rect 42236 24151 42294 24157
rect 42610 24148 42616 24160
rect 42668 24148 42674 24200
rect 34606 24120 34612 24132
rect 33980 24092 34612 24120
rect 34606 24080 34612 24092
rect 34664 24080 34670 24132
rect 35526 24080 35532 24132
rect 35584 24120 35590 24132
rect 37645 24123 37703 24129
rect 37645 24120 37657 24123
rect 35584 24092 37657 24120
rect 35584 24080 35590 24092
rect 37645 24089 37657 24092
rect 37691 24120 37703 24123
rect 37691 24092 38976 24120
rect 37691 24089 37703 24092
rect 37645 24083 37703 24089
rect 38948 24064 38976 24092
rect 39206 24080 39212 24132
rect 39264 24080 39270 24132
rect 30892 24024 31156 24052
rect 30892 24012 30898 24024
rect 35250 24012 35256 24064
rect 35308 24052 35314 24064
rect 38654 24052 38660 24064
rect 35308 24024 38660 24052
rect 35308 24012 35314 24024
rect 38654 24012 38660 24024
rect 38712 24012 38718 24064
rect 38930 24012 38936 24064
rect 38988 24012 38994 24064
rect 1104 23962 43884 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 43884 23962
rect 1104 23888 43884 23910
rect 14734 23808 14740 23860
rect 14792 23848 14798 23860
rect 14792 23820 15884 23848
rect 14792 23808 14798 23820
rect 11054 23780 11060 23792
rect 9232 23752 11060 23780
rect 9232 23721 9260 23752
rect 11054 23740 11060 23752
rect 11112 23740 11118 23792
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9484 23715 9542 23721
rect 9484 23681 9496 23715
rect 9530 23712 9542 23715
rect 9858 23712 9864 23724
rect 9530 23684 9864 23712
rect 9530 23681 9542 23684
rect 9484 23675 9542 23681
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 15028 23721 15056 23820
rect 15856 23721 15884 23820
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20312 23820 23796 23848
rect 20312 23808 20318 23820
rect 21177 23783 21235 23789
rect 21177 23780 21189 23783
rect 20824 23752 21189 23780
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23712 15255 23715
rect 15749 23715 15807 23721
rect 15749 23712 15761 23715
rect 15243 23684 15761 23712
rect 15243 23681 15255 23684
rect 15197 23675 15255 23681
rect 15749 23681 15761 23684
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23712 15899 23715
rect 15887 23684 17080 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 10226 23604 10232 23656
rect 10284 23644 10290 23656
rect 15212 23644 15240 23675
rect 10284 23616 15240 23644
rect 15289 23647 15347 23653
rect 10284 23604 10290 23616
rect 10612 23585 10640 23616
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 16206 23644 16212 23656
rect 15335 23616 16212 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 16301 23647 16359 23653
rect 16301 23613 16313 23647
rect 16347 23644 16359 23647
rect 16942 23644 16948 23656
rect 16347 23616 16948 23644
rect 16347 23613 16359 23616
rect 16301 23607 16359 23613
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17052 23644 17080 23684
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19889 23715 19947 23721
rect 19889 23712 19901 23715
rect 19484 23684 19901 23712
rect 19484 23672 19490 23684
rect 19889 23681 19901 23684
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 19981 23715 20039 23721
rect 19981 23681 19993 23715
rect 20027 23681 20039 23715
rect 19981 23675 20039 23681
rect 20073 23715 20131 23721
rect 20073 23681 20085 23715
rect 20119 23681 20131 23715
rect 20073 23675 20131 23681
rect 17052 23616 19748 23644
rect 10597 23579 10655 23585
rect 10597 23545 10609 23579
rect 10643 23545 10655 23579
rect 10597 23539 10655 23545
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 18104 23480 19625 23508
rect 18104 23468 18110 23480
rect 19613 23477 19625 23480
rect 19659 23477 19671 23511
rect 19720 23508 19748 23616
rect 19996 23576 20024 23675
rect 20088 23644 20116 23675
rect 20254 23672 20260 23724
rect 20312 23672 20318 23724
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 20824 23712 20852 23752
rect 21177 23749 21189 23752
rect 21223 23780 21235 23783
rect 22002 23780 22008 23792
rect 21223 23752 22008 23780
rect 21223 23749 21235 23752
rect 21177 23743 21235 23749
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 22462 23740 22468 23792
rect 22520 23740 22526 23792
rect 23768 23780 23796 23820
rect 24394 23808 24400 23860
rect 24452 23808 24458 23860
rect 24489 23851 24547 23857
rect 24489 23817 24501 23851
rect 24535 23848 24547 23851
rect 24578 23848 24584 23860
rect 24535 23820 24584 23848
rect 24535 23817 24547 23820
rect 24489 23811 24547 23817
rect 24504 23780 24532 23811
rect 24578 23808 24584 23820
rect 24636 23808 24642 23860
rect 26970 23808 26976 23860
rect 27028 23848 27034 23860
rect 27357 23851 27415 23857
rect 27357 23848 27369 23851
rect 27028 23820 27369 23848
rect 27028 23808 27034 23820
rect 27357 23817 27369 23820
rect 27403 23817 27415 23851
rect 27357 23811 27415 23817
rect 28074 23808 28080 23860
rect 28132 23808 28138 23860
rect 28258 23808 28264 23860
rect 28316 23848 28322 23860
rect 31202 23848 31208 23860
rect 28316 23820 31208 23848
rect 28316 23808 28322 23820
rect 31202 23808 31208 23820
rect 31260 23808 31266 23860
rect 31665 23851 31723 23857
rect 31665 23817 31677 23851
rect 31711 23848 31723 23851
rect 33134 23848 33140 23860
rect 31711 23820 33140 23848
rect 31711 23817 31723 23820
rect 31665 23811 31723 23817
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 39942 23848 39948 23860
rect 35176 23820 39948 23848
rect 23768 23752 24532 23780
rect 24670 23740 24676 23792
rect 24728 23740 24734 23792
rect 25590 23740 25596 23792
rect 25648 23740 25654 23792
rect 26694 23740 26700 23792
rect 26752 23780 26758 23792
rect 27154 23780 27160 23792
rect 26752 23752 27160 23780
rect 26752 23740 26758 23752
rect 27154 23740 27160 23752
rect 27212 23740 27218 23792
rect 35176 23789 35204 23820
rect 39942 23808 39948 23820
rect 40000 23808 40006 23860
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 27448 23752 32965 23780
rect 20588 23684 20852 23712
rect 20588 23672 20594 23684
rect 21082 23672 21088 23724
rect 21140 23672 21146 23724
rect 21542 23672 21548 23724
rect 21600 23712 21606 23724
rect 21600 23684 23428 23712
rect 21600 23672 21606 23684
rect 20990 23644 20996 23656
rect 20088 23616 20996 23644
rect 20990 23604 20996 23616
rect 21048 23604 21054 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23644 21419 23647
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21407 23616 22017 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 23400 23644 23428 23684
rect 23474 23672 23480 23724
rect 23532 23672 23538 23724
rect 24302 23672 24308 23724
rect 24360 23672 24366 23724
rect 27448 23712 27476 23752
rect 32953 23749 32965 23752
rect 32999 23749 33011 23783
rect 32953 23743 33011 23749
rect 35161 23783 35219 23789
rect 35161 23749 35173 23783
rect 35207 23749 35219 23783
rect 35161 23743 35219 23749
rect 35986 23740 35992 23792
rect 36044 23780 36050 23792
rect 36044 23752 36768 23780
rect 36044 23740 36050 23752
rect 24412 23684 27476 23712
rect 27985 23715 28043 23721
rect 24412 23644 24440 23684
rect 27985 23681 27997 23715
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 23400 23616 24440 23644
rect 22005 23607 22063 23613
rect 27154 23604 27160 23656
rect 27212 23644 27218 23656
rect 28000 23644 28028 23675
rect 28166 23672 28172 23724
rect 28224 23672 28230 23724
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23681 28871 23715
rect 28813 23675 28871 23681
rect 27212 23616 28028 23644
rect 27212 23604 27218 23616
rect 28074 23604 28080 23656
rect 28132 23644 28138 23656
rect 28828 23644 28856 23675
rect 28902 23672 28908 23724
rect 28960 23672 28966 23724
rect 29178 23672 29184 23724
rect 29236 23712 29242 23724
rect 30009 23715 30067 23721
rect 30009 23712 30021 23715
rect 29236 23684 30021 23712
rect 29236 23672 29242 23684
rect 30009 23681 30021 23684
rect 30055 23681 30067 23715
rect 30009 23675 30067 23681
rect 30377 23715 30435 23721
rect 30377 23681 30389 23715
rect 30423 23712 30435 23715
rect 30466 23712 30472 23724
rect 30423 23684 30472 23712
rect 30423 23681 30435 23684
rect 30377 23675 30435 23681
rect 30466 23672 30472 23684
rect 30524 23672 30530 23724
rect 30558 23672 30564 23724
rect 30616 23712 30622 23724
rect 31515 23715 31573 23721
rect 31515 23712 31527 23715
rect 30616 23684 31527 23712
rect 30616 23672 30622 23684
rect 31515 23681 31527 23684
rect 31561 23681 31573 23715
rect 31515 23675 31573 23681
rect 32582 23672 32588 23724
rect 32640 23672 32646 23724
rect 32678 23715 32736 23721
rect 32678 23681 32690 23715
rect 32724 23681 32736 23715
rect 32678 23675 32736 23681
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 32861 23675 32919 23681
rect 33091 23715 33149 23721
rect 33091 23681 33103 23715
rect 33137 23712 33149 23715
rect 33686 23712 33692 23724
rect 33137 23684 33692 23712
rect 33137 23681 33149 23684
rect 33091 23675 33149 23681
rect 31113 23647 31171 23653
rect 28132 23616 28856 23644
rect 28966 23616 31064 23644
rect 28132 23604 28138 23616
rect 20717 23579 20775 23585
rect 20717 23576 20729 23579
rect 19996 23548 20729 23576
rect 20717 23545 20729 23548
rect 20763 23545 20775 23579
rect 20717 23539 20775 23545
rect 21174 23536 21180 23588
rect 21232 23576 21238 23588
rect 22186 23576 22192 23588
rect 21232 23548 22192 23576
rect 21232 23536 21238 23548
rect 22186 23536 22192 23548
rect 22244 23536 22250 23588
rect 24118 23536 24124 23588
rect 24176 23536 24182 23588
rect 25314 23536 25320 23588
rect 25372 23536 25378 23588
rect 25406 23536 25412 23588
rect 25464 23576 25470 23588
rect 28966 23576 28994 23616
rect 25464 23548 28994 23576
rect 25464 23536 25470 23548
rect 29178 23536 29184 23588
rect 29236 23536 29242 23588
rect 29288 23548 30236 23576
rect 22738 23508 22744 23520
rect 19720 23480 22744 23508
rect 19613 23471 19671 23477
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 23569 23511 23627 23517
rect 23569 23477 23581 23511
rect 23615 23508 23627 23511
rect 25038 23508 25044 23520
rect 23615 23480 25044 23508
rect 23615 23477 23627 23480
rect 23569 23471 23627 23477
rect 25038 23468 25044 23480
rect 25096 23468 25102 23520
rect 25130 23468 25136 23520
rect 25188 23468 25194 23520
rect 27246 23468 27252 23520
rect 27304 23508 27310 23520
rect 27341 23511 27399 23517
rect 27341 23508 27353 23511
rect 27304 23480 27353 23508
rect 27304 23468 27310 23480
rect 27341 23477 27353 23480
rect 27387 23477 27399 23511
rect 27341 23471 27399 23477
rect 27525 23511 27583 23517
rect 27525 23477 27537 23511
rect 27571 23508 27583 23511
rect 28350 23508 28356 23520
rect 27571 23480 28356 23508
rect 27571 23477 27583 23480
rect 27525 23471 27583 23477
rect 28350 23468 28356 23480
rect 28408 23508 28414 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28408 23480 28917 23508
rect 28408 23468 28414 23480
rect 28905 23477 28917 23480
rect 28951 23508 28963 23511
rect 29288 23508 29316 23548
rect 28951 23480 29316 23508
rect 28951 23477 28963 23480
rect 28905 23471 28963 23477
rect 30098 23468 30104 23520
rect 30156 23468 30162 23520
rect 30208 23508 30236 23548
rect 30558 23536 30564 23588
rect 30616 23536 30622 23588
rect 30926 23508 30932 23520
rect 30208 23480 30932 23508
rect 30926 23468 30932 23480
rect 30984 23468 30990 23520
rect 31036 23508 31064 23616
rect 31113 23613 31125 23647
rect 31159 23613 31171 23647
rect 31113 23607 31171 23613
rect 31128 23576 31156 23607
rect 31202 23604 31208 23656
rect 31260 23644 31266 23656
rect 31260 23616 31754 23644
rect 31260 23604 31266 23616
rect 31294 23576 31300 23588
rect 31128 23548 31300 23576
rect 31294 23536 31300 23548
rect 31352 23536 31358 23588
rect 31726 23576 31754 23616
rect 32030 23604 32036 23656
rect 32088 23644 32094 23656
rect 32692 23644 32720 23675
rect 32088 23616 32720 23644
rect 32876 23644 32904 23675
rect 33686 23672 33692 23684
rect 33744 23712 33750 23724
rect 33962 23712 33968 23724
rect 33744 23684 33968 23712
rect 33744 23672 33750 23684
rect 33962 23672 33968 23684
rect 34020 23672 34026 23724
rect 34054 23672 34060 23724
rect 34112 23672 34118 23724
rect 34606 23672 34612 23724
rect 34664 23672 34670 23724
rect 34977 23715 35035 23721
rect 34977 23681 34989 23715
rect 35023 23712 35035 23715
rect 35342 23712 35348 23724
rect 35023 23684 35348 23712
rect 35023 23681 35035 23684
rect 34977 23675 35035 23681
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 35526 23672 35532 23724
rect 35584 23712 35590 23724
rect 36446 23712 36452 23724
rect 35584 23684 36452 23712
rect 35584 23672 35590 23684
rect 36446 23672 36452 23684
rect 36504 23712 36510 23724
rect 36740 23721 36768 23752
rect 36541 23715 36599 23721
rect 36541 23712 36553 23715
rect 36504 23684 36553 23712
rect 36504 23672 36510 23684
rect 36541 23681 36553 23684
rect 36587 23681 36599 23715
rect 36541 23675 36599 23681
rect 36725 23715 36783 23721
rect 36725 23681 36737 23715
rect 36771 23712 36783 23715
rect 37182 23712 37188 23724
rect 36771 23684 37188 23712
rect 36771 23681 36783 23684
rect 36725 23675 36783 23681
rect 37182 23672 37188 23684
rect 37240 23672 37246 23724
rect 42702 23672 42708 23724
rect 42760 23712 42766 23724
rect 42889 23715 42947 23721
rect 42889 23712 42901 23715
rect 42760 23684 42901 23712
rect 42760 23672 42766 23684
rect 42889 23681 42901 23684
rect 42935 23681 42947 23715
rect 42889 23675 42947 23681
rect 35894 23644 35900 23656
rect 32876 23616 35900 23644
rect 32088 23604 32094 23616
rect 35360 23588 35388 23616
rect 35894 23604 35900 23616
rect 35952 23604 35958 23656
rect 39022 23604 39028 23656
rect 39080 23644 39086 23656
rect 39206 23644 39212 23656
rect 39080 23616 39212 23644
rect 39080 23604 39086 23616
rect 39206 23604 39212 23616
rect 39264 23604 39270 23656
rect 43165 23647 43223 23653
rect 43165 23613 43177 23647
rect 43211 23644 43223 23647
rect 43990 23644 43996 23656
rect 43211 23616 43996 23644
rect 43211 23613 43223 23616
rect 43165 23607 43223 23613
rect 43990 23604 43996 23616
rect 44048 23604 44054 23656
rect 35250 23576 35256 23588
rect 31726 23548 35256 23576
rect 35250 23536 35256 23548
rect 35308 23536 35314 23588
rect 35342 23536 35348 23588
rect 35400 23536 35406 23588
rect 39574 23576 39580 23588
rect 35452 23548 39580 23576
rect 33042 23508 33048 23520
rect 31036 23480 33048 23508
rect 33042 23468 33048 23480
rect 33100 23468 33106 23520
rect 33229 23511 33287 23517
rect 33229 23477 33241 23511
rect 33275 23508 33287 23511
rect 33502 23508 33508 23520
rect 33275 23480 33508 23508
rect 33275 23477 33287 23480
rect 33229 23471 33287 23477
rect 33502 23468 33508 23480
rect 33560 23468 33566 23520
rect 34054 23468 34060 23520
rect 34112 23508 34118 23520
rect 34606 23508 34612 23520
rect 34112 23480 34612 23508
rect 34112 23468 34118 23480
rect 34606 23468 34612 23480
rect 34664 23508 34670 23520
rect 35452 23508 35480 23548
rect 39574 23536 39580 23548
rect 39632 23536 39638 23588
rect 34664 23480 35480 23508
rect 36633 23511 36691 23517
rect 34664 23468 34670 23480
rect 36633 23477 36645 23511
rect 36679 23508 36691 23511
rect 37642 23508 37648 23520
rect 36679 23480 37648 23508
rect 36679 23477 36691 23480
rect 36633 23471 36691 23477
rect 37642 23468 37648 23480
rect 37700 23468 37706 23520
rect 1104 23418 43884 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 43884 23418
rect 1104 23344 43884 23366
rect 10962 23304 10968 23316
rect 10704 23276 10968 23304
rect 10704 23180 10732 23276
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 17310 23264 17316 23316
rect 17368 23264 17374 23316
rect 22462 23304 22468 23316
rect 18524 23276 22468 23304
rect 10686 23128 10692 23180
rect 10744 23128 10750 23180
rect 15749 23171 15807 23177
rect 15749 23137 15761 23171
rect 15795 23168 15807 23171
rect 16850 23168 16856 23180
rect 15795 23140 16856 23168
rect 15795 23137 15807 23140
rect 15749 23131 15807 23137
rect 16850 23128 16856 23140
rect 16908 23128 16914 23180
rect 16022 23060 16028 23112
rect 16080 23060 16086 23112
rect 10956 23035 11014 23041
rect 10956 23001 10968 23035
rect 11002 23032 11014 23035
rect 12250 23032 12256 23044
rect 11002 23004 12256 23032
rect 11002 23001 11014 23004
rect 10956 22995 11014 23001
rect 12250 22992 12256 23004
rect 12308 22992 12314 23044
rect 16758 22992 16764 23044
rect 16816 23032 16822 23044
rect 18524 23032 18552 23276
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 24302 23264 24308 23316
rect 24360 23304 24366 23316
rect 24581 23307 24639 23313
rect 24581 23304 24593 23307
rect 24360 23276 24593 23304
rect 24360 23264 24366 23276
rect 24581 23273 24593 23276
rect 24627 23273 24639 23307
rect 24581 23267 24639 23273
rect 24762 23264 24768 23316
rect 24820 23304 24826 23316
rect 24820 23276 28994 23304
rect 24820 23264 24826 23276
rect 18782 23196 18788 23248
rect 18840 23236 18846 23248
rect 18877 23239 18935 23245
rect 18877 23236 18889 23239
rect 18840 23208 18889 23236
rect 18840 23196 18846 23208
rect 18877 23205 18889 23208
rect 18923 23205 18935 23239
rect 23385 23239 23443 23245
rect 23385 23236 23397 23239
rect 18877 23199 18935 23205
rect 19812 23208 21404 23236
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 18690 23100 18696 23112
rect 18647 23072 18696 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 18690 23060 18696 23072
rect 18748 23100 18754 23112
rect 19812 23100 19840 23208
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23168 20039 23171
rect 20438 23168 20444 23180
rect 20027 23140 20444 23168
rect 20027 23137 20039 23140
rect 19981 23131 20039 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 20990 23128 20996 23180
rect 21048 23128 21054 23180
rect 18748 23072 19840 23100
rect 18748 23060 18754 23072
rect 19886 23060 19892 23112
rect 19944 23100 19950 23112
rect 20073 23103 20131 23109
rect 20073 23100 20085 23103
rect 19944 23072 20085 23100
rect 19944 23060 19950 23072
rect 20073 23069 20085 23072
rect 20119 23100 20131 23103
rect 21082 23100 21088 23112
rect 20119 23072 21088 23100
rect 20119 23069 20131 23072
rect 20073 23063 20131 23069
rect 21082 23060 21088 23072
rect 21140 23060 21146 23112
rect 21174 23060 21180 23112
rect 21232 23060 21238 23112
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23069 21327 23103
rect 21376 23100 21404 23208
rect 23124 23208 23397 23236
rect 22373 23171 22431 23177
rect 22373 23137 22385 23171
rect 22419 23168 22431 23171
rect 23124 23168 23152 23208
rect 23385 23205 23397 23208
rect 23431 23236 23443 23239
rect 26602 23236 26608 23248
rect 23431 23208 26608 23236
rect 23431 23205 23443 23208
rect 23385 23199 23443 23205
rect 26602 23196 26608 23208
rect 26660 23196 26666 23248
rect 22419 23140 23152 23168
rect 22419 23137 22431 23140
rect 22373 23131 22431 23137
rect 22388 23100 22416 23131
rect 23198 23128 23204 23180
rect 23256 23128 23262 23180
rect 25038 23128 25044 23180
rect 25096 23128 25102 23180
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 26970 23128 26976 23180
rect 27028 23168 27034 23180
rect 27430 23168 27436 23180
rect 27028 23140 27436 23168
rect 27028 23128 27034 23140
rect 27430 23128 27436 23140
rect 27488 23128 27494 23180
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23168 27583 23171
rect 28166 23168 28172 23180
rect 27571 23140 28172 23168
rect 27571 23137 27583 23140
rect 27525 23131 27583 23137
rect 28166 23128 28172 23140
rect 28224 23128 28230 23180
rect 28966 23168 28994 23276
rect 30282 23264 30288 23316
rect 30340 23304 30346 23316
rect 31754 23304 31760 23316
rect 30340 23276 31760 23304
rect 30340 23264 30346 23276
rect 31754 23264 31760 23276
rect 31812 23304 31818 23316
rect 32490 23304 32496 23316
rect 31812 23276 32496 23304
rect 31812 23264 31818 23276
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 33042 23264 33048 23316
rect 33100 23304 33106 23316
rect 38194 23304 38200 23316
rect 33100 23276 38200 23304
rect 33100 23264 33106 23276
rect 38194 23264 38200 23276
rect 38252 23264 38258 23316
rect 43070 23304 43076 23316
rect 39408 23276 43076 23304
rect 30098 23196 30104 23248
rect 30156 23236 30162 23248
rect 34057 23239 34115 23245
rect 30156 23208 34008 23236
rect 30156 23196 30162 23208
rect 33980 23168 34008 23208
rect 34057 23205 34069 23239
rect 34103 23236 34115 23239
rect 37737 23239 37795 23245
rect 34103 23208 36860 23236
rect 34103 23205 34115 23208
rect 34057 23199 34115 23205
rect 35526 23168 35532 23180
rect 28966 23140 31754 23168
rect 33980 23140 35532 23168
rect 21376 23072 22416 23100
rect 21269 23063 21327 23069
rect 18877 23035 18935 23041
rect 18877 23032 18889 23035
rect 16816 23004 18889 23032
rect 16816 22992 16822 23004
rect 18877 23001 18889 23004
rect 18923 23001 18935 23035
rect 18877 22995 18935 23001
rect 19242 22992 19248 23044
rect 19300 23032 19306 23044
rect 21192 23032 21220 23060
rect 19300 23004 21220 23032
rect 19300 22992 19306 23004
rect 12066 22924 12072 22976
rect 12124 22924 12130 22976
rect 18693 22967 18751 22973
rect 18693 22933 18705 22967
rect 18739 22964 18751 22967
rect 19702 22964 19708 22976
rect 18739 22936 19708 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 19702 22924 19708 22936
rect 19760 22924 19766 22976
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22964 19855 22967
rect 19978 22964 19984 22976
rect 19843 22936 19984 22964
rect 19843 22933 19855 22936
rect 19797 22927 19855 22933
rect 19978 22924 19984 22936
rect 20036 22924 20042 22976
rect 20346 22924 20352 22976
rect 20404 22964 20410 22976
rect 20441 22967 20499 22973
rect 20441 22964 20453 22967
rect 20404 22936 20453 22964
rect 20404 22924 20410 22936
rect 20441 22933 20453 22936
rect 20487 22933 20499 22967
rect 20441 22927 20499 22933
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21284 22964 21312 23063
rect 22462 23060 22468 23112
rect 22520 23060 22526 23112
rect 22554 23060 22560 23112
rect 22612 23060 22618 23112
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23069 22707 23103
rect 22649 23063 22707 23069
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23100 23535 23103
rect 24762 23100 24768 23112
rect 23523 23072 24768 23100
rect 23523 23069 23535 23072
rect 23477 23063 23535 23069
rect 21637 23035 21695 23041
rect 21637 23001 21649 23035
rect 21683 23032 21695 23035
rect 22370 23032 22376 23044
rect 21683 23004 22376 23032
rect 21683 23001 21695 23004
rect 21637 22995 21695 23001
rect 22370 22992 22376 23004
rect 22428 22992 22434 23044
rect 22664 23032 22692 23063
rect 24762 23060 24768 23072
rect 24820 23100 24826 23112
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 24820 23072 24961 23100
rect 24820 23060 24826 23072
rect 24949 23069 24961 23072
rect 24995 23100 25007 23103
rect 26145 23103 26203 23109
rect 26145 23100 26157 23103
rect 24995 23072 26157 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 26145 23069 26157 23072
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 27157 23103 27215 23109
rect 27157 23069 27169 23103
rect 27203 23100 27215 23103
rect 27246 23100 27252 23112
rect 27203 23072 27252 23100
rect 27203 23069 27215 23072
rect 27157 23063 27215 23069
rect 27246 23060 27252 23072
rect 27304 23060 27310 23112
rect 30282 23060 30288 23112
rect 30340 23102 30346 23112
rect 30340 23074 30383 23102
rect 31726 23100 31754 23140
rect 35526 23128 35532 23140
rect 35584 23128 35590 23180
rect 36078 23168 36084 23180
rect 35728 23140 36084 23168
rect 33505 23103 33563 23109
rect 33505 23100 33517 23103
rect 30340 23060 30346 23074
rect 31726 23072 33517 23100
rect 33505 23069 33517 23072
rect 33551 23069 33563 23103
rect 33505 23063 33563 23069
rect 33686 23060 33692 23112
rect 33744 23060 33750 23112
rect 33873 23103 33931 23109
rect 33873 23069 33885 23103
rect 33919 23100 33931 23103
rect 34238 23100 34244 23112
rect 33919 23072 34244 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 34238 23060 34244 23072
rect 34296 23060 34302 23112
rect 35618 23060 35624 23112
rect 35676 23060 35682 23112
rect 35728 23109 35756 23140
rect 36078 23128 36084 23140
rect 36136 23128 36142 23180
rect 36538 23128 36544 23180
rect 36596 23128 36602 23180
rect 35713 23103 35771 23109
rect 35713 23069 35725 23103
rect 35759 23069 35771 23103
rect 35713 23063 35771 23069
rect 35802 23060 35808 23112
rect 35860 23060 35866 23112
rect 35897 23103 35955 23109
rect 35897 23069 35909 23103
rect 35943 23100 35955 23103
rect 36170 23100 36176 23112
rect 35943 23072 36176 23100
rect 35943 23069 35955 23072
rect 35897 23063 35955 23069
rect 36170 23060 36176 23072
rect 36228 23060 36234 23112
rect 36449 23103 36507 23109
rect 36449 23069 36461 23103
rect 36495 23100 36507 23103
rect 36630 23100 36636 23112
rect 36495 23072 36636 23100
rect 36495 23069 36507 23072
rect 36449 23063 36507 23069
rect 36630 23060 36636 23072
rect 36688 23060 36694 23112
rect 36722 23060 36728 23112
rect 36780 23060 36786 23112
rect 36832 23109 36860 23208
rect 37737 23205 37749 23239
rect 37783 23236 37795 23239
rect 38470 23236 38476 23248
rect 37783 23208 38476 23236
rect 37783 23205 37795 23208
rect 37737 23199 37795 23205
rect 38470 23196 38476 23208
rect 38528 23196 38534 23248
rect 37182 23128 37188 23180
rect 37240 23168 37246 23180
rect 38105 23171 38163 23177
rect 37240 23140 37964 23168
rect 37240 23128 37246 23140
rect 36817 23103 36875 23109
rect 36817 23069 36829 23103
rect 36863 23069 36875 23103
rect 36817 23063 36875 23069
rect 37642 23060 37648 23112
rect 37700 23060 37706 23112
rect 37936 23109 37964 23140
rect 38105 23137 38117 23171
rect 38151 23168 38163 23171
rect 39408 23168 39436 23276
rect 43070 23264 43076 23276
rect 43128 23264 43134 23316
rect 39485 23239 39543 23245
rect 39485 23205 39497 23239
rect 39531 23236 39543 23239
rect 39531 23208 40448 23236
rect 39531 23205 39543 23208
rect 39485 23199 39543 23205
rect 38151 23140 39436 23168
rect 40129 23171 40187 23177
rect 38151 23137 38163 23140
rect 38105 23131 38163 23137
rect 40129 23137 40141 23171
rect 40175 23168 40187 23171
rect 40218 23168 40224 23180
rect 40175 23140 40224 23168
rect 40175 23137 40187 23140
rect 40129 23131 40187 23137
rect 40218 23128 40224 23140
rect 40276 23128 40282 23180
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23069 37887 23103
rect 37829 23063 37887 23069
rect 37921 23103 37979 23109
rect 37921 23069 37933 23103
rect 37967 23069 37979 23103
rect 37921 23063 37979 23069
rect 23201 23035 23259 23041
rect 23201 23032 23213 23035
rect 22664 23004 23213 23032
rect 23201 23001 23213 23004
rect 23247 23001 23259 23035
rect 23201 22995 23259 23001
rect 25774 22992 25780 23044
rect 25832 22992 25838 23044
rect 25961 23035 26019 23041
rect 25961 23001 25973 23035
rect 26007 23001 26019 23035
rect 27264 23032 27292 23060
rect 28350 23032 28356 23044
rect 27264 23004 28356 23032
rect 25961 22995 26019 23001
rect 21232 22936 21312 22964
rect 21232 22924 21238 22936
rect 22186 22924 22192 22976
rect 22244 22924 22250 22976
rect 24854 22924 24860 22976
rect 24912 22964 24918 22976
rect 25498 22964 25504 22976
rect 24912 22936 25504 22964
rect 24912 22924 24918 22936
rect 25498 22924 25504 22936
rect 25556 22964 25562 22976
rect 25976 22964 26004 22995
rect 28350 22992 28356 23004
rect 28408 22992 28414 23044
rect 33781 23035 33839 23041
rect 33781 23001 33793 23035
rect 33827 23001 33839 23035
rect 33781 22995 33839 23001
rect 25556 22936 26004 22964
rect 30377 22967 30435 22973
rect 25556 22924 25562 22936
rect 30377 22933 30389 22967
rect 30423 22964 30435 22967
rect 30834 22964 30840 22976
rect 30423 22936 30840 22964
rect 30423 22933 30435 22936
rect 30377 22927 30435 22933
rect 30834 22924 30840 22936
rect 30892 22924 30898 22976
rect 33318 22924 33324 22976
rect 33376 22964 33382 22976
rect 33796 22964 33824 22995
rect 34146 22992 34152 23044
rect 34204 23032 34210 23044
rect 37844 23032 37872 23063
rect 38746 23060 38752 23112
rect 38804 23100 38810 23112
rect 39022 23109 39028 23112
rect 38841 23103 38899 23109
rect 38841 23100 38853 23103
rect 38804 23072 38853 23100
rect 38804 23060 38810 23072
rect 38841 23069 38853 23072
rect 38887 23069 38899 23103
rect 38841 23063 38899 23069
rect 38989 23103 39028 23109
rect 38989 23069 39001 23103
rect 38989 23063 39028 23069
rect 39022 23060 39028 23063
rect 39080 23060 39086 23112
rect 39390 23109 39396 23112
rect 39347 23103 39396 23109
rect 39347 23069 39359 23103
rect 39393 23069 39396 23103
rect 39347 23063 39396 23069
rect 39390 23060 39396 23063
rect 39448 23060 39454 23112
rect 40034 23060 40040 23112
rect 40092 23060 40098 23112
rect 40310 23060 40316 23112
rect 40368 23060 40374 23112
rect 40420 23109 40448 23208
rect 40589 23171 40647 23177
rect 40589 23137 40601 23171
rect 40635 23168 40647 23171
rect 42702 23168 42708 23180
rect 40635 23140 42708 23168
rect 40635 23137 40647 23140
rect 40589 23131 40647 23137
rect 42702 23128 42708 23140
rect 42760 23128 42766 23180
rect 42889 23171 42947 23177
rect 42889 23137 42901 23171
rect 42935 23168 42947 23171
rect 43254 23168 43260 23180
rect 42935 23140 43260 23168
rect 42935 23137 42947 23140
rect 42889 23131 42947 23137
rect 43254 23128 43260 23140
rect 43312 23128 43318 23180
rect 40405 23103 40463 23109
rect 40405 23069 40417 23103
rect 40451 23069 40463 23103
rect 40405 23063 40463 23069
rect 34204 23004 37872 23032
rect 34204 22992 34210 23004
rect 39114 22992 39120 23044
rect 39172 22992 39178 23044
rect 39209 23035 39267 23041
rect 39209 23001 39221 23035
rect 39255 23032 39267 23035
rect 39255 23004 42656 23032
rect 39255 23001 39267 23004
rect 39209 22995 39267 23001
rect 33376 22936 33824 22964
rect 33376 22924 33382 22936
rect 34606 22924 34612 22976
rect 34664 22964 34670 22976
rect 35437 22967 35495 22973
rect 35437 22964 35449 22967
rect 34664 22936 35449 22964
rect 34664 22924 34670 22936
rect 35437 22933 35449 22936
rect 35483 22933 35495 22967
rect 35437 22927 35495 22933
rect 36998 22924 37004 22976
rect 37056 22924 37062 22976
rect 39022 22924 39028 22976
rect 39080 22964 39086 22976
rect 39224 22964 39252 22995
rect 39080 22936 39252 22964
rect 39080 22924 39086 22936
rect 42058 22924 42064 22976
rect 42116 22964 42122 22976
rect 42628 22973 42656 23004
rect 42245 22967 42303 22973
rect 42245 22964 42257 22967
rect 42116 22936 42257 22964
rect 42116 22924 42122 22936
rect 42245 22933 42257 22936
rect 42291 22933 42303 22967
rect 42245 22927 42303 22933
rect 42613 22967 42671 22973
rect 42613 22933 42625 22967
rect 42659 22964 42671 22967
rect 43162 22964 43168 22976
rect 42659 22936 43168 22964
rect 42659 22933 42671 22936
rect 42613 22927 42671 22933
rect 43162 22924 43168 22936
rect 43220 22924 43226 22976
rect 1104 22874 43884 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 43884 22874
rect 1104 22800 43884 22822
rect 13909 22763 13967 22769
rect 13909 22729 13921 22763
rect 13955 22760 13967 22763
rect 15102 22760 15108 22772
rect 13955 22732 15108 22760
rect 13955 22729 13967 22732
rect 13909 22723 13967 22729
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 16942 22720 16948 22772
rect 17000 22720 17006 22772
rect 18325 22763 18383 22769
rect 18325 22729 18337 22763
rect 18371 22760 18383 22763
rect 18874 22760 18880 22772
rect 18371 22732 18880 22760
rect 18371 22729 18383 22732
rect 18325 22723 18383 22729
rect 18874 22720 18880 22732
rect 18932 22760 18938 22772
rect 19150 22760 19156 22772
rect 18932 22732 19156 22760
rect 18932 22720 18938 22732
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 20349 22763 20407 22769
rect 20349 22729 20361 22763
rect 20395 22760 20407 22763
rect 20530 22760 20536 22772
rect 20395 22732 20536 22760
rect 20395 22729 20407 22732
rect 20349 22723 20407 22729
rect 20530 22720 20536 22732
rect 20588 22720 20594 22772
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 23474 22760 23480 22772
rect 22612 22732 23480 22760
rect 22612 22720 22618 22732
rect 23474 22720 23480 22732
rect 23532 22760 23538 22772
rect 23661 22763 23719 22769
rect 23661 22760 23673 22763
rect 23532 22732 23673 22760
rect 23532 22720 23538 22732
rect 23661 22729 23673 22732
rect 23707 22729 23719 22763
rect 23661 22723 23719 22729
rect 24394 22720 24400 22772
rect 24452 22760 24458 22772
rect 24673 22763 24731 22769
rect 24673 22760 24685 22763
rect 24452 22732 24685 22760
rect 24452 22720 24458 22732
rect 24673 22729 24685 22732
rect 24719 22729 24731 22763
rect 24673 22723 24731 22729
rect 27982 22720 27988 22772
rect 28040 22760 28046 22772
rect 28553 22763 28611 22769
rect 28553 22760 28565 22763
rect 28040 22732 28565 22760
rect 28040 22720 28046 22732
rect 28553 22729 28565 22732
rect 28599 22729 28611 22763
rect 28553 22723 28611 22729
rect 31386 22720 31392 22772
rect 31444 22760 31450 22772
rect 35621 22763 35679 22769
rect 31444 22732 35572 22760
rect 31444 22720 31450 22732
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 16758 22584 16764 22636
rect 16816 22624 16822 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16816 22596 16865 22624
rect 16816 22584 16822 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16960 22624 16988 22720
rect 17129 22695 17187 22701
rect 17129 22661 17141 22695
rect 17175 22692 17187 22695
rect 18046 22692 18052 22704
rect 17175 22664 18052 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 18046 22652 18052 22664
rect 18104 22652 18110 22704
rect 22186 22692 22192 22704
rect 18708 22664 22192 22692
rect 18322 22633 18328 22636
rect 18266 22627 18328 22633
rect 18266 22624 18278 22627
rect 16960 22596 18278 22624
rect 16853 22587 16911 22593
rect 18266 22593 18278 22596
rect 18312 22593 18328 22627
rect 18266 22587 18328 22593
rect 13630 22516 13636 22568
rect 13688 22516 13694 22568
rect 16868 22556 16896 22587
rect 18322 22584 18328 22587
rect 18380 22584 18386 22636
rect 18708 22633 18736 22664
rect 22186 22652 22192 22664
rect 22244 22652 22250 22704
rect 25314 22652 25320 22704
rect 25372 22652 25378 22704
rect 27617 22695 27675 22701
rect 27617 22661 27629 22695
rect 27663 22692 27675 22695
rect 27663 22664 28304 22692
rect 27663 22661 27675 22664
rect 27617 22655 27675 22661
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 18782 22584 18788 22636
rect 18840 22584 18846 22636
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 20303 22596 21220 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 21192 22568 21220 22596
rect 23842 22584 23848 22636
rect 23900 22584 23906 22636
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22624 25007 22627
rect 25332 22624 25360 22652
rect 24995 22596 25360 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 27473 22627 27531 22633
rect 27473 22624 27485 22627
rect 27120 22596 27485 22624
rect 27120 22584 27126 22596
rect 27473 22593 27485 22596
rect 27519 22593 27531 22627
rect 27473 22587 27531 22593
rect 27706 22584 27712 22636
rect 27764 22584 27770 22636
rect 27890 22584 27896 22636
rect 27948 22584 27954 22636
rect 28276 22624 28304 22664
rect 28350 22652 28356 22704
rect 28408 22652 28414 22704
rect 33318 22692 33324 22704
rect 29656 22664 33324 22692
rect 29656 22624 29684 22664
rect 33318 22652 33324 22664
rect 33376 22652 33382 22704
rect 33686 22652 33692 22704
rect 33744 22692 33750 22704
rect 33873 22695 33931 22701
rect 33873 22692 33885 22695
rect 33744 22664 33885 22692
rect 33744 22652 33750 22664
rect 33873 22661 33885 22664
rect 33919 22661 33931 22695
rect 33873 22655 33931 22661
rect 35250 22652 35256 22704
rect 35308 22652 35314 22704
rect 35544 22692 35572 22732
rect 35621 22729 35633 22763
rect 35667 22760 35679 22763
rect 35802 22760 35808 22772
rect 35667 22732 35808 22760
rect 35667 22729 35679 22732
rect 35621 22723 35679 22729
rect 35802 22720 35808 22732
rect 35860 22720 35866 22772
rect 36170 22720 36176 22772
rect 36228 22720 36234 22772
rect 38105 22763 38163 22769
rect 38105 22729 38117 22763
rect 38151 22760 38163 22763
rect 40310 22760 40316 22772
rect 38151 22732 40316 22760
rect 38151 22729 38163 22732
rect 38105 22723 38163 22729
rect 40310 22720 40316 22732
rect 40368 22720 40374 22772
rect 37553 22695 37611 22701
rect 37553 22692 37565 22695
rect 35544 22664 37565 22692
rect 37553 22661 37565 22664
rect 37599 22692 37611 22695
rect 39301 22695 39359 22701
rect 39301 22692 39313 22695
rect 37599 22664 39313 22692
rect 37599 22661 37611 22664
rect 37553 22655 37611 22661
rect 39301 22661 39313 22664
rect 39347 22661 39359 22695
rect 39301 22655 39359 22661
rect 30098 22624 30104 22636
rect 28276 22596 29684 22624
rect 29840 22596 30104 22624
rect 17034 22556 17040 22568
rect 16868 22528 17040 22556
rect 17034 22516 17040 22528
rect 17092 22516 17098 22568
rect 20530 22516 20536 22568
rect 20588 22516 20594 22568
rect 21174 22516 21180 22568
rect 21232 22556 21238 22568
rect 24029 22559 24087 22565
rect 24029 22556 24041 22559
rect 21232 22528 24041 22556
rect 21232 22516 21238 22528
rect 24029 22525 24041 22528
rect 24075 22556 24087 22559
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 24075 22528 24869 22556
rect 24075 22525 24087 22528
rect 24029 22519 24087 22525
rect 24857 22525 24869 22528
rect 24903 22556 24915 22559
rect 25222 22556 25228 22568
rect 24903 22528 25228 22556
rect 24903 22525 24915 22528
rect 24857 22519 24915 22525
rect 25222 22516 25228 22528
rect 25280 22516 25286 22568
rect 25317 22559 25375 22565
rect 25317 22525 25329 22559
rect 25363 22556 25375 22559
rect 25590 22556 25596 22568
rect 25363 22528 25596 22556
rect 25363 22525 25375 22528
rect 25317 22519 25375 22525
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 26050 22516 26056 22568
rect 26108 22556 26114 22568
rect 29733 22559 29791 22565
rect 29733 22556 29745 22559
rect 26108 22528 29745 22556
rect 26108 22516 26114 22528
rect 29733 22525 29745 22528
rect 29779 22525 29791 22559
rect 29733 22519 29791 22525
rect 22002 22448 22008 22500
rect 22060 22488 22066 22500
rect 22186 22488 22192 22500
rect 22060 22460 22192 22488
rect 22060 22448 22066 22460
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 27341 22491 27399 22497
rect 27341 22488 27353 22491
rect 23584 22460 27353 22488
rect 17129 22423 17187 22429
rect 17129 22389 17141 22423
rect 17175 22420 17187 22423
rect 17218 22420 17224 22432
rect 17175 22392 17224 22420
rect 17175 22389 17187 22392
rect 17129 22383 17187 22389
rect 17218 22380 17224 22392
rect 17276 22380 17282 22432
rect 17310 22380 17316 22432
rect 17368 22420 17374 22432
rect 18141 22423 18199 22429
rect 18141 22420 18153 22423
rect 17368 22392 18153 22420
rect 17368 22380 17374 22392
rect 18141 22389 18153 22392
rect 18187 22389 18199 22423
rect 18141 22383 18199 22389
rect 19886 22380 19892 22432
rect 19944 22380 19950 22432
rect 20438 22380 20444 22432
rect 20496 22420 20502 22432
rect 23584 22420 23612 22460
rect 27341 22457 27353 22460
rect 27387 22457 27399 22491
rect 27341 22451 27399 22457
rect 27890 22448 27896 22500
rect 27948 22488 27954 22500
rect 27948 22460 29500 22488
rect 27948 22448 27954 22460
rect 20496 22392 23612 22420
rect 20496 22380 20502 22392
rect 24946 22380 24952 22432
rect 25004 22420 25010 22432
rect 25590 22420 25596 22432
rect 25004 22392 25596 22420
rect 25004 22380 25010 22392
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 27430 22380 27436 22432
rect 27488 22420 27494 22432
rect 28537 22423 28595 22429
rect 28537 22420 28549 22423
rect 27488 22392 28549 22420
rect 27488 22380 27494 22392
rect 28537 22389 28549 22392
rect 28583 22389 28595 22423
rect 28537 22383 28595 22389
rect 28721 22423 28779 22429
rect 28721 22389 28733 22423
rect 28767 22420 28779 22423
rect 28902 22420 28908 22432
rect 28767 22392 28908 22420
rect 28767 22389 28779 22392
rect 28721 22383 28779 22389
rect 28902 22380 28908 22392
rect 28960 22380 28966 22432
rect 29472 22420 29500 22460
rect 29546 22448 29552 22500
rect 29604 22488 29610 22500
rect 29840 22488 29868 22596
rect 30098 22584 30104 22596
rect 30156 22584 30162 22636
rect 30193 22627 30251 22633
rect 30193 22593 30205 22627
rect 30239 22624 30251 22627
rect 30282 22624 30288 22636
rect 30239 22596 30288 22624
rect 30239 22593 30251 22596
rect 30193 22587 30251 22593
rect 30282 22584 30288 22596
rect 30340 22584 30346 22636
rect 30834 22584 30840 22636
rect 30892 22584 30898 22636
rect 31110 22584 31116 22636
rect 31168 22624 31174 22636
rect 31205 22627 31263 22633
rect 31205 22624 31217 22627
rect 31168 22596 31217 22624
rect 31168 22584 31174 22596
rect 31205 22593 31217 22596
rect 31251 22593 31263 22627
rect 31205 22587 31263 22593
rect 32122 22584 32128 22636
rect 32180 22624 32186 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 32180 22596 33609 22624
rect 32180 22584 32186 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33778 22584 33784 22636
rect 33836 22584 33842 22636
rect 33965 22627 34023 22633
rect 33965 22593 33977 22627
rect 34011 22624 34023 22627
rect 34238 22624 34244 22636
rect 34011 22596 34244 22624
rect 34011 22593 34023 22596
rect 33965 22587 34023 22593
rect 34238 22584 34244 22596
rect 34296 22584 34302 22636
rect 34514 22584 34520 22636
rect 34572 22624 34578 22636
rect 35069 22627 35127 22633
rect 35069 22624 35081 22627
rect 34572 22596 35081 22624
rect 34572 22584 34578 22596
rect 35069 22593 35081 22596
rect 35115 22593 35127 22627
rect 35069 22587 35127 22593
rect 35342 22584 35348 22636
rect 35400 22584 35406 22636
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22593 35495 22627
rect 35437 22587 35495 22593
rect 29917 22559 29975 22565
rect 29917 22525 29929 22559
rect 29963 22556 29975 22559
rect 30374 22556 30380 22568
rect 29963 22528 30380 22556
rect 29963 22525 29975 22528
rect 29917 22519 29975 22525
rect 30374 22516 30380 22528
rect 30432 22516 30438 22568
rect 30653 22559 30711 22565
rect 30653 22525 30665 22559
rect 30699 22556 30711 22559
rect 31478 22556 31484 22568
rect 30699 22528 31484 22556
rect 30699 22525 30711 22528
rect 30653 22519 30711 22525
rect 31478 22516 31484 22528
rect 31536 22556 31542 22568
rect 34256 22556 34284 22584
rect 35452 22556 35480 22587
rect 35526 22584 35532 22636
rect 35584 22624 35590 22636
rect 36081 22627 36139 22633
rect 36081 22624 36093 22627
rect 35584 22596 36093 22624
rect 35584 22584 35590 22596
rect 36081 22593 36093 22596
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 36265 22627 36323 22633
rect 36265 22593 36277 22627
rect 36311 22593 36323 22627
rect 36265 22587 36323 22593
rect 31536 22528 31754 22556
rect 34256 22528 35480 22556
rect 31536 22516 31542 22528
rect 29604 22460 29868 22488
rect 29604 22448 29610 22460
rect 31110 22448 31116 22500
rect 31168 22448 31174 22500
rect 30098 22420 30104 22432
rect 29472 22392 30104 22420
rect 30098 22380 30104 22392
rect 30156 22380 30162 22432
rect 31726 22420 31754 22528
rect 35986 22516 35992 22568
rect 36044 22556 36050 22568
rect 36280 22556 36308 22587
rect 37826 22584 37832 22636
rect 37884 22584 37890 22636
rect 38654 22584 38660 22636
rect 38712 22624 38718 22636
rect 38838 22624 38844 22636
rect 38712 22596 38844 22624
rect 38712 22584 38718 22596
rect 38838 22584 38844 22596
rect 38896 22624 38902 22636
rect 38933 22627 38991 22633
rect 38933 22624 38945 22627
rect 38896 22596 38945 22624
rect 38896 22584 38902 22596
rect 38933 22593 38945 22596
rect 38979 22593 38991 22627
rect 38933 22587 38991 22593
rect 39022 22584 39028 22636
rect 39080 22624 39086 22636
rect 39080 22596 39125 22624
rect 39080 22584 39086 22596
rect 39206 22584 39212 22636
rect 39264 22584 39270 22636
rect 39439 22627 39497 22633
rect 39439 22624 39451 22627
rect 39316 22596 39451 22624
rect 39316 22568 39344 22596
rect 39439 22593 39451 22596
rect 39485 22624 39497 22627
rect 39574 22624 39580 22636
rect 39485 22596 39580 22624
rect 39485 22593 39497 22596
rect 39439 22587 39497 22593
rect 39574 22584 39580 22596
rect 39632 22584 39638 22636
rect 36044 22528 36308 22556
rect 36044 22516 36050 22528
rect 36538 22516 36544 22568
rect 36596 22556 36602 22568
rect 37274 22556 37280 22568
rect 36596 22528 37280 22556
rect 36596 22516 36602 22528
rect 37274 22516 37280 22528
rect 37332 22516 37338 22568
rect 37461 22559 37519 22565
rect 37461 22525 37473 22559
rect 37507 22556 37519 22559
rect 37550 22556 37556 22568
rect 37507 22528 37556 22556
rect 37507 22525 37519 22528
rect 37461 22519 37519 22525
rect 37550 22516 37556 22528
rect 37608 22516 37614 22568
rect 37921 22559 37979 22565
rect 37921 22525 37933 22559
rect 37967 22525 37979 22559
rect 37921 22519 37979 22525
rect 34146 22448 34152 22500
rect 34204 22448 34210 22500
rect 34238 22448 34244 22500
rect 34296 22488 34302 22500
rect 34296 22460 36860 22488
rect 34296 22448 34302 22460
rect 36538 22420 36544 22432
rect 31726 22392 36544 22420
rect 36538 22380 36544 22392
rect 36596 22380 36602 22432
rect 36832 22420 36860 22460
rect 37366 22448 37372 22500
rect 37424 22488 37430 22500
rect 37936 22488 37964 22519
rect 39298 22516 39304 22568
rect 39356 22516 39362 22568
rect 37424 22460 37964 22488
rect 37424 22448 37430 22460
rect 39206 22420 39212 22432
rect 36832 22392 39212 22420
rect 39206 22380 39212 22392
rect 39264 22380 39270 22432
rect 39574 22380 39580 22432
rect 39632 22380 39638 22432
rect 1104 22330 43884 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 43884 22330
rect 1104 22256 43884 22278
rect 13541 22219 13599 22225
rect 13541 22185 13553 22219
rect 13587 22216 13599 22219
rect 13630 22216 13636 22228
rect 13587 22188 13636 22216
rect 13587 22185 13599 22188
rect 13541 22179 13599 22185
rect 13630 22176 13636 22188
rect 13688 22176 13694 22228
rect 20530 22176 20536 22228
rect 20588 22216 20594 22228
rect 20625 22219 20683 22225
rect 20625 22216 20637 22219
rect 20588 22188 20637 22216
rect 20588 22176 20594 22188
rect 20625 22185 20637 22188
rect 20671 22185 20683 22219
rect 20625 22179 20683 22185
rect 23842 22176 23848 22228
rect 23900 22216 23906 22228
rect 25222 22216 25228 22228
rect 23900 22188 25228 22216
rect 23900 22176 23906 22188
rect 25222 22176 25228 22188
rect 25280 22216 25286 22228
rect 25774 22216 25780 22228
rect 25280 22188 25780 22216
rect 25280 22176 25286 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 31110 22216 31116 22228
rect 25884 22188 31116 22216
rect 20438 22108 20444 22160
rect 20496 22148 20502 22160
rect 20717 22151 20775 22157
rect 20717 22148 20729 22151
rect 20496 22120 20729 22148
rect 20496 22108 20502 22120
rect 20717 22117 20729 22120
rect 20763 22117 20775 22151
rect 20717 22111 20775 22117
rect 21913 22151 21971 22157
rect 21913 22117 21925 22151
rect 21959 22148 21971 22151
rect 22094 22148 22100 22160
rect 21959 22120 22100 22148
rect 21959 22117 21971 22120
rect 21913 22111 21971 22117
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 25884 22148 25912 22188
rect 31110 22176 31116 22188
rect 31168 22176 31174 22228
rect 34790 22216 34796 22228
rect 31726 22188 34796 22216
rect 22204 22120 25912 22148
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 17034 22080 17040 22092
rect 14292 22052 17040 22080
rect 10686 21972 10692 22024
rect 10744 22012 10750 22024
rect 10781 22015 10839 22021
rect 10781 22012 10793 22015
rect 10744 21984 10793 22012
rect 10744 21972 10750 21984
rect 10781 21981 10793 21984
rect 10827 22012 10839 22015
rect 11974 22012 11980 22024
rect 10827 21984 11980 22012
rect 10827 21981 10839 21984
rect 10781 21975 10839 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 13262 21972 13268 22024
rect 13320 21972 13326 22024
rect 11048 21947 11106 21953
rect 11048 21913 11060 21947
rect 11094 21944 11106 21947
rect 14292 21944 14320 22052
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 18690 22040 18696 22092
rect 18748 22080 18754 22092
rect 18785 22083 18843 22089
rect 18785 22080 18797 22083
rect 18748 22052 18797 22080
rect 18748 22040 18754 22052
rect 18785 22049 18797 22052
rect 18831 22049 18843 22083
rect 18785 22043 18843 22049
rect 20346 22040 20352 22092
rect 20404 22080 20410 22092
rect 21085 22083 21143 22089
rect 21085 22080 21097 22083
rect 20404 22052 21097 22080
rect 20404 22040 20410 22052
rect 21085 22049 21097 22052
rect 21131 22080 21143 22083
rect 22204 22080 22232 22120
rect 28626 22108 28632 22160
rect 28684 22148 28690 22160
rect 30193 22151 30251 22157
rect 30193 22148 30205 22151
rect 28684 22120 30205 22148
rect 28684 22108 28690 22120
rect 30193 22117 30205 22120
rect 30239 22148 30251 22151
rect 31726 22148 31754 22188
rect 34790 22176 34796 22188
rect 34848 22176 34854 22228
rect 35986 22176 35992 22228
rect 36044 22216 36050 22228
rect 36630 22216 36636 22228
rect 36044 22188 36636 22216
rect 36044 22176 36050 22188
rect 36630 22176 36636 22188
rect 36688 22176 36694 22228
rect 39485 22219 39543 22225
rect 39485 22185 39497 22219
rect 39531 22216 39543 22219
rect 40126 22216 40132 22228
rect 39531 22188 40132 22216
rect 39531 22185 39543 22188
rect 39485 22179 39543 22185
rect 40126 22176 40132 22188
rect 40184 22176 40190 22228
rect 43162 22176 43168 22228
rect 43220 22176 43226 22228
rect 30239 22120 31754 22148
rect 34885 22151 34943 22157
rect 30239 22117 30251 22120
rect 30193 22111 30251 22117
rect 34885 22117 34897 22151
rect 34931 22117 34943 22151
rect 34885 22111 34943 22117
rect 21131 22052 22232 22080
rect 27540 22052 29960 22080
rect 21131 22049 21143 22052
rect 21085 22043 21143 22049
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 22012 14703 22015
rect 15194 22012 15200 22024
rect 14691 21984 15200 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 15194 21972 15200 21984
rect 15252 22012 15258 22024
rect 15289 22015 15347 22021
rect 15289 22012 15301 22015
rect 15252 21984 15301 22012
rect 15252 21972 15258 21984
rect 15289 21981 15301 21984
rect 15335 22012 15347 22015
rect 17310 22012 17316 22024
rect 15335 21984 17316 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 19484 21984 19809 22012
rect 19484 21972 19490 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 19978 21972 19984 22024
rect 20036 21972 20042 22024
rect 20165 22015 20223 22021
rect 20165 21981 20177 22015
rect 20211 22012 20223 22015
rect 20254 22012 20260 22024
rect 20211 21984 20260 22012
rect 20211 21981 20223 21984
rect 20165 21975 20223 21981
rect 20254 21972 20260 21984
rect 20312 22012 20318 22024
rect 20622 22012 20628 22024
rect 20312 21984 20628 22012
rect 20312 21972 20318 21984
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 22097 22015 22155 22021
rect 22097 22012 22109 22015
rect 21508 21984 22109 22012
rect 21508 21972 21514 21984
rect 22097 21981 22109 21984
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 22186 21972 22192 22024
rect 22244 21972 22250 22024
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 22012 22523 22015
rect 22554 22012 22560 22024
rect 22511 21984 22560 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 11094 21916 14320 21944
rect 14369 21947 14427 21953
rect 11094 21913 11106 21916
rect 11048 21907 11106 21913
rect 14369 21913 14381 21947
rect 14415 21944 14427 21947
rect 15010 21944 15016 21956
rect 14415 21916 15016 21944
rect 14415 21913 14427 21916
rect 14369 21907 14427 21913
rect 15010 21904 15016 21916
rect 15068 21944 15074 21956
rect 15473 21947 15531 21953
rect 15068 21916 15240 21944
rect 15068 21904 15074 21916
rect 12158 21836 12164 21888
rect 12216 21836 12222 21888
rect 12250 21836 12256 21888
rect 12308 21876 12314 21888
rect 14467 21879 14525 21885
rect 14467 21876 14479 21879
rect 12308 21848 14479 21876
rect 12308 21836 12314 21848
rect 14467 21845 14479 21848
rect 14513 21845 14525 21879
rect 14467 21839 14525 21845
rect 14553 21879 14611 21885
rect 14553 21845 14565 21879
rect 14599 21876 14611 21879
rect 14642 21876 14648 21888
rect 14599 21848 14648 21876
rect 14599 21845 14611 21848
rect 14553 21839 14611 21845
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 15102 21836 15108 21888
rect 15160 21836 15166 21888
rect 15212 21876 15240 21916
rect 15473 21913 15485 21947
rect 15519 21913 15531 21947
rect 15473 21907 15531 21913
rect 18509 21947 18567 21953
rect 18509 21913 18521 21947
rect 18555 21944 18567 21947
rect 18690 21944 18696 21956
rect 18555 21916 18696 21944
rect 18555 21913 18567 21916
rect 18509 21907 18567 21913
rect 15488 21876 15516 21907
rect 18690 21904 18696 21916
rect 18748 21904 18754 21956
rect 21266 21944 21272 21956
rect 19444 21916 21272 21944
rect 18141 21879 18199 21885
rect 18141 21876 18153 21879
rect 15212 21848 18153 21876
rect 18141 21845 18153 21848
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 18601 21879 18659 21885
rect 18601 21845 18613 21879
rect 18647 21876 18659 21879
rect 19444 21876 19472 21916
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 21358 21904 21364 21956
rect 21416 21944 21422 21956
rect 22388 21944 22416 21975
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 24854 21972 24860 22024
rect 24912 21972 24918 22024
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 25225 22015 25283 22021
rect 25225 22012 25237 22015
rect 25188 21984 25237 22012
rect 25188 21972 25194 21984
rect 25225 21981 25237 21984
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 27062 21972 27068 22024
rect 27120 22012 27126 22024
rect 27540 22021 27568 22052
rect 27157 22015 27215 22021
rect 27157 22012 27169 22015
rect 27120 21984 27169 22012
rect 27120 21972 27126 21984
rect 27157 21981 27169 21984
rect 27203 21981 27215 22015
rect 27157 21975 27215 21981
rect 27249 22015 27307 22021
rect 27249 21981 27261 22015
rect 27295 22012 27307 22015
rect 27525 22015 27583 22021
rect 27295 21984 27476 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 23014 21944 23020 21956
rect 21416 21916 23020 21944
rect 21416 21904 21422 21916
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 24949 21947 25007 21953
rect 24949 21913 24961 21947
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 25041 21947 25099 21953
rect 25041 21913 25053 21947
rect 25087 21944 25099 21947
rect 25590 21944 25596 21956
rect 25087 21916 25596 21944
rect 25087 21913 25099 21916
rect 25041 21907 25099 21913
rect 18647 21848 19472 21876
rect 19521 21879 19579 21885
rect 18647 21845 18659 21848
rect 18601 21839 18659 21845
rect 19521 21845 19533 21879
rect 19567 21876 19579 21879
rect 19978 21876 19984 21888
rect 19567 21848 19984 21876
rect 19567 21845 19579 21848
rect 19521 21839 19579 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 23290 21876 23296 21888
rect 20220 21848 23296 21876
rect 20220 21836 20226 21848
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 24670 21836 24676 21888
rect 24728 21836 24734 21888
rect 24964 21876 24992 21907
rect 25590 21904 25596 21916
rect 25648 21904 25654 21956
rect 27341 21947 27399 21953
rect 27341 21913 27353 21947
rect 27387 21913 27399 21947
rect 27448 21944 27476 21984
rect 27525 21981 27537 22015
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27614 21972 27620 22024
rect 27672 22012 27678 22024
rect 27982 22012 27988 22024
rect 27672 21984 27988 22012
rect 27672 21972 27678 21984
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 28166 21972 28172 22024
rect 28224 21972 28230 22024
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 29825 22015 29883 22021
rect 29825 22012 29837 22015
rect 28316 21984 29837 22012
rect 28316 21972 28322 21984
rect 29825 21981 29837 21984
rect 29871 21981 29883 22015
rect 29932 22012 29960 22052
rect 30006 22040 30012 22092
rect 30064 22040 30070 22092
rect 31202 22080 31208 22092
rect 30208 22052 31208 22080
rect 30208 22012 30236 22052
rect 31202 22040 31208 22052
rect 31260 22040 31266 22092
rect 32677 22083 32735 22089
rect 32677 22049 32689 22083
rect 32723 22080 32735 22083
rect 33042 22080 33048 22092
rect 32723 22052 33048 22080
rect 32723 22049 32735 22052
rect 32677 22043 32735 22049
rect 33042 22040 33048 22052
rect 33100 22040 33106 22092
rect 29932 21984 30236 22012
rect 29825 21975 29883 21981
rect 30282 21972 30288 22024
rect 30340 21972 30346 22024
rect 33594 22012 33600 22024
rect 33336 21984 33600 22012
rect 30926 21944 30932 21956
rect 27448 21916 30932 21944
rect 27341 21907 27399 21913
rect 25866 21876 25872 21888
rect 24964 21848 25872 21876
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 26970 21836 26976 21888
rect 27028 21836 27034 21888
rect 27356 21876 27384 21907
rect 30926 21904 30932 21916
rect 30984 21904 30990 21956
rect 32306 21904 32312 21956
rect 32364 21944 32370 21956
rect 33336 21953 33364 21984
rect 33594 21972 33600 21984
rect 33652 21972 33658 22024
rect 34900 22012 34928 22111
rect 37918 22108 37924 22160
rect 37976 22148 37982 22160
rect 39114 22148 39120 22160
rect 37976 22120 39120 22148
rect 37976 22108 37982 22120
rect 39114 22108 39120 22120
rect 39172 22108 39178 22160
rect 34974 22040 34980 22092
rect 35032 22080 35038 22092
rect 35032 22052 39344 22080
rect 35032 22040 35038 22052
rect 39316 22021 39344 22052
rect 40402 22040 40408 22092
rect 40460 22080 40466 22092
rect 40497 22083 40555 22089
rect 40497 22080 40509 22083
rect 40460 22052 40509 22080
rect 40460 22040 40466 22052
rect 40497 22049 40509 22052
rect 40543 22049 40555 22083
rect 40497 22043 40555 22049
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 33704 21984 34928 22012
rect 34992 21984 35173 22012
rect 32410 21947 32468 21953
rect 32410 21944 32422 21947
rect 32364 21916 32422 21944
rect 32364 21904 32370 21916
rect 32410 21913 32422 21916
rect 32456 21913 32468 21947
rect 32410 21907 32468 21913
rect 33321 21947 33379 21953
rect 33321 21913 33333 21947
rect 33367 21913 33379 21947
rect 33321 21907 33379 21913
rect 33410 21904 33416 21956
rect 33468 21944 33474 21956
rect 33505 21947 33563 21953
rect 33505 21944 33517 21947
rect 33468 21916 33517 21944
rect 33468 21904 33474 21916
rect 33505 21913 33517 21916
rect 33551 21944 33563 21947
rect 33704 21944 33732 21984
rect 33551 21916 33732 21944
rect 33551 21913 33563 21916
rect 33505 21907 33563 21913
rect 34054 21904 34060 21956
rect 34112 21944 34118 21956
rect 34238 21944 34244 21956
rect 34112 21916 34244 21944
rect 34112 21904 34118 21916
rect 34238 21904 34244 21916
rect 34296 21904 34302 21956
rect 34330 21904 34336 21956
rect 34388 21944 34394 21956
rect 34885 21947 34943 21953
rect 34885 21944 34897 21947
rect 34388 21916 34897 21944
rect 34388 21904 34394 21916
rect 34885 21913 34897 21916
rect 34931 21913 34943 21947
rect 34885 21907 34943 21913
rect 27706 21876 27712 21888
rect 27356 21848 27712 21876
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 28261 21879 28319 21885
rect 28261 21845 28273 21879
rect 28307 21876 28319 21879
rect 29638 21876 29644 21888
rect 28307 21848 29644 21876
rect 28307 21845 28319 21848
rect 28261 21839 28319 21845
rect 29638 21836 29644 21848
rect 29696 21836 29702 21888
rect 31110 21836 31116 21888
rect 31168 21876 31174 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 31168 21848 31309 21876
rect 31168 21836 31174 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 31297 21839 31355 21845
rect 33689 21879 33747 21885
rect 33689 21845 33701 21879
rect 33735 21876 33747 21879
rect 33778 21876 33784 21888
rect 33735 21848 33784 21876
rect 33735 21845 33747 21848
rect 33689 21839 33747 21845
rect 33778 21836 33784 21848
rect 33836 21836 33842 21888
rect 34422 21836 34428 21888
rect 34480 21876 34486 21888
rect 34992 21876 35020 21984
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 39209 22015 39267 22021
rect 39209 21981 39221 22015
rect 39255 21981 39267 22015
rect 39209 21975 39267 21981
rect 39301 22015 39359 22021
rect 39301 21981 39313 22015
rect 39347 22012 39359 22015
rect 40034 22012 40040 22024
rect 39347 21984 40040 22012
rect 39347 21981 39359 21984
rect 39301 21975 39359 21981
rect 39224 21944 39252 21975
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 41785 22015 41843 22021
rect 41785 21981 41797 22015
rect 41831 22012 41843 22015
rect 41874 22012 41880 22024
rect 41831 21984 41880 22012
rect 41831 21981 41843 21984
rect 41785 21975 41843 21981
rect 41874 21972 41880 21984
rect 41932 21972 41938 22024
rect 42058 22021 42064 22024
rect 42052 22012 42064 22021
rect 42019 21984 42064 22012
rect 42052 21975 42064 21984
rect 42058 21972 42064 21975
rect 42116 21972 42122 22024
rect 39485 21947 39543 21953
rect 39224 21916 39344 21944
rect 39316 21888 39344 21916
rect 39485 21913 39497 21947
rect 39531 21913 39543 21947
rect 39485 21907 39543 21913
rect 34480 21848 35020 21876
rect 34480 21836 34486 21848
rect 35066 21836 35072 21888
rect 35124 21876 35130 21888
rect 35342 21876 35348 21888
rect 35124 21848 35348 21876
rect 35124 21836 35130 21848
rect 35342 21836 35348 21848
rect 35400 21836 35406 21888
rect 39298 21836 39304 21888
rect 39356 21836 39362 21888
rect 39500 21876 39528 21907
rect 40126 21904 40132 21956
rect 40184 21904 40190 21956
rect 40313 21947 40371 21953
rect 40313 21913 40325 21947
rect 40359 21913 40371 21947
rect 40313 21907 40371 21913
rect 39574 21876 39580 21888
rect 39500 21848 39580 21876
rect 39574 21836 39580 21848
rect 39632 21836 39638 21888
rect 39758 21836 39764 21888
rect 39816 21876 39822 21888
rect 40328 21876 40356 21907
rect 39816 21848 40356 21876
rect 39816 21836 39822 21848
rect 1104 21786 43884 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 43884 21786
rect 1104 21712 43884 21734
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 23198 21672 23204 21684
rect 16264 21644 23204 21672
rect 16264 21632 16270 21644
rect 20180 21613 20208 21644
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 24670 21632 24676 21684
rect 24728 21672 24734 21684
rect 24949 21675 25007 21681
rect 24949 21672 24961 21675
rect 24728 21644 24961 21672
rect 24728 21632 24734 21644
rect 24949 21641 24961 21644
rect 24995 21641 25007 21675
rect 24949 21635 25007 21641
rect 25590 21632 25596 21684
rect 25648 21632 25654 21684
rect 27522 21632 27528 21684
rect 27580 21672 27586 21684
rect 27982 21672 27988 21684
rect 27580 21644 27988 21672
rect 27580 21632 27586 21644
rect 27982 21632 27988 21644
rect 28040 21632 28046 21684
rect 31110 21672 31116 21684
rect 28276 21644 31116 21672
rect 15197 21607 15255 21613
rect 15197 21573 15209 21607
rect 15243 21604 15255 21607
rect 20165 21607 20223 21613
rect 15243 21576 15884 21604
rect 15243 21573 15255 21576
rect 15197 21567 15255 21573
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 14642 21496 14648 21548
rect 14700 21536 14706 21548
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 14700 21508 14933 21536
rect 14700 21496 14706 21508
rect 14921 21505 14933 21508
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 15010 21496 15016 21548
rect 15068 21496 15074 21548
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 15856 21545 15884 21576
rect 20165 21573 20177 21607
rect 20211 21573 20223 21607
rect 20165 21567 20223 21573
rect 20346 21564 20352 21616
rect 20404 21564 20410 21616
rect 21177 21607 21235 21613
rect 21177 21573 21189 21607
rect 21223 21604 21235 21607
rect 28074 21604 28080 21616
rect 21223 21576 22416 21604
rect 21223 21573 21235 21576
rect 21177 21567 21235 21573
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 15160 21508 15669 21536
rect 15160 21496 15166 21508
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 16114 21496 16120 21548
rect 16172 21536 16178 21548
rect 21358 21536 21364 21548
rect 16172 21508 21364 21536
rect 16172 21496 16178 21508
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 22094 21496 22100 21548
rect 22152 21496 22158 21548
rect 22388 21545 22416 21576
rect 24320 21576 28080 21604
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22646 21496 22652 21548
rect 22704 21496 22710 21548
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 12158 21428 12164 21480
rect 12216 21428 12222 21480
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21468 12495 21471
rect 13538 21468 13544 21480
rect 12483 21440 13544 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 15194 21428 15200 21480
rect 15252 21428 15258 21480
rect 16850 21428 16856 21480
rect 16908 21428 16914 21480
rect 17126 21428 17132 21480
rect 17184 21428 17190 21480
rect 21174 21428 21180 21480
rect 21232 21428 21238 21480
rect 21468 21468 21496 21496
rect 22940 21468 22968 21499
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 24320 21536 24348 21576
rect 28074 21564 28080 21576
rect 28132 21564 28138 21616
rect 23072 21508 24348 21536
rect 23072 21496 23078 21508
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25682 21536 25688 21548
rect 24912 21508 25688 21536
rect 24912 21496 24918 21508
rect 25682 21496 25688 21508
rect 25740 21536 25746 21548
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25740 21508 25789 21536
rect 25740 21496 25746 21508
rect 25777 21505 25789 21508
rect 25823 21505 25835 21539
rect 25777 21499 25835 21505
rect 25866 21496 25872 21548
rect 25924 21496 25930 21548
rect 27433 21539 27491 21545
rect 27433 21505 27445 21539
rect 27479 21536 27491 21539
rect 27522 21536 27528 21548
rect 27479 21508 27528 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 27706 21496 27712 21548
rect 27764 21536 27770 21548
rect 27890 21536 27896 21548
rect 27764 21508 27896 21536
rect 27764 21496 27770 21508
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21536 28227 21539
rect 28276 21536 28304 21644
rect 31110 21632 31116 21644
rect 31168 21672 31174 21684
rect 31168 21644 34376 21672
rect 31168 21632 31174 21644
rect 31202 21564 31208 21616
rect 31260 21564 31266 21616
rect 31294 21564 31300 21616
rect 31352 21604 31358 21616
rect 31389 21607 31447 21613
rect 31389 21604 31401 21607
rect 31352 21576 31401 21604
rect 31352 21564 31358 21576
rect 31389 21573 31401 21576
rect 31435 21573 31447 21607
rect 31389 21567 31447 21573
rect 32232 21576 33916 21604
rect 28215 21508 28304 21536
rect 28629 21539 28687 21545
rect 28215 21505 28227 21508
rect 28169 21499 28227 21505
rect 28629 21505 28641 21539
rect 28675 21505 28687 21539
rect 28629 21499 28687 21505
rect 21468 21440 23060 21468
rect 13262 21360 13268 21412
rect 13320 21400 13326 21412
rect 13722 21400 13728 21412
rect 13320 21372 13728 21400
rect 13320 21360 13326 21372
rect 13722 21360 13728 21372
rect 13780 21400 13786 21412
rect 20162 21400 20168 21412
rect 13780 21372 15884 21400
rect 13780 21360 13786 21372
rect 15746 21292 15752 21344
rect 15804 21292 15810 21344
rect 15856 21332 15884 21372
rect 17788 21372 20168 21400
rect 17788 21332 17816 21372
rect 20162 21360 20168 21372
rect 20220 21360 20226 21412
rect 23032 21400 23060 21440
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 24471 21471 24529 21477
rect 24471 21468 24483 21471
rect 23256 21440 24483 21468
rect 23256 21428 23262 21440
rect 24471 21437 24483 21440
rect 24517 21437 24529 21471
rect 24471 21431 24529 21437
rect 24946 21428 24952 21480
rect 25004 21428 25010 21480
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 25590 21428 25596 21480
rect 25648 21428 25654 21480
rect 27062 21428 27068 21480
rect 27120 21468 27126 21480
rect 28534 21468 28540 21480
rect 27120 21440 28540 21468
rect 27120 21428 27126 21440
rect 28534 21428 28540 21440
rect 28592 21468 28598 21480
rect 28644 21468 28672 21499
rect 28592 21440 28672 21468
rect 28592 21428 28598 21440
rect 30466 21428 30472 21480
rect 30524 21468 30530 21480
rect 31110 21468 31116 21480
rect 30524 21440 31116 21468
rect 30524 21428 30530 21440
rect 31110 21428 31116 21440
rect 31168 21428 31174 21480
rect 32232 21468 32260 21576
rect 32677 21539 32735 21545
rect 32677 21505 32689 21539
rect 32723 21536 32735 21539
rect 33410 21536 33416 21548
rect 32723 21508 33416 21536
rect 32723 21505 32735 21508
rect 32677 21499 32735 21505
rect 33410 21496 33416 21508
rect 33468 21496 33474 21548
rect 31726 21440 32260 21468
rect 27249 21403 27307 21409
rect 27249 21400 27261 21403
rect 23032 21372 27261 21400
rect 27249 21369 27261 21372
rect 27295 21369 27307 21403
rect 27249 21363 27307 21369
rect 29362 21360 29368 21412
rect 29420 21400 29426 21412
rect 31726 21400 31754 21440
rect 32306 21428 32312 21480
rect 32364 21428 32370 21480
rect 32769 21471 32827 21477
rect 32769 21437 32781 21471
rect 32815 21468 32827 21471
rect 33594 21468 33600 21480
rect 32815 21440 33600 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 33594 21428 33600 21440
rect 33652 21428 33658 21480
rect 29420 21372 31754 21400
rect 29420 21360 29426 21372
rect 15856 21304 17816 21332
rect 18414 21292 18420 21344
rect 18472 21292 18478 21344
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 22738 21292 22744 21344
rect 22796 21332 22802 21344
rect 23385 21335 23443 21341
rect 23385 21332 23397 21335
rect 22796 21304 23397 21332
rect 22796 21292 22802 21304
rect 23385 21301 23397 21304
rect 23431 21301 23443 21335
rect 23385 21295 23443 21301
rect 24854 21292 24860 21344
rect 24912 21332 24918 21344
rect 25590 21332 25596 21344
rect 24912 21304 25596 21332
rect 24912 21292 24918 21304
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 31665 21335 31723 21341
rect 31665 21301 31677 21335
rect 31711 21332 31723 21335
rect 33134 21332 33140 21344
rect 31711 21304 33140 21332
rect 31711 21301 31723 21304
rect 31665 21295 31723 21301
rect 33134 21292 33140 21304
rect 33192 21292 33198 21344
rect 33704 21332 33732 21576
rect 33781 21539 33839 21545
rect 33781 21505 33793 21539
rect 33827 21505 33839 21539
rect 33888 21536 33916 21576
rect 33962 21564 33968 21616
rect 34020 21564 34026 21616
rect 34348 21604 34376 21644
rect 34698 21632 34704 21684
rect 34756 21672 34762 21684
rect 35618 21672 35624 21684
rect 34756 21644 35624 21672
rect 34756 21632 34762 21644
rect 35618 21632 35624 21644
rect 35676 21632 35682 21684
rect 37458 21632 37464 21684
rect 37516 21672 37522 21684
rect 39206 21672 39212 21684
rect 37516 21644 37872 21672
rect 37516 21632 37522 21644
rect 35066 21604 35072 21616
rect 34348 21576 35072 21604
rect 35066 21564 35072 21576
rect 35124 21604 35130 21616
rect 35713 21607 35771 21613
rect 35713 21604 35725 21607
rect 35124 21576 35725 21604
rect 35124 21564 35130 21576
rect 35713 21573 35725 21576
rect 35759 21573 35771 21607
rect 35713 21567 35771 21573
rect 37274 21564 37280 21616
rect 37332 21604 37338 21616
rect 37737 21607 37795 21613
rect 37737 21604 37749 21607
rect 37332 21576 37749 21604
rect 37332 21564 37338 21576
rect 37737 21573 37749 21576
rect 37783 21573 37795 21607
rect 37737 21567 37795 21573
rect 34057 21539 34115 21545
rect 34057 21536 34069 21539
rect 33888 21508 34069 21536
rect 33781 21499 33839 21505
rect 34057 21505 34069 21508
rect 34103 21505 34115 21539
rect 34057 21499 34115 21505
rect 33796 21400 33824 21499
rect 34146 21496 34152 21548
rect 34204 21496 34210 21548
rect 35437 21539 35495 21545
rect 35437 21505 35449 21539
rect 35483 21536 35495 21539
rect 35483 21508 36216 21536
rect 35483 21505 35495 21508
rect 35437 21499 35495 21505
rect 34514 21468 34520 21480
rect 34440 21440 34520 21468
rect 34238 21400 34244 21412
rect 33796 21372 34244 21400
rect 34238 21360 34244 21372
rect 34296 21360 34302 21412
rect 34330 21360 34336 21412
rect 34388 21360 34394 21412
rect 34440 21332 34468 21440
rect 34514 21428 34520 21440
rect 34572 21468 34578 21480
rect 34698 21468 34704 21480
rect 34572 21440 34704 21468
rect 34572 21428 34578 21440
rect 34698 21428 34704 21440
rect 34756 21428 34762 21480
rect 34790 21428 34796 21480
rect 34848 21468 34854 21480
rect 35345 21471 35403 21477
rect 35345 21468 35357 21471
rect 34848 21440 35357 21468
rect 34848 21428 34854 21440
rect 35345 21437 35357 21440
rect 35391 21468 35403 21471
rect 35526 21468 35532 21480
rect 35391 21440 35532 21468
rect 35391 21437 35403 21440
rect 35345 21431 35403 21437
rect 35526 21428 35532 21440
rect 35584 21428 35590 21480
rect 35805 21471 35863 21477
rect 35805 21437 35817 21471
rect 35851 21468 35863 21471
rect 36078 21468 36084 21480
rect 35851 21440 36084 21468
rect 35851 21437 35863 21440
rect 35805 21431 35863 21437
rect 36078 21428 36084 21440
rect 36136 21428 36142 21480
rect 36188 21468 36216 21508
rect 36262 21496 36268 21548
rect 36320 21536 36326 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 36320 21508 37473 21536
rect 36320 21496 36326 21508
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 37461 21499 37519 21505
rect 37550 21496 37556 21548
rect 37608 21536 37614 21548
rect 37844 21545 37872 21644
rect 38948 21644 39212 21672
rect 38948 21613 38976 21644
rect 39206 21632 39212 21644
rect 39264 21632 39270 21684
rect 39298 21632 39304 21684
rect 39356 21672 39362 21684
rect 39942 21672 39948 21684
rect 39356 21644 39948 21672
rect 39356 21632 39362 21644
rect 39942 21632 39948 21644
rect 40000 21632 40006 21684
rect 40034 21632 40040 21684
rect 40092 21672 40098 21684
rect 40681 21675 40739 21681
rect 40681 21672 40693 21675
rect 40092 21644 40693 21672
rect 40092 21632 40098 21644
rect 40681 21641 40693 21644
rect 40727 21641 40739 21675
rect 40681 21635 40739 21641
rect 38933 21607 38991 21613
rect 38933 21573 38945 21607
rect 38979 21573 38991 21607
rect 38933 21567 38991 21573
rect 43162 21564 43168 21616
rect 43220 21564 43226 21616
rect 37645 21539 37703 21545
rect 37645 21536 37657 21539
rect 37608 21508 37657 21536
rect 37608 21496 37614 21508
rect 37645 21505 37657 21508
rect 37691 21505 37703 21539
rect 37645 21499 37703 21505
rect 37829 21539 37887 21545
rect 37829 21505 37841 21539
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 38654 21496 38660 21548
rect 38712 21496 38718 21548
rect 38746 21496 38752 21548
rect 38804 21536 38810 21548
rect 39025 21539 39083 21545
rect 38804 21508 38849 21536
rect 38804 21496 38810 21508
rect 39025 21505 39037 21539
rect 39071 21505 39083 21539
rect 39025 21499 39083 21505
rect 39163 21539 39221 21545
rect 39163 21505 39175 21539
rect 39209 21536 39221 21539
rect 39390 21536 39396 21548
rect 39209 21508 39396 21536
rect 39209 21505 39221 21508
rect 39163 21499 39221 21505
rect 37182 21468 37188 21480
rect 36188 21440 37188 21468
rect 37182 21428 37188 21440
rect 37240 21468 37246 21480
rect 37734 21468 37740 21480
rect 37240 21440 37740 21468
rect 37240 21428 37246 21440
rect 37734 21428 37740 21440
rect 37792 21428 37798 21480
rect 39040 21468 39068 21499
rect 39390 21496 39396 21508
rect 39448 21496 39454 21548
rect 40586 21496 40592 21548
rect 40644 21536 40650 21548
rect 41794 21539 41852 21545
rect 41794 21536 41806 21539
rect 40644 21508 41806 21536
rect 40644 21496 40650 21508
rect 41794 21505 41806 21508
rect 41840 21505 41852 21539
rect 41794 21499 41852 21505
rect 41966 21496 41972 21548
rect 42024 21536 42030 21548
rect 42061 21539 42119 21545
rect 42061 21536 42073 21539
rect 42024 21508 42073 21536
rect 42024 21496 42030 21508
rect 42061 21505 42073 21508
rect 42107 21505 42119 21539
rect 42061 21499 42119 21505
rect 42702 21496 42708 21548
rect 42760 21536 42766 21548
rect 42889 21539 42947 21545
rect 42889 21536 42901 21539
rect 42760 21508 42901 21536
rect 42760 21496 42766 21508
rect 42889 21505 42901 21508
rect 42935 21505 42947 21539
rect 42889 21499 42947 21505
rect 37844 21440 39068 21468
rect 37844 21412 37872 21440
rect 37826 21360 37832 21412
rect 37884 21360 37890 21412
rect 38013 21403 38071 21409
rect 38013 21369 38025 21403
rect 38059 21400 38071 21403
rect 40310 21400 40316 21412
rect 38059 21372 40316 21400
rect 38059 21369 38071 21372
rect 38013 21363 38071 21369
rect 40310 21360 40316 21372
rect 40368 21360 40374 21412
rect 33704 21304 34468 21332
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 35161 21335 35219 21341
rect 35161 21332 35173 21335
rect 34572 21304 35173 21332
rect 34572 21292 34578 21304
rect 35161 21301 35173 21304
rect 35207 21301 35219 21335
rect 35161 21295 35219 21301
rect 36722 21292 36728 21344
rect 36780 21332 36786 21344
rect 38378 21332 38384 21344
rect 36780 21304 38384 21332
rect 36780 21292 36786 21304
rect 38378 21292 38384 21304
rect 38436 21292 38442 21344
rect 39301 21335 39359 21341
rect 39301 21301 39313 21335
rect 39347 21332 39359 21335
rect 39390 21332 39396 21344
rect 39347 21304 39396 21332
rect 39347 21301 39359 21304
rect 39301 21295 39359 21301
rect 39390 21292 39396 21304
rect 39448 21292 39454 21344
rect 1104 21242 43884 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 43884 21242
rect 1104 21168 43884 21190
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 16758 21128 16764 21140
rect 13412 21100 16764 21128
rect 13412 21088 13418 21100
rect 16758 21088 16764 21100
rect 16816 21088 16822 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 17126 21128 17132 21140
rect 16991 21100 17132 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 18414 21088 18420 21140
rect 18472 21128 18478 21140
rect 24762 21128 24768 21140
rect 18472 21100 24768 21128
rect 18472 21088 18478 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 25004 21100 25084 21128
rect 25004 21088 25010 21100
rect 14642 21020 14648 21072
rect 14700 21060 14706 21072
rect 16666 21060 16672 21072
rect 14700 21032 16672 21060
rect 14700 21020 14706 21032
rect 16666 21020 16672 21032
rect 16724 21020 16730 21072
rect 19334 21020 19340 21072
rect 19392 21060 19398 21072
rect 19521 21063 19579 21069
rect 19521 21060 19533 21063
rect 19392 21032 19533 21060
rect 19392 21020 19398 21032
rect 19521 21029 19533 21032
rect 19567 21029 19579 21063
rect 19521 21023 19579 21029
rect 20898 21020 20904 21072
rect 20956 21060 20962 21072
rect 20993 21063 21051 21069
rect 20993 21060 21005 21063
rect 20956 21032 21005 21060
rect 20956 21020 20962 21032
rect 20993 21029 21005 21032
rect 21039 21029 21051 21063
rect 25056 21060 25084 21100
rect 25130 21088 25136 21140
rect 25188 21088 25194 21140
rect 25682 21088 25688 21140
rect 25740 21088 25746 21140
rect 28994 21088 29000 21140
rect 29052 21128 29058 21140
rect 29730 21128 29736 21140
rect 29052 21100 29736 21128
rect 29052 21088 29058 21100
rect 29730 21088 29736 21100
rect 29788 21088 29794 21140
rect 30101 21131 30159 21137
rect 30101 21097 30113 21131
rect 30147 21128 30159 21131
rect 30374 21128 30380 21140
rect 30147 21100 30380 21128
rect 30147 21097 30159 21100
rect 30101 21091 30159 21097
rect 30374 21088 30380 21100
rect 30432 21088 30438 21140
rect 32214 21088 32220 21140
rect 32272 21128 32278 21140
rect 32272 21100 38332 21128
rect 32272 21088 32278 21100
rect 25056 21032 25912 21060
rect 20993 21023 21051 21029
rect 25884 21004 25912 21032
rect 27430 21020 27436 21072
rect 27488 21060 27494 21072
rect 27525 21063 27583 21069
rect 27525 21060 27537 21063
rect 27488 21032 27537 21060
rect 27488 21020 27494 21032
rect 27525 21029 27537 21032
rect 27571 21029 27583 21063
rect 27525 21023 27583 21029
rect 27798 21020 27804 21072
rect 27856 21060 27862 21072
rect 29362 21060 29368 21072
rect 27856 21032 29368 21060
rect 27856 21020 27862 21032
rect 29362 21020 29368 21032
rect 29420 21020 29426 21072
rect 29454 21020 29460 21072
rect 29512 21060 29518 21072
rect 30282 21060 30288 21072
rect 29512 21032 30288 21060
rect 29512 21020 29518 21032
rect 30282 21020 30288 21032
rect 30340 21020 30346 21072
rect 31570 21060 31576 21072
rect 31312 21032 31576 21060
rect 16025 20995 16083 21001
rect 16025 20992 16037 20995
rect 15212 20964 16037 20992
rect 15212 20936 15240 20964
rect 16025 20961 16037 20964
rect 16071 20992 16083 20995
rect 16071 20964 16436 20992
rect 16071 20961 16083 20964
rect 16025 20955 16083 20961
rect 11974 20884 11980 20936
rect 12032 20884 12038 20936
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 13262 20924 13268 20936
rect 12299 20896 13268 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 14918 20884 14924 20936
rect 14976 20884 14982 20936
rect 15013 20927 15071 20933
rect 15013 20893 15025 20927
rect 15059 20924 15071 20927
rect 15102 20924 15108 20936
rect 15059 20896 15108 20924
rect 15059 20893 15071 20896
rect 15013 20887 15071 20893
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 15286 20884 15292 20936
rect 15344 20924 15350 20936
rect 16114 20924 16120 20936
rect 15344 20896 16120 20924
rect 15344 20884 15350 20896
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 16206 20884 16212 20936
rect 16264 20884 16270 20936
rect 16408 20856 16436 20964
rect 17126 20952 17132 21004
rect 17184 20952 17190 21004
rect 19429 20995 19487 21001
rect 19429 20992 19441 20995
rect 17236 20964 19441 20992
rect 17236 20933 17264 20964
rect 19429 20961 19441 20964
rect 19475 20961 19487 20995
rect 19429 20955 19487 20961
rect 21450 20952 21456 21004
rect 21508 20992 21514 21004
rect 21545 20995 21603 21001
rect 21545 20992 21557 20995
rect 21508 20964 21557 20992
rect 21508 20952 21514 20964
rect 21545 20961 21557 20964
rect 21591 20961 21603 20995
rect 21545 20955 21603 20961
rect 25866 20952 25872 21004
rect 25924 20992 25930 21004
rect 31205 20995 31263 21001
rect 31205 20992 31217 20995
rect 25924 20964 31217 20992
rect 25924 20952 25930 20964
rect 31205 20961 31217 20964
rect 31251 20961 31263 20995
rect 31205 20955 31263 20961
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20893 17279 20927
rect 17221 20887 17279 20893
rect 21266 20884 21272 20936
rect 21324 20884 21330 20936
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22244 20896 22845 20924
rect 22244 20884 22250 20896
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 23017 20927 23075 20933
rect 23017 20893 23029 20927
rect 23063 20924 23075 20927
rect 23382 20924 23388 20936
rect 23063 20896 23388 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 19889 20859 19947 20865
rect 16408 20828 19334 20856
rect 14734 20748 14740 20800
rect 14792 20748 14798 20800
rect 19306 20788 19334 20828
rect 19889 20825 19901 20859
rect 19935 20856 19947 20859
rect 20162 20856 20168 20868
rect 19935 20828 20168 20856
rect 19935 20825 19947 20828
rect 19889 20819 19947 20825
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 24596 20856 24624 20887
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 24949 20927 25007 20933
rect 24949 20924 24961 20927
rect 24912 20896 24961 20924
rect 24912 20884 24918 20896
rect 24949 20893 24961 20896
rect 24995 20924 25007 20927
rect 25222 20924 25228 20936
rect 24995 20896 25228 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 25593 20927 25651 20933
rect 25593 20924 25605 20927
rect 25372 20896 25605 20924
rect 25372 20884 25378 20896
rect 25593 20893 25605 20896
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 25777 20927 25835 20933
rect 25777 20893 25789 20927
rect 25823 20924 25835 20927
rect 26970 20924 26976 20936
rect 25823 20896 26976 20924
rect 25823 20893 25835 20896
rect 25777 20887 25835 20893
rect 25792 20856 25820 20887
rect 26970 20884 26976 20896
rect 27028 20884 27034 20936
rect 27080 20896 28212 20924
rect 22848 20828 25820 20856
rect 22848 20800 22876 20828
rect 25866 20816 25872 20868
rect 25924 20856 25930 20868
rect 27080 20856 27108 20896
rect 27798 20856 27804 20868
rect 25924 20828 27108 20856
rect 27172 20828 27804 20856
rect 25924 20816 25930 20828
rect 20622 20788 20628 20800
rect 19306 20760 20628 20788
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 21453 20791 21511 20797
rect 21453 20788 21465 20791
rect 21416 20760 21465 20788
rect 21416 20748 21422 20760
rect 21453 20757 21465 20760
rect 21499 20757 21511 20791
rect 21453 20751 21511 20757
rect 22830 20748 22836 20800
rect 22888 20748 22894 20800
rect 22925 20791 22983 20797
rect 22925 20757 22937 20791
rect 22971 20788 22983 20791
rect 23290 20788 23296 20800
rect 22971 20760 23296 20788
rect 22971 20757 22983 20760
rect 22925 20751 22983 20757
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 27172 20788 27200 20828
rect 27798 20816 27804 20828
rect 27856 20816 27862 20868
rect 28074 20816 28080 20868
rect 28132 20816 28138 20868
rect 28184 20856 28212 20896
rect 29638 20884 29644 20936
rect 29696 20924 29702 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29696 20896 29745 20924
rect 29696 20884 29702 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 29917 20927 29975 20933
rect 29917 20893 29929 20927
rect 29963 20924 29975 20927
rect 30006 20924 30012 20936
rect 29963 20896 30012 20924
rect 29963 20893 29975 20896
rect 29917 20887 29975 20893
rect 30006 20884 30012 20896
rect 30064 20924 30070 20936
rect 31312 20924 31340 21032
rect 31570 21020 31576 21032
rect 31628 21020 31634 21072
rect 36722 21060 36728 21072
rect 34992 21032 36728 21060
rect 31389 20995 31447 21001
rect 31389 20961 31401 20995
rect 31435 20992 31447 20995
rect 31846 20992 31852 21004
rect 31435 20964 31852 20992
rect 31435 20961 31447 20964
rect 31389 20955 31447 20961
rect 31846 20952 31852 20964
rect 31904 20952 31910 21004
rect 32398 20952 32404 21004
rect 32456 20952 32462 21004
rect 32585 20995 32643 21001
rect 32585 20961 32597 20995
rect 32631 20992 32643 20995
rect 33594 20992 33600 21004
rect 32631 20964 33600 20992
rect 32631 20961 32643 20964
rect 32585 20955 32643 20961
rect 33594 20952 33600 20964
rect 33652 20952 33658 21004
rect 34422 20992 34428 21004
rect 33980 20964 34428 20992
rect 30064 20896 31340 20924
rect 30064 20884 30070 20896
rect 31570 20884 31576 20936
rect 31628 20884 31634 20936
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20924 31723 20927
rect 31754 20924 31760 20936
rect 31711 20896 31760 20924
rect 31711 20893 31723 20896
rect 31665 20887 31723 20893
rect 31754 20884 31760 20896
rect 31812 20924 31818 20936
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 31812 20896 32689 20924
rect 31812 20884 31818 20896
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 33686 20884 33692 20936
rect 33744 20924 33750 20936
rect 33781 20927 33839 20933
rect 33781 20924 33793 20927
rect 33744 20896 33793 20924
rect 33744 20884 33750 20896
rect 33781 20893 33793 20896
rect 33827 20893 33839 20927
rect 33781 20887 33839 20893
rect 32217 20859 32275 20865
rect 32217 20856 32229 20859
rect 28184 20828 32229 20856
rect 32217 20825 32229 20828
rect 32263 20825 32275 20859
rect 32217 20819 32275 20825
rect 33870 20816 33876 20868
rect 33928 20856 33934 20868
rect 33980 20865 34008 20964
rect 34422 20952 34428 20964
rect 34480 20952 34486 21004
rect 34146 20884 34152 20936
rect 34204 20884 34210 20936
rect 34992 20924 35020 21032
rect 36722 21020 36728 21032
rect 36780 21020 36786 21072
rect 36538 20952 36544 21004
rect 36596 20992 36602 21004
rect 37093 20995 37151 21001
rect 37093 20992 37105 20995
rect 36596 20964 37105 20992
rect 36596 20952 36602 20964
rect 37093 20961 37105 20964
rect 37139 20961 37151 20995
rect 37093 20955 37151 20961
rect 37826 20952 37832 21004
rect 37884 20952 37890 21004
rect 34624 20896 35020 20924
rect 35069 20927 35127 20933
rect 33965 20859 34023 20865
rect 33965 20856 33977 20859
rect 33928 20828 33977 20856
rect 33928 20816 33934 20828
rect 33965 20825 33977 20828
rect 34011 20825 34023 20859
rect 33965 20819 34023 20825
rect 34057 20859 34115 20865
rect 34057 20825 34069 20859
rect 34103 20856 34115 20859
rect 34624 20856 34652 20896
rect 35069 20893 35081 20927
rect 35115 20924 35127 20927
rect 35115 20896 35388 20924
rect 35115 20893 35127 20896
rect 35069 20887 35127 20893
rect 34103 20828 34652 20856
rect 34103 20825 34115 20828
rect 34057 20819 34115 20825
rect 24820 20760 27200 20788
rect 24820 20748 24826 20760
rect 27522 20748 27528 20800
rect 27580 20788 27586 20800
rect 27985 20791 28043 20797
rect 27985 20788 27997 20791
rect 27580 20760 27997 20788
rect 27580 20748 27586 20760
rect 27985 20757 27997 20760
rect 28031 20788 28043 20791
rect 29914 20788 29920 20800
rect 28031 20760 29920 20788
rect 28031 20757 28043 20760
rect 27985 20751 28043 20757
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 30282 20748 30288 20800
rect 30340 20788 30346 20800
rect 34072 20788 34100 20819
rect 34698 20816 34704 20868
rect 34756 20856 34762 20868
rect 35161 20859 35219 20865
rect 35161 20856 35173 20859
rect 34756 20828 35173 20856
rect 34756 20816 34762 20828
rect 35161 20825 35173 20828
rect 35207 20825 35219 20859
rect 35161 20819 35219 20825
rect 35253 20859 35311 20865
rect 35253 20825 35265 20859
rect 35299 20825 35311 20859
rect 35360 20856 35388 20896
rect 35434 20884 35440 20936
rect 35492 20884 35498 20936
rect 37001 20927 37059 20933
rect 36648 20896 36952 20924
rect 36648 20865 36676 20896
rect 36633 20859 36691 20865
rect 36633 20856 36645 20859
rect 35360 20828 36645 20856
rect 35253 20819 35311 20825
rect 36633 20825 36645 20828
rect 36679 20825 36691 20859
rect 36633 20819 36691 20825
rect 30340 20760 34100 20788
rect 34333 20791 34391 20797
rect 30340 20748 30346 20760
rect 34333 20757 34345 20791
rect 34379 20788 34391 20791
rect 34790 20788 34796 20800
rect 34379 20760 34796 20788
rect 34379 20757 34391 20760
rect 34333 20751 34391 20757
rect 34790 20748 34796 20760
rect 34848 20748 34854 20800
rect 34882 20748 34888 20800
rect 34940 20748 34946 20800
rect 35268 20788 35296 20819
rect 36722 20816 36728 20868
rect 36780 20816 36786 20868
rect 36924 20856 36952 20896
rect 37001 20893 37013 20927
rect 37047 20924 37059 20927
rect 37182 20924 37188 20936
rect 37047 20896 37188 20924
rect 37047 20893 37059 20896
rect 37001 20887 37059 20893
rect 37182 20884 37188 20896
rect 37240 20924 37246 20936
rect 38105 20927 38163 20933
rect 38105 20924 38117 20927
rect 37240 20896 38117 20924
rect 37240 20884 37246 20896
rect 38105 20893 38117 20896
rect 38151 20893 38163 20927
rect 38105 20887 38163 20893
rect 38194 20884 38200 20936
rect 38252 20884 38258 20936
rect 38304 20924 38332 21100
rect 40586 21088 40592 21140
rect 40644 21088 40650 21140
rect 38381 21063 38439 21069
rect 38381 21029 38393 21063
rect 38427 21060 38439 21063
rect 40402 21060 40408 21072
rect 38427 21032 40408 21060
rect 38427 21029 38439 21032
rect 38381 21023 38439 21029
rect 40402 21020 40408 21032
rect 40460 21020 40466 21072
rect 38841 20995 38899 21001
rect 38841 20961 38853 20995
rect 38887 20992 38899 20995
rect 39298 20992 39304 21004
rect 38887 20964 39304 20992
rect 38887 20961 38899 20964
rect 38841 20955 38899 20961
rect 39298 20952 39304 20964
rect 39356 20952 39362 21004
rect 39390 20952 39396 21004
rect 39448 20952 39454 21004
rect 40126 20952 40132 21004
rect 40184 20952 40190 21004
rect 43165 20995 43223 21001
rect 43165 20961 43177 20995
rect 43211 20992 43223 20995
rect 43254 20992 43260 21004
rect 43211 20964 43260 20992
rect 43211 20961 43223 20964
rect 43165 20955 43223 20961
rect 43254 20952 43260 20964
rect 43312 20952 43318 21004
rect 39025 20927 39083 20933
rect 39025 20924 39037 20927
rect 38304 20896 39037 20924
rect 39025 20893 39037 20896
rect 39071 20893 39083 20927
rect 39025 20887 39083 20893
rect 37550 20856 37556 20868
rect 36924 20828 37556 20856
rect 37550 20816 37556 20828
rect 37608 20856 37614 20868
rect 37737 20859 37795 20865
rect 37737 20856 37749 20859
rect 37608 20828 37749 20856
rect 37608 20816 37614 20828
rect 37737 20825 37749 20828
rect 37783 20825 37795 20859
rect 39040 20856 39068 20887
rect 39758 20884 39764 20936
rect 39816 20924 39822 20936
rect 40221 20927 40279 20933
rect 40221 20924 40233 20927
rect 39816 20896 40233 20924
rect 39816 20884 39822 20896
rect 40221 20893 40233 20896
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 40126 20856 40132 20868
rect 39040 20828 40132 20856
rect 37737 20819 37795 20825
rect 40126 20816 40132 20828
rect 40184 20816 40190 20868
rect 42702 20816 42708 20868
rect 42760 20856 42766 20868
rect 42981 20859 43039 20865
rect 42981 20856 42993 20859
rect 42760 20828 42993 20856
rect 42760 20816 42766 20828
rect 42981 20825 42993 20828
rect 43027 20825 43039 20859
rect 42981 20819 43039 20825
rect 37182 20788 37188 20800
rect 35268 20760 37188 20788
rect 37182 20748 37188 20760
rect 37240 20748 37246 20800
rect 37277 20791 37335 20797
rect 37277 20757 37289 20791
rect 37323 20788 37335 20791
rect 37642 20788 37648 20800
rect 37323 20760 37648 20788
rect 37323 20757 37335 20760
rect 37277 20751 37335 20757
rect 37642 20748 37648 20760
rect 37700 20748 37706 20800
rect 39298 20748 39304 20800
rect 39356 20748 39362 20800
rect 42518 20748 42524 20800
rect 42576 20748 42582 20800
rect 42794 20748 42800 20800
rect 42852 20788 42858 20800
rect 42889 20791 42947 20797
rect 42889 20788 42901 20791
rect 42852 20760 42901 20788
rect 42852 20748 42858 20760
rect 42889 20757 42901 20760
rect 42935 20757 42947 20791
rect 42889 20751 42947 20757
rect 1104 20698 43884 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 43884 20698
rect 1104 20624 43884 20646
rect 13262 20544 13268 20596
rect 13320 20584 13326 20596
rect 13909 20587 13967 20593
rect 13909 20584 13921 20587
rect 13320 20556 13921 20584
rect 13320 20544 13326 20556
rect 13909 20553 13921 20556
rect 13955 20553 13967 20587
rect 13909 20547 13967 20553
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14734 20584 14740 20596
rect 14323 20556 14740 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 17126 20544 17132 20596
rect 17184 20584 17190 20596
rect 17681 20587 17739 20593
rect 17681 20584 17693 20587
rect 17184 20556 17693 20584
rect 17184 20544 17190 20556
rect 17681 20553 17693 20556
rect 17727 20553 17739 20587
rect 17681 20547 17739 20553
rect 27890 20544 27896 20596
rect 27948 20584 27954 20596
rect 28718 20584 28724 20596
rect 27948 20556 28724 20584
rect 27948 20544 27954 20556
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 29914 20544 29920 20596
rect 29972 20584 29978 20596
rect 30374 20584 30380 20596
rect 29972 20556 30047 20584
rect 29972 20544 29978 20556
rect 14829 20519 14887 20525
rect 14829 20516 14841 20519
rect 14384 20488 14841 20516
rect 14090 20408 14096 20460
rect 14148 20408 14154 20460
rect 14384 20457 14412 20488
rect 14829 20485 14841 20488
rect 14875 20485 14887 20519
rect 18785 20519 18843 20525
rect 14829 20479 14887 20485
rect 17696 20488 18000 20516
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20448 15071 20451
rect 15102 20448 15108 20460
rect 15059 20420 15108 20448
rect 15059 20417 15071 20420
rect 15013 20411 15071 20417
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 17696 20457 17724 20488
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 15252 20420 15301 20448
rect 15252 20408 15258 20420
rect 15289 20417 15301 20420
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17972 20448 18000 20488
rect 18785 20485 18797 20519
rect 18831 20516 18843 20519
rect 20162 20516 20168 20528
rect 18831 20488 20168 20516
rect 18831 20485 18843 20488
rect 18785 20479 18843 20485
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 22738 20516 22744 20528
rect 20640 20488 22744 20516
rect 18874 20448 18880 20460
rect 17972 20420 18880 20448
rect 17865 20411 17923 20417
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 14918 20380 14924 20392
rect 14608 20352 14924 20380
rect 14608 20340 14614 20352
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 17880 20380 17908 20411
rect 18874 20408 18880 20420
rect 18932 20448 18938 20460
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 18932 20420 19165 20448
rect 18932 20408 18938 20420
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 18138 20380 18144 20392
rect 17880 20352 18144 20380
rect 18138 20340 18144 20352
rect 18196 20380 18202 20392
rect 19061 20383 19119 20389
rect 19061 20380 19073 20383
rect 18196 20352 19073 20380
rect 18196 20340 18202 20352
rect 19061 20349 19073 20352
rect 19107 20349 19119 20383
rect 19260 20380 19288 20411
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 20128 20420 20269 20448
rect 20128 20408 20134 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20346 20408 20352 20460
rect 20404 20448 20410 20460
rect 20640 20457 20668 20488
rect 22738 20476 22744 20488
rect 22796 20476 22802 20528
rect 23293 20519 23351 20525
rect 23293 20485 23305 20519
rect 23339 20516 23351 20519
rect 24210 20516 24216 20528
rect 23339 20488 24216 20516
rect 23339 20485 23351 20488
rect 23293 20479 23351 20485
rect 24210 20476 24216 20488
rect 24268 20476 24274 20528
rect 27525 20519 27583 20525
rect 27525 20485 27537 20519
rect 27571 20516 27583 20519
rect 27571 20488 29960 20516
rect 27571 20485 27583 20488
rect 27525 20479 27583 20485
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20404 20420 20637 20448
rect 20404 20408 20410 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 20898 20408 20904 20460
rect 20956 20408 20962 20460
rect 21361 20451 21419 20457
rect 21361 20417 21373 20451
rect 21407 20448 21419 20451
rect 22094 20448 22100 20460
rect 21407 20420 22100 20448
rect 21407 20417 21419 20420
rect 21361 20411 21419 20417
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22704 20420 23121 20448
rect 22704 20408 22710 20420
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 23934 20448 23940 20460
rect 23431 20420 23940 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 19334 20380 19340 20392
rect 19260 20352 19340 20380
rect 19061 20343 19119 20349
rect 19334 20340 19340 20352
rect 19392 20380 19398 20392
rect 19981 20383 20039 20389
rect 19981 20380 19993 20383
rect 19392 20352 19993 20380
rect 19392 20340 19398 20352
rect 19981 20349 19993 20352
rect 20027 20349 20039 20383
rect 23124 20380 23152 20411
rect 23934 20408 23940 20420
rect 23992 20408 23998 20460
rect 24854 20408 24860 20460
rect 24912 20408 24918 20460
rect 25041 20451 25099 20457
rect 25041 20417 25053 20451
rect 25087 20448 25099 20451
rect 25682 20448 25688 20460
rect 25087 20420 25688 20448
rect 25087 20417 25099 20420
rect 25041 20411 25099 20417
rect 25682 20408 25688 20420
rect 25740 20448 25746 20460
rect 26050 20448 26056 20460
rect 25740 20420 26056 20448
rect 25740 20408 25746 20420
rect 26050 20408 26056 20420
rect 26108 20408 26114 20460
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27381 20451 27439 20457
rect 27381 20448 27393 20451
rect 27120 20420 27393 20448
rect 27120 20408 27126 20420
rect 27381 20417 27393 20420
rect 27427 20417 27439 20451
rect 27381 20411 27439 20417
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20417 27675 20451
rect 27617 20411 27675 20417
rect 25314 20380 25320 20392
rect 23124 20352 25320 20380
rect 19981 20343 20039 20349
rect 25314 20340 25320 20352
rect 25372 20340 25378 20392
rect 27632 20380 27660 20411
rect 27798 20408 27804 20460
rect 27856 20408 27862 20460
rect 28534 20457 28540 20460
rect 28532 20448 28540 20457
rect 28495 20420 28540 20448
rect 28532 20411 28540 20420
rect 28534 20408 28540 20411
rect 28592 20408 28598 20460
rect 28629 20451 28687 20457
rect 28629 20417 28641 20451
rect 28675 20417 28687 20451
rect 28629 20411 28687 20417
rect 27890 20380 27896 20392
rect 27632 20352 27896 20380
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 15197 20315 15255 20321
rect 15197 20281 15209 20315
rect 15243 20312 15255 20315
rect 15286 20312 15292 20324
rect 15243 20284 15292 20312
rect 15243 20281 15255 20284
rect 15197 20275 15255 20281
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 18506 20272 18512 20324
rect 18564 20272 18570 20324
rect 23382 20272 23388 20324
rect 23440 20312 23446 20324
rect 24026 20312 24032 20324
rect 23440 20284 24032 20312
rect 23440 20272 23446 20284
rect 24026 20272 24032 20284
rect 24084 20312 24090 20324
rect 28644 20312 28672 20411
rect 28718 20408 28724 20460
rect 28776 20408 28782 20460
rect 28902 20408 28908 20460
rect 28960 20408 28966 20460
rect 29932 20380 29960 20488
rect 30019 20457 30047 20556
rect 30208 20556 30380 20584
rect 30098 20476 30104 20528
rect 30156 20476 30162 20528
rect 30208 20525 30236 20556
rect 30374 20544 30380 20556
rect 30432 20544 30438 20596
rect 34054 20544 34060 20596
rect 34112 20584 34118 20596
rect 34112 20556 35756 20584
rect 34112 20544 34118 20556
rect 30193 20519 30251 20525
rect 30193 20485 30205 20519
rect 30239 20485 30251 20519
rect 34882 20516 34888 20528
rect 30193 20479 30251 20485
rect 34440 20488 34888 20516
rect 30004 20451 30062 20457
rect 30004 20417 30016 20451
rect 30050 20417 30062 20451
rect 30004 20411 30062 20417
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20448 30435 20451
rect 30650 20448 30656 20460
rect 30423 20420 30656 20448
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 30650 20408 30656 20420
rect 30708 20408 30714 20460
rect 34149 20451 34207 20457
rect 34149 20417 34161 20451
rect 34195 20417 34207 20451
rect 34149 20411 34207 20417
rect 33686 20380 33692 20392
rect 29932 20352 33692 20380
rect 33686 20340 33692 20352
rect 33744 20340 33750 20392
rect 34164 20312 34192 20411
rect 34238 20408 34244 20460
rect 34296 20408 34302 20460
rect 34440 20457 34468 20488
rect 34882 20476 34888 20488
rect 34940 20476 34946 20528
rect 35342 20476 35348 20528
rect 35400 20476 35406 20528
rect 34425 20451 34483 20457
rect 34425 20417 34437 20451
rect 34471 20417 34483 20451
rect 34425 20411 34483 20417
rect 34514 20408 34520 20460
rect 34572 20408 34578 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 34977 20451 35035 20457
rect 34977 20448 34989 20451
rect 34848 20420 34989 20448
rect 34848 20408 34854 20420
rect 34977 20417 34989 20420
rect 35023 20417 35035 20451
rect 34977 20411 35035 20417
rect 35250 20408 35256 20460
rect 35308 20408 35314 20460
rect 35728 20457 35756 20556
rect 39022 20544 39028 20596
rect 39080 20584 39086 20596
rect 39669 20587 39727 20593
rect 39080 20556 39344 20584
rect 39080 20544 39086 20556
rect 39316 20525 39344 20556
rect 39669 20553 39681 20587
rect 39715 20553 39727 20587
rect 39669 20547 39727 20553
rect 40681 20587 40739 20593
rect 40681 20553 40693 20587
rect 40727 20584 40739 20587
rect 42702 20584 42708 20596
rect 40727 20556 42708 20584
rect 40727 20553 40739 20556
rect 40681 20547 40739 20553
rect 39301 20519 39359 20525
rect 39301 20485 39313 20519
rect 39347 20485 39359 20519
rect 39684 20516 39712 20547
rect 42702 20544 42708 20556
rect 42760 20544 42766 20596
rect 39684 20488 40540 20516
rect 39301 20479 39359 20485
rect 35529 20451 35587 20457
rect 35529 20417 35541 20451
rect 35575 20417 35587 20451
rect 35529 20411 35587 20417
rect 35713 20451 35771 20457
rect 35713 20417 35725 20451
rect 35759 20417 35771 20451
rect 35713 20411 35771 20417
rect 35544 20312 35572 20411
rect 38838 20408 38844 20460
rect 38896 20448 38902 20460
rect 39025 20451 39083 20457
rect 39025 20448 39037 20451
rect 38896 20420 39037 20448
rect 38896 20408 38902 20420
rect 39025 20417 39037 20420
rect 39071 20417 39083 20451
rect 39025 20411 39083 20417
rect 39114 20408 39120 20460
rect 39172 20408 39178 20460
rect 39393 20451 39451 20457
rect 39393 20417 39405 20451
rect 39439 20417 39451 20451
rect 39393 20411 39451 20417
rect 37366 20340 37372 20392
rect 37424 20380 37430 20392
rect 37734 20380 37740 20392
rect 37424 20352 37740 20380
rect 37424 20340 37430 20352
rect 37734 20340 37740 20352
rect 37792 20340 37798 20392
rect 38746 20340 38752 20392
rect 38804 20380 38810 20392
rect 39408 20380 39436 20411
rect 39482 20408 39488 20460
rect 39540 20457 39546 20460
rect 39540 20448 39548 20457
rect 39540 20420 39585 20448
rect 39540 20411 39548 20420
rect 39540 20408 39546 20411
rect 40126 20408 40132 20460
rect 40184 20408 40190 20460
rect 40402 20408 40408 20460
rect 40460 20408 40466 20460
rect 40512 20457 40540 20488
rect 40497 20451 40555 20457
rect 40497 20417 40509 20451
rect 40543 20417 40555 20451
rect 40497 20411 40555 20417
rect 42702 20408 42708 20460
rect 42760 20448 42766 20460
rect 42889 20451 42947 20457
rect 42889 20448 42901 20451
rect 42760 20420 42901 20448
rect 42760 20408 42766 20420
rect 42889 20417 42901 20420
rect 42935 20417 42947 20451
rect 42889 20411 42947 20417
rect 42794 20380 42800 20392
rect 38804 20352 42800 20380
rect 38804 20340 38810 20352
rect 42794 20340 42800 20352
rect 42852 20340 42858 20392
rect 43162 20340 43168 20392
rect 43220 20340 43226 20392
rect 37458 20312 37464 20324
rect 24084 20284 27384 20312
rect 28644 20284 31754 20312
rect 34164 20284 35480 20312
rect 35544 20284 37464 20312
rect 24084 20272 24090 20284
rect 22925 20247 22983 20253
rect 22925 20213 22937 20247
rect 22971 20244 22983 20247
rect 23014 20244 23020 20256
rect 22971 20216 23020 20244
rect 22971 20213 22983 20216
rect 22925 20207 22983 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 24946 20204 24952 20256
rect 25004 20244 25010 20256
rect 25041 20247 25099 20253
rect 25041 20244 25053 20247
rect 25004 20216 25053 20244
rect 25004 20204 25010 20216
rect 25041 20213 25053 20216
rect 25087 20213 25099 20247
rect 25041 20207 25099 20213
rect 27246 20204 27252 20256
rect 27304 20204 27310 20256
rect 27356 20244 27384 20284
rect 28353 20247 28411 20253
rect 28353 20244 28365 20247
rect 27356 20216 28365 20244
rect 28353 20213 28365 20216
rect 28399 20213 28411 20247
rect 28353 20207 28411 20213
rect 29822 20204 29828 20256
rect 29880 20204 29886 20256
rect 31726 20244 31754 20284
rect 32214 20244 32220 20256
rect 31726 20216 32220 20244
rect 32214 20204 32220 20216
rect 32272 20204 32278 20256
rect 33965 20247 34023 20253
rect 33965 20213 33977 20247
rect 34011 20244 34023 20247
rect 34698 20244 34704 20256
rect 34011 20216 34704 20244
rect 34011 20213 34023 20216
rect 33965 20207 34023 20213
rect 34698 20204 34704 20216
rect 34756 20204 34762 20256
rect 35452 20244 35480 20284
rect 37458 20272 37464 20284
rect 37516 20312 37522 20324
rect 42978 20312 42984 20324
rect 37516 20284 42984 20312
rect 37516 20272 37522 20284
rect 42978 20272 42984 20284
rect 43036 20272 43042 20324
rect 37550 20244 37556 20256
rect 35452 20216 37556 20244
rect 37550 20204 37556 20216
rect 37608 20204 37614 20256
rect 40126 20204 40132 20256
rect 40184 20244 40190 20256
rect 40221 20247 40279 20253
rect 40221 20244 40233 20247
rect 40184 20216 40233 20244
rect 40184 20204 40190 20216
rect 40221 20213 40233 20216
rect 40267 20213 40279 20247
rect 40221 20207 40279 20213
rect 1104 20154 43884 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 43884 20154
rect 1104 20080 43884 20102
rect 14090 20000 14096 20052
rect 14148 20040 14154 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14148 20012 14657 20040
rect 14148 20000 14154 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 15289 20043 15347 20049
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 15378 20040 15384 20052
rect 15335 20012 15384 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 18138 20000 18144 20052
rect 18196 20000 18202 20052
rect 23201 20043 23259 20049
rect 23201 20009 23213 20043
rect 23247 20040 23259 20043
rect 24854 20040 24860 20052
rect 23247 20012 24860 20040
rect 23247 20009 23259 20012
rect 23201 20003 23259 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 28350 20000 28356 20052
rect 28408 20040 28414 20052
rect 29454 20040 29460 20052
rect 28408 20012 29460 20040
rect 28408 20000 28414 20012
rect 18322 19972 18328 19984
rect 17972 19944 18328 19972
rect 15381 19907 15439 19913
rect 15381 19873 15393 19907
rect 15427 19904 15439 19907
rect 15470 19904 15476 19916
rect 15427 19876 15476 19904
rect 15427 19873 15439 19876
rect 15381 19867 15439 19873
rect 15470 19864 15476 19876
rect 15528 19904 15534 19916
rect 16022 19904 16028 19916
rect 15528 19876 16028 19904
rect 15528 19864 15534 19876
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 17972 19845 18000 19944
rect 18322 19932 18328 19944
rect 18380 19972 18386 19984
rect 22646 19972 22652 19984
rect 18380 19944 22652 19972
rect 18380 19932 18386 19944
rect 22646 19932 22652 19944
rect 22704 19932 22710 19984
rect 24670 19972 24676 19984
rect 23768 19944 24676 19972
rect 23768 19916 23796 19944
rect 24670 19932 24676 19944
rect 24728 19932 24734 19984
rect 24762 19932 24768 19984
rect 24820 19972 24826 19984
rect 25225 19975 25283 19981
rect 25225 19972 25237 19975
rect 24820 19944 25237 19972
rect 24820 19932 24826 19944
rect 25225 19941 25237 19944
rect 25271 19941 25283 19975
rect 25225 19935 25283 19941
rect 19981 19907 20039 19913
rect 19981 19873 19993 19907
rect 20027 19904 20039 19907
rect 20346 19904 20352 19916
rect 20027 19876 20352 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 20898 19904 20904 19916
rect 20579 19876 20904 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 23750 19864 23756 19916
rect 23808 19864 23814 19916
rect 25038 19904 25044 19916
rect 23860 19876 25044 19904
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 14884 19808 14933 19836
rect 14884 19796 14890 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 18414 19836 18420 19848
rect 18187 19808 18420 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 20070 19796 20076 19848
rect 20128 19836 20134 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 20128 19808 20177 19836
rect 20128 19796 20134 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 22922 19796 22928 19848
rect 22980 19796 22986 19848
rect 23014 19796 23020 19848
rect 23072 19796 23078 19848
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19836 23351 19839
rect 23860 19836 23888 19876
rect 25038 19864 25044 19876
rect 25096 19864 25102 19916
rect 27798 19864 27804 19916
rect 27856 19904 27862 19916
rect 27856 19876 28580 19904
rect 27856 19864 27862 19876
rect 23339 19808 23888 19836
rect 23339 19805 23351 19808
rect 23293 19799 23351 19805
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 15105 19771 15163 19777
rect 15105 19768 15117 19771
rect 14608 19740 15117 19768
rect 14608 19728 14614 19740
rect 15105 19737 15117 19740
rect 15151 19737 15163 19771
rect 15105 19731 15163 19737
rect 20622 19728 20628 19780
rect 20680 19768 20686 19780
rect 23308 19768 23336 19799
rect 23934 19796 23940 19848
rect 23992 19796 23998 19848
rect 24029 19839 24087 19845
rect 24029 19805 24041 19839
rect 24075 19836 24087 19839
rect 24210 19836 24216 19848
rect 24075 19808 24216 19836
rect 24075 19805 24087 19808
rect 24029 19799 24087 19805
rect 24210 19796 24216 19808
rect 24268 19836 24274 19848
rect 24854 19836 24860 19848
rect 24268 19808 24860 19836
rect 24268 19796 24274 19808
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 24946 19796 24952 19848
rect 25004 19796 25010 19848
rect 25498 19796 25504 19848
rect 25556 19836 25562 19848
rect 25685 19839 25743 19845
rect 25685 19836 25697 19839
rect 25556 19808 25697 19836
rect 25556 19796 25562 19808
rect 25685 19805 25697 19808
rect 25731 19805 25743 19839
rect 25685 19799 25743 19805
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19836 25927 19839
rect 27246 19836 27252 19848
rect 25915 19808 27252 19836
rect 25915 19805 25927 19808
rect 25869 19799 25927 19805
rect 20680 19740 23336 19768
rect 20680 19728 20686 19740
rect 23382 19728 23388 19780
rect 23440 19768 23446 19780
rect 25041 19771 25099 19777
rect 25041 19768 25053 19771
rect 23440 19740 25053 19768
rect 23440 19728 23446 19740
rect 25041 19737 25053 19740
rect 25087 19737 25099 19771
rect 25041 19731 25099 19737
rect 15013 19703 15071 19709
rect 15013 19669 15025 19703
rect 15059 19700 15071 19703
rect 19426 19700 19432 19712
rect 15059 19672 19432 19700
rect 15059 19669 15071 19672
rect 15013 19663 15071 19669
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 20162 19660 20168 19712
rect 20220 19660 20226 19712
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22741 19703 22799 19709
rect 22741 19700 22753 19703
rect 22612 19672 22753 19700
rect 22612 19660 22618 19672
rect 22741 19669 22753 19672
rect 22787 19669 22799 19703
rect 22741 19663 22799 19669
rect 23106 19660 23112 19712
rect 23164 19700 23170 19712
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23164 19672 23765 19700
rect 23164 19660 23170 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 25056 19700 25084 19731
rect 25222 19728 25228 19780
rect 25280 19728 25286 19780
rect 25884 19768 25912 19799
rect 27246 19796 27252 19808
rect 27304 19796 27310 19848
rect 28074 19845 28080 19848
rect 28057 19839 28080 19845
rect 28057 19805 28069 19839
rect 28057 19799 28080 19805
rect 28074 19796 28080 19799
rect 28132 19796 28138 19848
rect 28166 19796 28172 19848
rect 28224 19796 28230 19848
rect 25700 19740 25912 19768
rect 25700 19700 25728 19740
rect 28442 19728 28448 19780
rect 28500 19728 28506 19780
rect 28552 19777 28580 19876
rect 28828 19836 28856 20012
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 29638 20000 29644 20052
rect 29696 20040 29702 20052
rect 29825 20043 29883 20049
rect 29825 20040 29837 20043
rect 29696 20012 29837 20040
rect 29696 20000 29702 20012
rect 29825 20009 29837 20012
rect 29871 20009 29883 20043
rect 29825 20003 29883 20009
rect 30650 20000 30656 20052
rect 30708 20000 30714 20052
rect 33686 20000 33692 20052
rect 33744 20040 33750 20052
rect 37366 20040 37372 20052
rect 33744 20012 37372 20040
rect 33744 20000 33750 20012
rect 37366 20000 37372 20012
rect 37424 20000 37430 20052
rect 40034 20000 40040 20052
rect 40092 20040 40098 20052
rect 41414 20040 41420 20052
rect 40092 20012 41420 20040
rect 40092 20000 40098 20012
rect 41414 20000 41420 20012
rect 41472 20000 41478 20052
rect 42794 20000 42800 20052
rect 42852 20040 42858 20052
rect 43257 20043 43315 20049
rect 43257 20040 43269 20043
rect 42852 20012 43269 20040
rect 42852 20000 42858 20012
rect 43257 20009 43269 20012
rect 43303 20009 43315 20043
rect 43257 20003 43315 20009
rect 28902 19932 28908 19984
rect 28960 19972 28966 19984
rect 31846 19972 31852 19984
rect 28960 19944 31852 19972
rect 28960 19932 28966 19944
rect 31846 19932 31852 19944
rect 31904 19932 31910 19984
rect 37274 19932 37280 19984
rect 37332 19972 37338 19984
rect 37918 19972 37924 19984
rect 37332 19944 37924 19972
rect 37332 19932 37338 19944
rect 37918 19932 37924 19944
rect 37976 19972 37982 19984
rect 39022 19972 39028 19984
rect 37976 19944 39028 19972
rect 37976 19932 37982 19944
rect 39022 19932 39028 19944
rect 39080 19932 39086 19984
rect 39224 19944 41414 19972
rect 29730 19904 29736 19916
rect 29196 19876 29736 19904
rect 28997 19839 29055 19845
rect 28997 19836 29009 19839
rect 28828 19808 29009 19836
rect 28997 19805 29009 19808
rect 29043 19805 29055 19839
rect 28997 19799 29055 19805
rect 29086 19796 29092 19848
rect 29144 19836 29150 19848
rect 29196 19845 29224 19876
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 29914 19864 29920 19916
rect 29972 19904 29978 19916
rect 31110 19904 31116 19916
rect 29972 19876 31116 19904
rect 29972 19864 29978 19876
rect 29181 19839 29239 19845
rect 29181 19836 29193 19839
rect 29144 19808 29193 19836
rect 29144 19796 29150 19808
rect 29181 19805 29193 19808
rect 29227 19805 29239 19839
rect 29181 19799 29239 19805
rect 29454 19796 29460 19848
rect 29512 19836 29518 19848
rect 30006 19836 30012 19848
rect 29512 19808 30012 19836
rect 29512 19796 29518 19808
rect 30006 19796 30012 19808
rect 30064 19796 30070 19848
rect 30098 19796 30104 19848
rect 30156 19836 30162 19848
rect 30852 19845 30880 19876
rect 31110 19864 31116 19876
rect 31168 19904 31174 19916
rect 39224 19904 39252 19944
rect 31168 19876 32076 19904
rect 31168 19864 31174 19876
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 30156 19808 30205 19836
rect 30156 19796 30162 19808
rect 30193 19805 30205 19808
rect 30239 19836 30251 19839
rect 30653 19839 30711 19845
rect 30653 19836 30665 19839
rect 30239 19808 30665 19836
rect 30239 19805 30251 19808
rect 30193 19799 30251 19805
rect 30653 19805 30665 19808
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19805 30895 19839
rect 30837 19799 30895 19805
rect 31754 19796 31760 19848
rect 31812 19796 31818 19848
rect 31846 19796 31852 19848
rect 31904 19796 31910 19848
rect 32048 19845 32076 19876
rect 34256 19876 39252 19904
rect 33870 19845 33876 19848
rect 32033 19839 32091 19845
rect 32033 19805 32045 19839
rect 32079 19805 32091 19839
rect 32033 19799 32091 19805
rect 33868 19799 33876 19845
rect 33870 19796 33876 19799
rect 33928 19796 33934 19848
rect 34054 19796 34060 19848
rect 34112 19796 34118 19848
rect 34256 19845 34284 19876
rect 34240 19839 34298 19845
rect 34240 19805 34252 19839
rect 34286 19805 34298 19839
rect 34240 19799 34298 19805
rect 34330 19796 34336 19848
rect 34388 19796 34394 19848
rect 36078 19796 36084 19848
rect 36136 19836 36142 19848
rect 37093 19839 37151 19845
rect 37093 19836 37105 19839
rect 36136 19808 37105 19836
rect 36136 19796 36142 19808
rect 37093 19805 37105 19808
rect 37139 19805 37151 19839
rect 37093 19799 37151 19805
rect 28537 19771 28595 19777
rect 28537 19737 28549 19771
rect 28583 19768 28595 19771
rect 30374 19768 30380 19780
rect 28583 19740 30380 19768
rect 28583 19737 28595 19740
rect 28537 19731 28595 19737
rect 30374 19728 30380 19740
rect 30432 19728 30438 19780
rect 32493 19771 32551 19777
rect 32493 19737 32505 19771
rect 32539 19768 32551 19771
rect 32582 19768 32588 19780
rect 32539 19740 32588 19768
rect 32539 19737 32551 19740
rect 32493 19731 32551 19737
rect 32582 19728 32588 19740
rect 32640 19728 32646 19780
rect 33410 19728 33416 19780
rect 33468 19768 33474 19780
rect 33965 19771 34023 19777
rect 33965 19768 33977 19771
rect 33468 19740 33977 19768
rect 33468 19728 33474 19740
rect 33965 19737 33977 19740
rect 34011 19768 34023 19771
rect 34422 19768 34428 19780
rect 34011 19740 34428 19768
rect 34011 19737 34023 19740
rect 33965 19731 34023 19737
rect 34422 19728 34428 19740
rect 34480 19728 34486 19780
rect 25056 19672 25728 19700
rect 25777 19703 25835 19709
rect 23753 19663 23811 19669
rect 25777 19669 25789 19703
rect 25823 19700 25835 19703
rect 26050 19700 26056 19712
rect 25823 19672 26056 19700
rect 25823 19669 25835 19672
rect 25777 19663 25835 19669
rect 26050 19660 26056 19672
rect 26108 19660 26114 19712
rect 27890 19660 27896 19712
rect 27948 19660 27954 19712
rect 28718 19660 28724 19712
rect 28776 19700 28782 19712
rect 28997 19703 29055 19709
rect 28997 19700 29009 19703
rect 28776 19672 29009 19700
rect 28776 19660 28782 19672
rect 28997 19669 29009 19672
rect 29043 19669 29055 19703
rect 28997 19663 29055 19669
rect 33686 19660 33692 19712
rect 33744 19660 33750 19712
rect 37108 19700 37136 19799
rect 37182 19796 37188 19848
rect 37240 19796 37246 19848
rect 37274 19796 37280 19848
rect 37332 19836 37338 19848
rect 37369 19839 37427 19845
rect 37369 19836 37381 19839
rect 37332 19808 37381 19836
rect 37332 19796 37338 19808
rect 37369 19805 37381 19808
rect 37415 19805 37427 19839
rect 37369 19799 37427 19805
rect 37458 19796 37464 19848
rect 37516 19796 37522 19848
rect 37550 19796 37556 19848
rect 37608 19845 37614 19848
rect 37608 19836 37616 19845
rect 38746 19836 38752 19848
rect 37608 19808 38752 19836
rect 37608 19799 37616 19808
rect 37608 19796 37614 19799
rect 38746 19796 38752 19808
rect 38804 19796 38810 19848
rect 38838 19796 38844 19848
rect 38896 19796 38902 19848
rect 38930 19796 38936 19848
rect 38988 19796 38994 19848
rect 39022 19796 39028 19848
rect 39080 19836 39086 19848
rect 39224 19845 39252 19876
rect 40126 19864 40132 19916
rect 40184 19864 40190 19916
rect 39117 19839 39175 19845
rect 39117 19836 39129 19839
rect 39080 19808 39129 19836
rect 39080 19796 39086 19808
rect 39117 19805 39129 19808
rect 39163 19805 39175 19839
rect 39117 19799 39175 19805
rect 39209 19839 39267 19845
rect 39209 19805 39221 19839
rect 39255 19805 39267 19839
rect 39209 19799 39267 19805
rect 39306 19839 39364 19845
rect 39306 19805 39318 19839
rect 39352 19836 39364 19839
rect 39482 19836 39488 19848
rect 39352 19808 39488 19836
rect 39352 19805 39364 19808
rect 39306 19799 39364 19805
rect 38856 19768 38884 19796
rect 37660 19740 38884 19768
rect 37660 19700 37688 19740
rect 37108 19672 37688 19700
rect 37737 19703 37795 19709
rect 37737 19669 37749 19703
rect 37783 19700 37795 19703
rect 37826 19700 37832 19712
rect 37783 19672 37832 19700
rect 37783 19669 37795 19672
rect 37737 19663 37795 19669
rect 37826 19660 37832 19672
rect 37884 19660 37890 19712
rect 38746 19660 38752 19712
rect 38804 19700 38810 19712
rect 39316 19700 39344 19799
rect 39482 19796 39488 19808
rect 39540 19796 39546 19848
rect 39666 19796 39672 19848
rect 39724 19836 39730 19848
rect 40037 19839 40095 19845
rect 40037 19836 40049 19839
rect 39724 19808 40049 19836
rect 39724 19796 39730 19808
rect 40037 19805 40049 19808
rect 40083 19805 40095 19839
rect 40037 19799 40095 19805
rect 40310 19796 40316 19848
rect 40368 19796 40374 19848
rect 40405 19839 40463 19845
rect 40405 19805 40417 19839
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 40420 19768 40448 19799
rect 39500 19740 40448 19768
rect 41386 19768 41414 19944
rect 41506 19796 41512 19848
rect 41564 19836 41570 19848
rect 41877 19839 41935 19845
rect 41877 19836 41889 19839
rect 41564 19808 41889 19836
rect 41564 19796 41570 19808
rect 41877 19805 41889 19808
rect 41923 19805 41935 19839
rect 41877 19799 41935 19805
rect 42144 19839 42202 19845
rect 42144 19805 42156 19839
rect 42190 19836 42202 19839
rect 42518 19836 42524 19848
rect 42190 19808 42524 19836
rect 42190 19805 42202 19808
rect 42144 19799 42202 19805
rect 42518 19796 42524 19808
rect 42576 19796 42582 19848
rect 41598 19768 41604 19780
rect 41386 19740 41604 19768
rect 39500 19709 39528 19740
rect 41598 19728 41604 19740
rect 41656 19728 41662 19780
rect 38804 19672 39344 19700
rect 39485 19703 39543 19709
rect 38804 19660 38810 19672
rect 39485 19669 39497 19703
rect 39531 19669 39543 19703
rect 39485 19663 39543 19669
rect 40589 19703 40647 19709
rect 40589 19669 40601 19703
rect 40635 19700 40647 19703
rect 41690 19700 41696 19712
rect 40635 19672 41696 19700
rect 40635 19669 40647 19672
rect 40589 19663 40647 19669
rect 41690 19660 41696 19672
rect 41748 19660 41754 19712
rect 1104 19610 43884 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 43884 19610
rect 1104 19536 43884 19558
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 15102 19496 15108 19508
rect 14875 19468 15108 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 15102 19456 15108 19468
rect 15160 19496 15166 19508
rect 16301 19499 16359 19505
rect 16301 19496 16313 19499
rect 15160 19468 16313 19496
rect 15160 19456 15166 19468
rect 16301 19465 16313 19468
rect 16347 19496 16359 19499
rect 16945 19499 17003 19505
rect 16945 19496 16957 19499
rect 16347 19468 16957 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 16945 19465 16957 19468
rect 16991 19465 17003 19499
rect 16945 19459 17003 19465
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 20254 19496 20260 19508
rect 19484 19468 20260 19496
rect 19484 19456 19490 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 22922 19456 22928 19508
rect 22980 19456 22986 19508
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 23842 19496 23848 19508
rect 23072 19468 23848 19496
rect 23072 19456 23078 19468
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 23934 19456 23940 19508
rect 23992 19456 23998 19508
rect 25498 19496 25504 19508
rect 24044 19468 25504 19496
rect 15746 19428 15752 19440
rect 14660 19400 15752 19428
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 14660 19369 14688 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 17218 19428 17224 19440
rect 15948 19400 17224 19428
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 12032 19332 12173 19360
rect 12032 19320 12038 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 14918 19320 14924 19372
rect 14976 19320 14982 19372
rect 15948 19369 15976 19400
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 24044 19428 24072 19468
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 28718 19456 28724 19508
rect 28776 19456 28782 19508
rect 28902 19456 28908 19508
rect 28960 19496 28966 19508
rect 29914 19496 29920 19508
rect 28960 19468 29920 19496
rect 28960 19456 28966 19468
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 31754 19456 31760 19508
rect 31812 19456 31818 19508
rect 32309 19499 32367 19505
rect 32309 19465 32321 19499
rect 32355 19465 32367 19499
rect 34149 19499 34207 19505
rect 34149 19496 34161 19499
rect 32309 19459 32367 19465
rect 33612 19468 34161 19496
rect 25593 19431 25651 19437
rect 25593 19428 25605 19431
rect 23860 19400 24072 19428
rect 24872 19400 25605 19428
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 17000 19332 17325 19360
rect 17000 19320 17006 19332
rect 17313 19329 17325 19332
rect 17359 19360 17371 19363
rect 17359 19332 17908 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 14274 19292 14280 19304
rect 12483 19264 14280 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 17221 19295 17279 19301
rect 17221 19261 17233 19295
rect 17267 19292 17279 19295
rect 17267 19264 17816 19292
rect 17267 19261 17279 19264
rect 17221 19255 17279 19261
rect 13722 19184 13728 19236
rect 13780 19184 13786 19236
rect 14461 19159 14519 19165
rect 14461 19125 14473 19159
rect 14507 19156 14519 19159
rect 14550 19156 14556 19168
rect 14507 19128 14556 19156
rect 14507 19125 14519 19128
rect 14461 19119 14519 19125
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 15657 19159 15715 19165
rect 15657 19156 15669 19159
rect 15344 19128 15669 19156
rect 15344 19116 15350 19128
rect 15657 19125 15669 19128
rect 15703 19125 15715 19159
rect 15657 19119 15715 19125
rect 17218 19116 17224 19168
rect 17276 19116 17282 19168
rect 17788 19156 17816 19264
rect 17880 19233 17908 19332
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18598 19360 18604 19372
rect 18371 19332 18604 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18598 19320 18604 19332
rect 18656 19360 18662 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 18656 19332 19441 19360
rect 18656 19320 18662 19332
rect 19429 19329 19441 19332
rect 19475 19360 19487 19363
rect 19475 19332 20668 19360
rect 19475 19329 19487 19332
rect 19429 19323 19487 19329
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 19242 19292 19248 19304
rect 18555 19264 19248 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 20640 19292 20668 19332
rect 23106 19320 23112 19372
rect 23164 19320 23170 19372
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 23860 19369 23888 19400
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 24762 19320 24768 19372
rect 24820 19320 24826 19372
rect 24872 19369 24900 19400
rect 25593 19397 25605 19400
rect 25639 19397 25651 19431
rect 25593 19391 25651 19397
rect 25682 19388 25688 19440
rect 25740 19428 25746 19440
rect 25961 19431 26019 19437
rect 25961 19428 25973 19431
rect 25740 19400 25973 19428
rect 25740 19388 25746 19400
rect 25961 19397 25973 19400
rect 26007 19397 26019 19431
rect 25961 19391 26019 19397
rect 28261 19431 28319 19437
rect 28261 19397 28273 19431
rect 28307 19428 28319 19431
rect 29086 19428 29092 19440
rect 28307 19400 29092 19428
rect 28307 19397 28319 19400
rect 28261 19391 28319 19397
rect 29086 19388 29092 19400
rect 29144 19388 29150 19440
rect 32122 19428 32128 19440
rect 30392 19400 32128 19428
rect 24857 19363 24915 19369
rect 24857 19329 24869 19363
rect 24903 19329 24915 19363
rect 24857 19323 24915 19329
rect 25038 19320 25044 19372
rect 25096 19360 25102 19372
rect 25133 19363 25191 19369
rect 25133 19360 25145 19363
rect 25096 19332 25145 19360
rect 25096 19320 25102 19332
rect 25133 19329 25145 19332
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 25314 19320 25320 19372
rect 25372 19360 25378 19372
rect 25777 19363 25835 19369
rect 25777 19360 25789 19363
rect 25372 19332 25789 19360
rect 25372 19320 25378 19332
rect 25777 19329 25789 19332
rect 25823 19329 25835 19363
rect 25777 19323 25835 19329
rect 26050 19320 26056 19372
rect 26108 19320 26114 19372
rect 27798 19320 27804 19372
rect 27856 19360 27862 19372
rect 28077 19363 28135 19369
rect 28077 19360 28089 19363
rect 27856 19332 28089 19360
rect 27856 19320 27862 19332
rect 28077 19329 28089 19332
rect 28123 19360 28135 19363
rect 28350 19360 28356 19372
rect 28123 19332 28356 19360
rect 28123 19329 28135 19332
rect 28077 19323 28135 19329
rect 28350 19320 28356 19332
rect 28408 19320 28414 19372
rect 28442 19320 28448 19372
rect 28500 19360 28506 19372
rect 28902 19360 28908 19372
rect 28500 19332 28908 19360
rect 28500 19320 28506 19332
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29181 19363 29239 19369
rect 29181 19360 29193 19363
rect 29012 19332 29193 19360
rect 29012 19304 29040 19332
rect 29181 19329 29193 19332
rect 29227 19329 29239 19363
rect 29181 19323 29239 19329
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 30392 19369 30420 19400
rect 32122 19388 32128 19400
rect 32180 19388 32186 19440
rect 30377 19363 30435 19369
rect 29696 19332 30328 19360
rect 29696 19320 29702 19332
rect 21266 19292 21272 19304
rect 20640 19264 21272 19292
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 23385 19295 23443 19301
rect 23385 19261 23397 19295
rect 23431 19292 23443 19295
rect 27893 19295 27951 19301
rect 23431 19264 24900 19292
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 24872 19236 24900 19264
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 28994 19292 29000 19304
rect 27939 19264 29000 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 28994 19252 29000 19264
rect 29052 19252 29058 19304
rect 29086 19252 29092 19304
rect 29144 19292 29150 19304
rect 30098 19292 30104 19304
rect 29144 19264 30104 19292
rect 29144 19252 29150 19264
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30300 19301 30328 19332
rect 30377 19329 30389 19363
rect 30423 19329 30435 19363
rect 31389 19363 31447 19369
rect 31389 19360 31401 19363
rect 30377 19323 30435 19329
rect 30484 19332 31401 19360
rect 30285 19295 30343 19301
rect 30285 19261 30297 19295
rect 30331 19261 30343 19295
rect 30285 19255 30343 19261
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19193 17923 19227
rect 24581 19227 24639 19233
rect 24581 19224 24593 19227
rect 17865 19187 17923 19193
rect 23768 19196 24593 19224
rect 18414 19156 18420 19168
rect 17788 19128 18420 19156
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19156 19579 19159
rect 19702 19156 19708 19168
rect 19567 19128 19708 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 23768 19156 23796 19196
rect 24581 19193 24593 19196
rect 24627 19193 24639 19227
rect 24581 19187 24639 19193
rect 24854 19184 24860 19236
rect 24912 19224 24918 19236
rect 25041 19227 25099 19233
rect 25041 19224 25053 19227
rect 24912 19196 25053 19224
rect 24912 19184 24918 19196
rect 25041 19193 25053 19196
rect 25087 19224 25099 19227
rect 25866 19224 25872 19236
rect 25087 19196 25872 19224
rect 25087 19193 25099 19196
rect 25041 19187 25099 19193
rect 25866 19184 25872 19196
rect 25924 19184 25930 19236
rect 29365 19227 29423 19233
rect 29365 19193 29377 19227
rect 29411 19224 29423 19227
rect 30484 19224 30512 19332
rect 31389 19329 31401 19332
rect 31435 19329 31447 19363
rect 32324 19360 32352 19459
rect 33444 19431 33502 19437
rect 33444 19397 33456 19431
rect 33490 19428 33502 19431
rect 33612 19428 33640 19468
rect 34149 19465 34161 19468
rect 34195 19465 34207 19499
rect 34149 19459 34207 19465
rect 34422 19456 34428 19508
rect 34480 19496 34486 19508
rect 38838 19496 38844 19508
rect 34480 19468 38844 19496
rect 34480 19456 34486 19468
rect 38838 19456 38844 19468
rect 38896 19496 38902 19508
rect 39666 19496 39672 19508
rect 38896 19468 39672 19496
rect 38896 19456 38902 19468
rect 39666 19456 39672 19468
rect 39724 19456 39730 19508
rect 39758 19456 39764 19508
rect 39816 19456 39822 19508
rect 41598 19456 41604 19508
rect 41656 19456 41662 19508
rect 41690 19456 41696 19508
rect 41748 19496 41754 19508
rect 42886 19496 42892 19508
rect 41748 19468 42892 19496
rect 41748 19456 41754 19468
rect 42886 19456 42892 19468
rect 42944 19456 42950 19508
rect 42978 19456 42984 19508
rect 43036 19456 43042 19508
rect 35710 19428 35716 19440
rect 33490 19400 33640 19428
rect 33704 19400 35716 19428
rect 33490 19397 33502 19400
rect 33444 19391 33502 19397
rect 33704 19369 33732 19400
rect 35710 19388 35716 19400
rect 35768 19388 35774 19440
rect 39298 19388 39304 19440
rect 39356 19428 39362 19440
rect 39393 19431 39451 19437
rect 39393 19428 39405 19431
rect 39356 19400 39405 19428
rect 39356 19388 39362 19400
rect 39393 19397 39405 19400
rect 39439 19397 39451 19431
rect 39393 19391 39451 19397
rect 42702 19388 42708 19440
rect 42760 19428 42766 19440
rect 43073 19431 43131 19437
rect 43073 19428 43085 19431
rect 42760 19400 43085 19428
rect 42760 19388 42766 19400
rect 43073 19397 43085 19400
rect 43119 19397 43131 19431
rect 43073 19391 43131 19397
rect 33689 19363 33747 19369
rect 32324 19332 33640 19360
rect 31389 19323 31447 19329
rect 31297 19295 31355 19301
rect 31297 19292 31309 19295
rect 30760 19264 31309 19292
rect 30760 19233 30788 19264
rect 31297 19261 31309 19264
rect 31343 19261 31355 19295
rect 33612 19292 33640 19332
rect 33689 19329 33701 19363
rect 33735 19329 33747 19363
rect 34238 19360 34244 19372
rect 33689 19323 33747 19329
rect 33796 19332 34244 19360
rect 33796 19292 33824 19332
rect 34238 19320 34244 19332
rect 34296 19360 34302 19372
rect 34517 19363 34575 19369
rect 34517 19360 34529 19363
rect 34296 19332 34529 19360
rect 34296 19320 34302 19332
rect 34517 19329 34529 19332
rect 34563 19329 34575 19363
rect 34517 19323 34575 19329
rect 37366 19320 37372 19372
rect 37424 19360 37430 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37424 19332 37473 19360
rect 37424 19320 37430 19332
rect 37461 19329 37473 19332
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 37642 19320 37648 19372
rect 37700 19360 37706 19372
rect 37737 19363 37795 19369
rect 37737 19360 37749 19363
rect 37700 19332 37749 19360
rect 37700 19320 37706 19332
rect 37737 19329 37749 19332
rect 37783 19329 37795 19363
rect 37737 19323 37795 19329
rect 37826 19320 37832 19372
rect 37884 19320 37890 19372
rect 39574 19320 39580 19372
rect 39632 19320 39638 19372
rect 33612 19264 33824 19292
rect 34609 19295 34667 19301
rect 31297 19255 31355 19261
rect 34609 19261 34621 19295
rect 34655 19292 34667 19295
rect 34698 19292 34704 19304
rect 34655 19264 34704 19292
rect 34655 19261 34667 19264
rect 34609 19255 34667 19261
rect 34698 19252 34704 19264
rect 34756 19252 34762 19304
rect 34793 19295 34851 19301
rect 34793 19261 34805 19295
rect 34839 19292 34851 19295
rect 41785 19295 41843 19301
rect 41785 19292 41797 19295
rect 34839 19264 41797 19292
rect 34839 19261 34851 19264
rect 34793 19255 34851 19261
rect 41785 19261 41797 19264
rect 41831 19292 41843 19295
rect 43165 19295 43223 19301
rect 43165 19292 43177 19295
rect 41831 19264 43177 19292
rect 41831 19261 41843 19264
rect 41785 19255 41843 19261
rect 43165 19261 43177 19264
rect 43211 19292 43223 19295
rect 43254 19292 43260 19304
rect 43211 19264 43260 19292
rect 43211 19261 43223 19264
rect 43165 19255 43223 19261
rect 43254 19252 43260 19264
rect 43312 19252 43318 19304
rect 29411 19196 30512 19224
rect 30745 19227 30803 19233
rect 29411 19193 29423 19196
rect 29365 19187 29423 19193
rect 30745 19193 30757 19227
rect 30791 19193 30803 19227
rect 30745 19187 30803 19193
rect 38013 19227 38071 19233
rect 38013 19193 38025 19227
rect 38059 19224 38071 19227
rect 42702 19224 42708 19236
rect 38059 19196 42708 19224
rect 38059 19193 38071 19196
rect 38013 19187 38071 19193
rect 42702 19184 42708 19196
rect 42760 19184 42766 19236
rect 20956 19128 23796 19156
rect 37553 19159 37611 19165
rect 20956 19116 20962 19128
rect 37553 19125 37565 19159
rect 37599 19156 37611 19159
rect 40126 19156 40132 19168
rect 37599 19128 40132 19156
rect 37599 19125 37611 19128
rect 37553 19119 37611 19125
rect 40126 19116 40132 19128
rect 40184 19116 40190 19168
rect 41230 19116 41236 19168
rect 41288 19116 41294 19168
rect 42610 19116 42616 19168
rect 42668 19116 42674 19168
rect 1104 19066 43884 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 43884 19066
rect 1104 18992 43884 19014
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 16485 18955 16543 18961
rect 16485 18952 16497 18955
rect 15896 18924 16497 18952
rect 15896 18912 15902 18924
rect 16485 18921 16497 18924
rect 16531 18921 16543 18955
rect 16485 18915 16543 18921
rect 22066 18924 23520 18952
rect 22066 18884 22094 18924
rect 23382 18884 23388 18896
rect 18616 18856 22094 18884
rect 23216 18856 23388 18884
rect 18616 18825 18644 18856
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 20622 18816 20628 18828
rect 18601 18779 18659 18785
rect 20364 18788 20628 18816
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 14476 18612 14504 18711
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 15102 18708 15108 18760
rect 15160 18708 15166 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 15746 18748 15752 18760
rect 15427 18720 15752 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 16942 18748 16948 18760
rect 16899 18720 16948 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 18138 18748 18144 18760
rect 17543 18720 18144 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19392 18720 19533 18748
rect 19392 18708 19398 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 19978 18748 19984 18760
rect 19760 18720 19984 18748
rect 19760 18708 19766 18720
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20364 18757 20392 18788
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 21453 18819 21511 18825
rect 21453 18816 21465 18819
rect 21324 18788 21465 18816
rect 21324 18776 21330 18788
rect 21453 18785 21465 18788
rect 21499 18785 21511 18819
rect 21453 18779 21511 18785
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 23216 18816 23244 18856
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 23492 18884 23520 18924
rect 25222 18912 25228 18964
rect 25280 18912 25286 18964
rect 25593 18955 25651 18961
rect 25593 18921 25605 18955
rect 25639 18952 25651 18955
rect 26050 18952 26056 18964
rect 25639 18924 26056 18952
rect 25639 18921 25651 18924
rect 25593 18915 25651 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 28166 18912 28172 18964
rect 28224 18952 28230 18964
rect 28445 18955 28503 18961
rect 28445 18952 28457 18955
rect 28224 18924 28457 18952
rect 28224 18912 28230 18924
rect 28445 18921 28457 18924
rect 28491 18921 28503 18955
rect 28445 18915 28503 18921
rect 33778 18912 33784 18964
rect 33836 18952 33842 18964
rect 35345 18955 35403 18961
rect 35345 18952 35357 18955
rect 33836 18924 35357 18952
rect 33836 18912 33842 18924
rect 35345 18921 35357 18924
rect 35391 18952 35403 18955
rect 35434 18952 35440 18964
rect 35391 18924 35440 18952
rect 35391 18921 35403 18924
rect 35345 18915 35403 18921
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 42978 18912 42984 18964
rect 43036 18952 43042 18964
rect 43165 18955 43223 18961
rect 43165 18952 43177 18955
rect 43036 18924 43177 18952
rect 43036 18912 43042 18924
rect 43165 18921 43177 18924
rect 43211 18921 43223 18955
rect 43165 18915 43223 18921
rect 25406 18884 25412 18896
rect 23492 18856 25412 18884
rect 25406 18844 25412 18856
rect 25464 18844 25470 18896
rect 28718 18884 28724 18896
rect 28644 18856 28724 18884
rect 28644 18825 28672 18856
rect 28718 18844 28724 18856
rect 28776 18844 28782 18896
rect 34698 18844 34704 18896
rect 34756 18884 34762 18896
rect 34756 18856 39712 18884
rect 34756 18844 34762 18856
rect 21683 18788 23244 18816
rect 23293 18819 23351 18825
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 23293 18785 23305 18819
rect 23339 18785 23351 18819
rect 23293 18779 23351 18785
rect 28629 18819 28687 18825
rect 28629 18785 28641 18819
rect 28675 18785 28687 18819
rect 28994 18816 29000 18828
rect 28629 18779 28687 18785
rect 28736 18788 29000 18816
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18748 20591 18751
rect 22646 18748 22652 18760
rect 20579 18720 22652 18748
rect 20579 18717 20591 18720
rect 20533 18711 20591 18717
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 23308 18748 23336 18779
rect 22888 18720 23336 18748
rect 22888 18708 22894 18720
rect 23750 18708 23756 18760
rect 23808 18748 23814 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 23808 18720 25421 18748
rect 23808 18708 23814 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 25682 18708 25688 18760
rect 25740 18708 25746 18760
rect 28736 18757 28764 18788
rect 28994 18776 29000 18788
rect 29052 18776 29058 18828
rect 35342 18776 35348 18828
rect 35400 18776 35406 18828
rect 28721 18751 28779 18757
rect 28721 18717 28733 18751
rect 28767 18717 28779 18751
rect 28721 18711 28779 18717
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 14918 18640 14924 18692
rect 14976 18680 14982 18692
rect 15197 18683 15255 18689
rect 15197 18680 15209 18683
rect 14976 18652 15209 18680
rect 14976 18640 14982 18652
rect 15197 18649 15209 18652
rect 15243 18649 15255 18683
rect 15197 18643 15255 18649
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 17328 18680 17356 18708
rect 16724 18652 17356 18680
rect 17405 18683 17463 18689
rect 16724 18640 16730 18652
rect 17405 18649 17417 18683
rect 17451 18680 17463 18683
rect 18230 18680 18236 18692
rect 17451 18652 18236 18680
rect 17451 18649 17463 18652
rect 17405 18643 17463 18649
rect 18230 18640 18236 18652
rect 18288 18680 18294 18692
rect 18325 18683 18383 18689
rect 18325 18680 18337 18683
rect 18288 18652 18337 18680
rect 18288 18640 18294 18652
rect 18325 18649 18337 18652
rect 18371 18649 18383 18683
rect 18432 18680 18460 18708
rect 19429 18683 19487 18689
rect 19429 18680 19441 18683
rect 18432 18652 19441 18680
rect 18325 18643 18383 18649
rect 19429 18649 19441 18652
rect 19475 18649 19487 18683
rect 23109 18683 23167 18689
rect 23109 18680 23121 18683
rect 19429 18643 19487 18649
rect 21376 18652 23121 18680
rect 21376 18624 21404 18652
rect 23109 18649 23121 18652
rect 23155 18649 23167 18683
rect 28828 18680 28856 18711
rect 28902 18708 28908 18760
rect 28960 18708 28966 18760
rect 33686 18708 33692 18760
rect 33744 18748 33750 18760
rect 34790 18748 34796 18760
rect 33744 18720 34796 18748
rect 33744 18708 33750 18720
rect 34790 18708 34796 18720
rect 34848 18748 34854 18760
rect 34977 18751 35035 18757
rect 34977 18748 34989 18751
rect 34848 18720 34989 18748
rect 34848 18708 34854 18720
rect 34977 18717 34989 18720
rect 35023 18717 35035 18751
rect 34977 18711 35035 18717
rect 36262 18708 36268 18760
rect 36320 18708 36326 18760
rect 36446 18708 36452 18760
rect 36504 18708 36510 18760
rect 29086 18680 29092 18692
rect 28828 18652 29092 18680
rect 23109 18643 23167 18649
rect 29086 18640 29092 18652
rect 29144 18640 29150 18692
rect 39574 18680 39580 18692
rect 35176 18652 39580 18680
rect 14826 18612 14832 18624
rect 14476 18584 14832 18612
rect 14826 18572 14832 18584
rect 14884 18612 14890 18624
rect 15105 18615 15163 18621
rect 15105 18612 15117 18615
rect 14884 18584 15117 18612
rect 14884 18572 14890 18584
rect 15105 18581 15117 18584
rect 15151 18581 15163 18615
rect 15105 18575 15163 18581
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 18417 18615 18475 18621
rect 18417 18612 18429 18615
rect 18196 18584 18429 18612
rect 18196 18572 18202 18584
rect 18417 18581 18429 18584
rect 18463 18612 18475 18615
rect 18598 18612 18604 18624
rect 18463 18584 18604 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 20990 18572 20996 18624
rect 21048 18572 21054 18624
rect 21358 18572 21364 18624
rect 21416 18572 21422 18624
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 35176 18621 35204 18652
rect 39574 18640 39580 18652
rect 39632 18640 39638 18692
rect 39684 18680 39712 18856
rect 40678 18708 40684 18760
rect 40736 18748 40742 18760
rect 41506 18748 41512 18760
rect 40736 18720 41512 18748
rect 40736 18708 40742 18720
rect 41506 18708 41512 18720
rect 41564 18748 41570 18760
rect 41785 18751 41843 18757
rect 41785 18748 41797 18751
rect 41564 18720 41797 18748
rect 41564 18708 41570 18720
rect 41785 18717 41797 18720
rect 41831 18717 41843 18751
rect 41785 18711 41843 18717
rect 42052 18751 42110 18757
rect 42052 18717 42064 18751
rect 42098 18748 42110 18751
rect 42610 18748 42616 18760
rect 42098 18720 42616 18748
rect 42098 18717 42110 18720
rect 42052 18711 42110 18717
rect 42610 18708 42616 18720
rect 42668 18708 42674 18760
rect 42794 18680 42800 18692
rect 39684 18652 42800 18680
rect 42794 18640 42800 18652
rect 42852 18640 42858 18692
rect 23201 18615 23259 18621
rect 23201 18612 23213 18615
rect 22980 18584 23213 18612
rect 22980 18572 22986 18584
rect 23201 18581 23213 18584
rect 23247 18581 23259 18615
rect 23201 18575 23259 18581
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18581 35219 18615
rect 35161 18575 35219 18581
rect 36357 18615 36415 18621
rect 36357 18581 36369 18615
rect 36403 18612 36415 18615
rect 37550 18612 37556 18624
rect 36403 18584 37556 18612
rect 36403 18581 36415 18584
rect 36357 18575 36415 18581
rect 37550 18572 37556 18584
rect 37608 18572 37614 18624
rect 1104 18522 43884 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 43884 18522
rect 1104 18448 43884 18470
rect 15381 18411 15439 18417
rect 15381 18377 15393 18411
rect 15427 18408 15439 18411
rect 15470 18408 15476 18420
rect 15427 18380 15476 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 18690 18368 18696 18420
rect 18748 18368 18754 18420
rect 19889 18411 19947 18417
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 19978 18408 19984 18420
rect 19935 18380 19984 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 21266 18368 21272 18420
rect 21324 18408 21330 18420
rect 22922 18408 22928 18420
rect 21324 18380 22928 18408
rect 21324 18368 21330 18380
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 28629 18411 28687 18417
rect 28629 18377 28641 18411
rect 28675 18408 28687 18411
rect 28994 18408 29000 18420
rect 28675 18380 29000 18408
rect 28675 18377 28687 18380
rect 28629 18371 28687 18377
rect 28994 18368 29000 18380
rect 29052 18368 29058 18420
rect 38838 18368 38844 18420
rect 38896 18368 38902 18420
rect 41598 18368 41604 18420
rect 41656 18408 41662 18420
rect 42061 18411 42119 18417
rect 42061 18408 42073 18411
rect 41656 18380 42073 18408
rect 41656 18368 41662 18380
rect 42061 18377 42073 18380
rect 42107 18377 42119 18411
rect 42061 18371 42119 18377
rect 17313 18343 17371 18349
rect 17313 18309 17325 18343
rect 17359 18340 17371 18343
rect 17954 18340 17960 18352
rect 17359 18312 17960 18340
rect 17359 18309 17371 18312
rect 17313 18303 17371 18309
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 18230 18300 18236 18352
rect 18288 18340 18294 18352
rect 18708 18340 18736 18368
rect 21358 18340 21364 18352
rect 18288 18312 18644 18340
rect 18708 18312 21364 18340
rect 18288 18300 18294 18312
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14976 18244 15025 18272
rect 14976 18232 14982 18244
rect 15013 18241 15025 18244
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18414 18272 18420 18284
rect 17543 18244 18420 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18616 18281 18644 18312
rect 20824 18281 20852 18312
rect 21358 18300 21364 18312
rect 21416 18340 21422 18352
rect 22741 18343 22799 18349
rect 22741 18340 22753 18343
rect 21416 18312 22753 18340
rect 21416 18300 21422 18312
rect 22741 18309 22753 18312
rect 22787 18309 22799 18343
rect 22741 18303 22799 18309
rect 23014 18300 23020 18352
rect 23072 18300 23078 18352
rect 28445 18343 28503 18349
rect 28445 18309 28457 18343
rect 28491 18340 28503 18343
rect 29086 18340 29092 18352
rect 28491 18312 29092 18340
rect 28491 18309 28503 18312
rect 28445 18303 28503 18309
rect 29086 18300 29092 18312
rect 29144 18300 29150 18352
rect 30190 18300 30196 18352
rect 30248 18340 30254 18352
rect 30650 18340 30656 18352
rect 30248 18312 30656 18340
rect 30248 18300 30254 18312
rect 30650 18300 30656 18312
rect 30708 18340 30714 18352
rect 34793 18343 34851 18349
rect 34793 18340 34805 18343
rect 30708 18312 34805 18340
rect 30708 18300 30714 18312
rect 34793 18309 34805 18312
rect 34839 18340 34851 18343
rect 35802 18340 35808 18352
rect 34839 18312 35808 18340
rect 34839 18309 34851 18312
rect 34793 18303 34851 18309
rect 35802 18300 35808 18312
rect 35860 18300 35866 18352
rect 40948 18343 41006 18349
rect 35912 18312 40080 18340
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18272 19855 18275
rect 20717 18275 20775 18281
rect 20717 18272 20729 18275
rect 19843 18244 20729 18272
rect 19843 18241 19855 18244
rect 19797 18235 19855 18241
rect 20717 18241 20729 18244
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 22646 18232 22652 18284
rect 22704 18272 22710 18284
rect 25682 18272 25688 18284
rect 22704 18244 25688 18272
rect 22704 18232 22710 18244
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 28718 18232 28724 18284
rect 28776 18232 28782 18284
rect 33778 18232 33784 18284
rect 33836 18272 33842 18284
rect 33873 18275 33931 18281
rect 33873 18272 33885 18275
rect 33836 18244 33885 18272
rect 33836 18232 33842 18244
rect 33873 18241 33885 18244
rect 33919 18241 33931 18275
rect 33873 18235 33931 18241
rect 35621 18275 35679 18281
rect 35621 18241 35633 18275
rect 35667 18272 35679 18275
rect 35710 18272 35716 18284
rect 35667 18244 35716 18272
rect 35667 18241 35679 18244
rect 35621 18235 35679 18241
rect 35710 18232 35716 18244
rect 35768 18272 35774 18284
rect 35912 18272 35940 18312
rect 35768 18244 35940 18272
rect 36357 18275 36415 18281
rect 35768 18232 35774 18244
rect 36357 18241 36369 18275
rect 36403 18272 36415 18275
rect 36446 18272 36452 18284
rect 36403 18244 36452 18272
rect 36403 18241 36415 18244
rect 36357 18235 36415 18241
rect 20073 18207 20131 18213
rect 20073 18173 20085 18207
rect 20119 18204 20131 18207
rect 20346 18204 20352 18216
rect 20119 18176 20352 18204
rect 20119 18173 20131 18176
rect 20073 18167 20131 18173
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 29362 18164 29368 18216
rect 29420 18164 29426 18216
rect 35342 18164 35348 18216
rect 35400 18204 35406 18216
rect 36265 18207 36323 18213
rect 36265 18204 36277 18207
rect 35400 18176 36277 18204
rect 35400 18164 35406 18176
rect 36265 18173 36277 18176
rect 36311 18173 36323 18207
rect 36265 18167 36323 18173
rect 16942 18096 16948 18148
rect 17000 18136 17006 18148
rect 17129 18139 17187 18145
rect 17129 18136 17141 18139
rect 17000 18108 17141 18136
rect 17000 18096 17006 18108
rect 17129 18105 17141 18108
rect 17175 18105 17187 18139
rect 17129 18099 17187 18105
rect 22278 18096 22284 18148
rect 22336 18136 22342 18148
rect 23106 18136 23112 18148
rect 22336 18108 23112 18136
rect 22336 18096 22342 18108
rect 23106 18096 23112 18108
rect 23164 18096 23170 18148
rect 28074 18096 28080 18148
rect 28132 18136 28138 18148
rect 28445 18139 28503 18145
rect 28445 18136 28457 18139
rect 28132 18108 28457 18136
rect 28132 18096 28138 18108
rect 28445 18105 28457 18108
rect 28491 18105 28503 18139
rect 28445 18099 28503 18105
rect 33686 18096 33692 18148
rect 33744 18136 33750 18148
rect 34149 18139 34207 18145
rect 34149 18136 34161 18139
rect 33744 18108 34161 18136
rect 33744 18096 33750 18108
rect 34149 18105 34161 18108
rect 34195 18105 34207 18139
rect 34149 18099 34207 18105
rect 34333 18139 34391 18145
rect 34333 18105 34345 18139
rect 34379 18136 34391 18139
rect 36372 18136 36400 18235
rect 36446 18232 36452 18244
rect 36504 18232 36510 18284
rect 37476 18281 37504 18312
rect 40052 18284 40080 18312
rect 40948 18309 40960 18343
rect 40994 18340 41006 18343
rect 41230 18340 41236 18352
rect 40994 18312 41236 18340
rect 40994 18309 41006 18312
rect 40948 18303 41006 18309
rect 41230 18300 41236 18312
rect 41288 18300 41294 18352
rect 43162 18300 43168 18352
rect 43220 18300 43226 18352
rect 37461 18275 37519 18281
rect 37461 18241 37473 18275
rect 37507 18241 37519 18275
rect 37461 18235 37519 18241
rect 37550 18232 37556 18284
rect 37608 18272 37614 18284
rect 37717 18275 37775 18281
rect 37717 18272 37729 18275
rect 37608 18244 37729 18272
rect 37608 18232 37614 18244
rect 37717 18241 37729 18244
rect 37763 18241 37775 18275
rect 37717 18235 37775 18241
rect 39574 18232 39580 18284
rect 39632 18232 39638 18284
rect 40034 18232 40040 18284
rect 40092 18272 40098 18284
rect 40678 18272 40684 18284
rect 40092 18244 40684 18272
rect 40092 18232 40098 18244
rect 40678 18232 40684 18244
rect 40736 18232 40742 18284
rect 42886 18232 42892 18284
rect 42944 18232 42950 18284
rect 39298 18164 39304 18216
rect 39356 18204 39362 18216
rect 39485 18207 39543 18213
rect 39485 18204 39497 18207
rect 39356 18176 39497 18204
rect 39356 18164 39362 18176
rect 39485 18173 39497 18176
rect 39531 18173 39543 18207
rect 39485 18167 39543 18173
rect 34379 18108 36400 18136
rect 34379 18105 34391 18108
rect 34333 18099 34391 18105
rect 19426 18028 19432 18080
rect 19484 18028 19490 18080
rect 22465 18071 22523 18077
rect 22465 18037 22477 18071
rect 22511 18068 22523 18071
rect 23382 18068 23388 18080
rect 22511 18040 23388 18068
rect 22511 18037 22523 18040
rect 22465 18031 22523 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 36538 18028 36544 18080
rect 36596 18068 36602 18080
rect 36633 18071 36691 18077
rect 36633 18068 36645 18071
rect 36596 18040 36645 18068
rect 36596 18028 36602 18040
rect 36633 18037 36645 18040
rect 36679 18037 36691 18071
rect 36633 18031 36691 18037
rect 39945 18071 40003 18077
rect 39945 18037 39957 18071
rect 39991 18068 40003 18071
rect 40310 18068 40316 18080
rect 39991 18040 40316 18068
rect 39991 18037 40003 18040
rect 39945 18031 40003 18037
rect 40310 18028 40316 18040
rect 40368 18028 40374 18080
rect 1104 17978 43884 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 43884 17978
rect 1104 17904 43884 17926
rect 14645 17867 14703 17873
rect 14645 17833 14657 17867
rect 14691 17864 14703 17867
rect 15194 17864 15200 17876
rect 14691 17836 15200 17864
rect 14691 17833 14703 17836
rect 14645 17827 14703 17833
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 22373 17867 22431 17873
rect 22373 17833 22385 17867
rect 22419 17864 22431 17867
rect 22738 17864 22744 17876
rect 22419 17836 22744 17864
rect 22419 17833 22431 17836
rect 22373 17827 22431 17833
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 37458 17824 37464 17876
rect 37516 17864 37522 17876
rect 37645 17867 37703 17873
rect 37645 17864 37657 17867
rect 37516 17836 37657 17864
rect 37516 17824 37522 17836
rect 37645 17833 37657 17836
rect 37691 17833 37703 17867
rect 37645 17827 37703 17833
rect 41414 17824 41420 17876
rect 41472 17824 41478 17876
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 15105 17799 15163 17805
rect 15105 17796 15117 17799
rect 14976 17768 15117 17796
rect 14976 17756 14982 17768
rect 15105 17765 15117 17768
rect 15151 17765 15163 17799
rect 17770 17796 17776 17808
rect 15105 17759 15163 17765
rect 16684 17768 17776 17796
rect 16684 17737 16712 17768
rect 17770 17756 17776 17768
rect 17828 17796 17834 17808
rect 24118 17796 24124 17808
rect 17828 17768 24124 17796
rect 17828 17756 17834 17768
rect 24118 17756 24124 17768
rect 24176 17756 24182 17808
rect 28258 17756 28264 17808
rect 28316 17796 28322 17808
rect 28353 17799 28411 17805
rect 28353 17796 28365 17799
rect 28316 17768 28365 17796
rect 28316 17756 28322 17768
rect 28353 17765 28365 17768
rect 28399 17765 28411 17799
rect 28353 17759 28411 17765
rect 33781 17799 33839 17805
rect 33781 17765 33793 17799
rect 33827 17796 33839 17799
rect 33870 17796 33876 17808
rect 33827 17768 33876 17796
rect 33827 17765 33839 17768
rect 33781 17759 33839 17765
rect 33870 17756 33876 17768
rect 33928 17756 33934 17808
rect 16669 17731 16727 17737
rect 14568 17700 15608 17728
rect 14568 17669 14596 17700
rect 15580 17672 15608 17700
rect 16669 17697 16681 17731
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19334 17728 19340 17740
rect 18831 17700 19340 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19334 17688 19340 17700
rect 19392 17728 19398 17740
rect 19392 17700 19840 17728
rect 19392 17688 19398 17700
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17561 14427 17595
rect 14660 17592 14688 17623
rect 15286 17620 15292 17672
rect 15344 17620 15350 17672
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 17368 17632 18705 17660
rect 17368 17620 17374 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 14660 17564 15485 17592
rect 14369 17555 14427 17561
rect 15473 17561 15485 17564
rect 15519 17592 15531 17595
rect 16022 17592 16028 17604
rect 15519 17564 16028 17592
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 14384 17524 14412 17555
rect 16022 17552 16028 17564
rect 16080 17592 16086 17604
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 16080 17564 16773 17592
rect 16080 17552 16086 17564
rect 16761 17561 16773 17564
rect 16807 17592 16819 17595
rect 17126 17592 17132 17604
rect 16807 17564 17132 17592
rect 16807 17561 16819 17564
rect 16761 17555 16819 17561
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 18708 17592 18736 17623
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19812 17669 19840 17700
rect 22094 17688 22100 17740
rect 22152 17728 22158 17740
rect 22465 17731 22523 17737
rect 22465 17728 22477 17731
rect 22152 17700 22477 17728
rect 22152 17688 22158 17700
rect 22465 17697 22477 17700
rect 22511 17728 22523 17731
rect 22646 17728 22652 17740
rect 22511 17700 22652 17728
rect 22511 17697 22523 17700
rect 22465 17691 22523 17697
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 29362 17728 29368 17740
rect 27540 17700 29368 17728
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19484 17632 19717 17660
rect 19484 17620 19490 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 19978 17620 19984 17672
rect 20036 17620 20042 17672
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20438 17660 20444 17672
rect 20119 17632 20444 17660
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22094 17592 22100 17604
rect 18708 17564 22100 17592
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22204 17592 22232 17623
rect 22738 17620 22744 17672
rect 22796 17660 22802 17672
rect 23017 17663 23075 17669
rect 23017 17660 23029 17663
rect 22796 17632 23029 17660
rect 22796 17620 22802 17632
rect 23017 17629 23029 17632
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 23198 17620 23204 17672
rect 23256 17620 23262 17672
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 26513 17663 26571 17669
rect 26513 17660 26525 17663
rect 26384 17632 26525 17660
rect 26384 17620 26390 17632
rect 26513 17629 26525 17632
rect 26559 17660 26571 17663
rect 27540 17660 27568 17700
rect 29362 17688 29368 17700
rect 29420 17728 29426 17740
rect 29733 17731 29791 17737
rect 29733 17728 29745 17731
rect 29420 17700 29745 17728
rect 29420 17688 29426 17700
rect 29733 17697 29745 17700
rect 29779 17697 29791 17731
rect 29733 17691 29791 17697
rect 31754 17688 31760 17740
rect 31812 17688 31818 17740
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17728 33011 17731
rect 35710 17728 35716 17740
rect 32999 17700 35716 17728
rect 32999 17697 33011 17700
rect 32953 17691 33011 17697
rect 35710 17688 35716 17700
rect 35768 17728 35774 17740
rect 36265 17731 36323 17737
rect 36265 17728 36277 17731
rect 35768 17700 36277 17728
rect 35768 17688 35774 17700
rect 36265 17697 36277 17700
rect 36311 17697 36323 17731
rect 36265 17691 36323 17697
rect 28629 17663 28687 17669
rect 28629 17660 28641 17663
rect 26559 17632 27568 17660
rect 27632 17632 28641 17660
rect 26559 17629 26571 17632
rect 26513 17623 26571 17629
rect 23216 17592 23244 17620
rect 22204 17564 23244 17592
rect 26780 17595 26838 17601
rect 26780 17561 26792 17595
rect 26826 17592 26838 17595
rect 27154 17592 27160 17604
rect 26826 17564 27160 17592
rect 26826 17561 26838 17564
rect 26780 17555 26838 17561
rect 27154 17552 27160 17564
rect 27212 17552 27218 17604
rect 27246 17552 27252 17604
rect 27304 17592 27310 17604
rect 27632 17592 27660 17632
rect 28629 17629 28641 17632
rect 28675 17629 28687 17663
rect 31772 17660 31800 17688
rect 31772 17632 32812 17660
rect 28629 17623 28687 17629
rect 27304 17564 27660 17592
rect 27304 17552 27310 17564
rect 28350 17552 28356 17604
rect 28408 17552 28414 17604
rect 30006 17601 30012 17604
rect 30000 17555 30012 17601
rect 30006 17552 30012 17555
rect 30064 17552 30070 17604
rect 31754 17552 31760 17604
rect 31812 17592 31818 17604
rect 32686 17595 32744 17601
rect 32686 17592 32698 17595
rect 31812 17564 32698 17592
rect 31812 17552 31818 17564
rect 32686 17561 32698 17564
rect 32732 17561 32744 17595
rect 32784 17592 32812 17632
rect 33410 17620 33416 17672
rect 33468 17620 33474 17672
rect 33781 17663 33839 17669
rect 33781 17629 33793 17663
rect 33827 17660 33839 17663
rect 33965 17663 34023 17669
rect 33827 17632 33916 17660
rect 33827 17629 33839 17632
rect 33781 17623 33839 17629
rect 33888 17592 33916 17632
rect 33965 17629 33977 17663
rect 34011 17660 34023 17663
rect 34011 17632 35664 17660
rect 34011 17629 34023 17632
rect 33965 17623 34023 17629
rect 32784 17564 33916 17592
rect 32686 17555 32744 17561
rect 15286 17524 15292 17536
rect 14384 17496 15292 17524
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 18656 17496 19533 17524
rect 18656 17484 18662 17496
rect 19521 17493 19533 17496
rect 19567 17493 19579 17527
rect 19521 17487 19579 17493
rect 22002 17484 22008 17536
rect 22060 17484 22066 17536
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22244 17496 23029 17524
rect 22244 17484 22250 17496
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 23017 17487 23075 17493
rect 27522 17484 27528 17536
rect 27580 17524 27586 17536
rect 27893 17527 27951 17533
rect 27893 17524 27905 17527
rect 27580 17496 27905 17524
rect 27580 17484 27586 17496
rect 27893 17493 27905 17496
rect 27939 17524 27951 17527
rect 28537 17527 28595 17533
rect 28537 17524 28549 17527
rect 27939 17496 28549 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 28537 17493 28549 17496
rect 28583 17493 28595 17527
rect 28537 17487 28595 17493
rect 31110 17484 31116 17536
rect 31168 17484 31174 17536
rect 31573 17527 31631 17533
rect 31573 17493 31585 17527
rect 31619 17524 31631 17527
rect 31846 17524 31852 17536
rect 31619 17496 31852 17524
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 31846 17484 31852 17496
rect 31904 17484 31910 17536
rect 33888 17524 33916 17564
rect 35069 17595 35127 17601
rect 35069 17561 35081 17595
rect 35115 17592 35127 17595
rect 35526 17592 35532 17604
rect 35115 17564 35532 17592
rect 35115 17561 35127 17564
rect 35069 17555 35127 17561
rect 35526 17552 35532 17564
rect 35584 17552 35590 17604
rect 35636 17592 35664 17632
rect 35802 17620 35808 17672
rect 35860 17620 35866 17672
rect 36538 17669 36544 17672
rect 36532 17660 36544 17669
rect 36499 17632 36544 17660
rect 36532 17623 36544 17632
rect 36538 17620 36544 17623
rect 36596 17620 36602 17672
rect 40034 17620 40040 17672
rect 40092 17620 40098 17672
rect 40310 17669 40316 17672
rect 40293 17663 40316 17669
rect 40293 17629 40305 17663
rect 40293 17623 40316 17629
rect 40310 17620 40316 17623
rect 40368 17620 40374 17672
rect 42794 17620 42800 17672
rect 42852 17660 42858 17672
rect 42889 17663 42947 17669
rect 42889 17660 42901 17663
rect 42852 17632 42901 17660
rect 42852 17620 42858 17632
rect 42889 17629 42901 17632
rect 42935 17629 42947 17663
rect 42889 17623 42947 17629
rect 35986 17592 35992 17604
rect 35636 17564 35992 17592
rect 35986 17552 35992 17564
rect 36044 17552 36050 17604
rect 43162 17552 43168 17604
rect 43220 17552 43226 17604
rect 37550 17524 37556 17536
rect 33888 17496 37556 17524
rect 37550 17484 37556 17496
rect 37608 17484 37614 17536
rect 1104 17434 43884 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 43884 17434
rect 1104 17360 43884 17382
rect 15289 17323 15347 17329
rect 15289 17289 15301 17323
rect 15335 17320 15347 17323
rect 15378 17320 15384 17332
rect 15335 17292 15384 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 18248 17292 22232 17320
rect 18248 17252 18276 17292
rect 22204 17264 22232 17292
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 23290 17320 23296 17332
rect 22520 17292 23296 17320
rect 22520 17280 22526 17292
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 23566 17280 23572 17332
rect 23624 17320 23630 17332
rect 23624 17292 27108 17320
rect 23624 17280 23630 17292
rect 19978 17252 19984 17264
rect 16316 17224 18276 17252
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15151 17156 15761 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 15028 17048 15056 17147
rect 15948 17116 15976 17147
rect 16022 17144 16028 17196
rect 16080 17144 16086 17196
rect 16206 17144 16212 17196
rect 16264 17144 16270 17196
rect 16316 17193 16344 17224
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 18248 17193 18276 17224
rect 19536 17224 19984 17252
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17184 19395 17187
rect 19426 17184 19432 17196
rect 19383 17156 19432 17184
rect 19383 17153 19395 17156
rect 19337 17147 19395 17153
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 15948 17088 17417 17116
rect 17405 17085 17417 17088
rect 17451 17116 17463 17119
rect 17586 17116 17592 17128
rect 17451 17088 17592 17116
rect 17451 17085 17463 17088
rect 17405 17079 17463 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17880 17116 17908 17147
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19536 17193 19564 17224
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 20990 17212 20996 17264
rect 21048 17252 21054 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 21048 17224 21097 17252
rect 21048 17212 21054 17224
rect 21085 17221 21097 17224
rect 21131 17221 21143 17255
rect 21085 17215 21143 17221
rect 22002 17212 22008 17264
rect 22060 17212 22066 17264
rect 22186 17212 22192 17264
rect 22244 17212 22250 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 25593 17255 25651 17261
rect 22336 17224 23060 17252
rect 22336 17212 22342 17224
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17184 19671 17187
rect 20438 17184 20444 17196
rect 19659 17156 20444 17184
rect 19659 17153 19671 17156
rect 19613 17147 19671 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 22462 17144 22468 17196
rect 22520 17184 22526 17196
rect 23032 17193 23060 17224
rect 25593 17221 25605 17255
rect 25639 17252 25651 17255
rect 25774 17252 25780 17264
rect 25639 17224 25780 17252
rect 25639 17221 25651 17224
rect 25593 17215 25651 17221
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22520 17156 22845 17184
rect 22520 17144 22526 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23017 17187 23075 17193
rect 23017 17153 23029 17187
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23566 17144 23572 17196
rect 23624 17184 23630 17196
rect 24213 17187 24271 17193
rect 24213 17184 24225 17187
rect 23624 17156 24225 17184
rect 23624 17144 23630 17156
rect 24213 17153 24225 17156
rect 24259 17153 24271 17187
rect 27080 17184 27108 17292
rect 27154 17280 27160 17332
rect 27212 17280 27218 17332
rect 27522 17280 27528 17332
rect 27580 17280 27586 17332
rect 27706 17280 27712 17332
rect 27764 17320 27770 17332
rect 29914 17320 29920 17332
rect 27764 17292 29920 17320
rect 27764 17280 27770 17292
rect 29914 17280 29920 17292
rect 29972 17320 29978 17332
rect 31297 17323 31355 17329
rect 31297 17320 31309 17323
rect 29972 17292 31309 17320
rect 29972 17280 29978 17292
rect 31297 17289 31309 17292
rect 31343 17289 31355 17323
rect 31297 17283 31355 17289
rect 31754 17280 31760 17332
rect 31812 17280 31818 17332
rect 35713 17323 35771 17329
rect 35713 17289 35725 17323
rect 35759 17320 35771 17323
rect 36262 17320 36268 17332
rect 35759 17292 36268 17320
rect 35759 17289 35771 17292
rect 35713 17283 35771 17289
rect 36262 17280 36268 17292
rect 36320 17280 36326 17332
rect 27430 17212 27436 17264
rect 27488 17252 27494 17264
rect 27617 17255 27675 17261
rect 27617 17252 27629 17255
rect 27488 17224 27629 17252
rect 27488 17212 27494 17224
rect 27617 17221 27629 17224
rect 27663 17221 27675 17255
rect 27617 17215 27675 17221
rect 34790 17212 34796 17264
rect 34848 17252 34854 17264
rect 35253 17255 35311 17261
rect 35253 17252 35265 17255
rect 34848 17224 35265 17252
rect 34848 17212 34854 17224
rect 35253 17221 35265 17224
rect 35299 17221 35311 17255
rect 35253 17215 35311 17221
rect 30377 17187 30435 17193
rect 30377 17184 30389 17187
rect 27080 17156 30389 17184
rect 24213 17147 24271 17153
rect 30377 17153 30389 17156
rect 30423 17184 30435 17187
rect 31389 17187 31447 17193
rect 30423 17156 31340 17184
rect 30423 17153 30435 17156
rect 30377 17147 30435 17153
rect 17880 17088 19656 17116
rect 15562 17048 15568 17060
rect 15028 17020 15568 17048
rect 15562 17008 15568 17020
rect 15620 17048 15626 17060
rect 16853 17051 16911 17057
rect 16853 17048 16865 17051
rect 15620 17020 16865 17048
rect 15620 17008 15626 17020
rect 16853 17017 16865 17020
rect 16899 17017 16911 17051
rect 16853 17011 16911 17017
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 17880 16980 17908 17088
rect 16264 16952 17908 16980
rect 16264 16940 16270 16952
rect 18782 16940 18788 16992
rect 18840 16980 18846 16992
rect 19153 16983 19211 16989
rect 19153 16980 19165 16983
rect 18840 16952 19165 16980
rect 18840 16940 18846 16952
rect 19153 16949 19165 16952
rect 19199 16949 19211 16983
rect 19628 16980 19656 17088
rect 20530 17076 20536 17128
rect 20588 17076 20594 17128
rect 23934 17116 23940 17128
rect 22066 17088 23940 17116
rect 22066 17060 22094 17088
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17116 27859 17119
rect 31202 17116 31208 17128
rect 27847 17088 31208 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 31202 17076 31208 17088
rect 31260 17076 31266 17128
rect 31312 17116 31340 17156
rect 31389 17153 31401 17187
rect 31435 17184 31447 17187
rect 31846 17184 31852 17196
rect 31435 17156 31852 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 31846 17144 31852 17156
rect 31904 17184 31910 17196
rect 32398 17184 32404 17196
rect 31904 17156 32404 17184
rect 31904 17144 31910 17156
rect 32398 17144 32404 17156
rect 32456 17144 32462 17196
rect 33502 17144 33508 17196
rect 33560 17144 33566 17196
rect 33594 17144 33600 17196
rect 33652 17184 33658 17196
rect 34333 17187 34391 17193
rect 34333 17184 34345 17187
rect 33652 17156 34345 17184
rect 33652 17144 33658 17156
rect 34333 17153 34345 17156
rect 34379 17184 34391 17187
rect 37274 17184 37280 17196
rect 34379 17156 37280 17184
rect 34379 17153 34391 17156
rect 34333 17147 34391 17153
rect 37274 17144 37280 17156
rect 37332 17184 37338 17196
rect 38194 17184 38200 17196
rect 37332 17156 38200 17184
rect 37332 17144 37338 17156
rect 38194 17144 38200 17156
rect 38252 17144 38258 17196
rect 31570 17116 31576 17128
rect 31312 17088 31576 17116
rect 31570 17076 31576 17088
rect 31628 17076 31634 17128
rect 34793 17119 34851 17125
rect 34793 17085 34805 17119
rect 34839 17116 34851 17119
rect 35986 17116 35992 17128
rect 34839 17088 35992 17116
rect 34839 17085 34851 17088
rect 34793 17079 34851 17085
rect 35986 17076 35992 17088
rect 36044 17076 36050 17128
rect 22002 17008 22008 17060
rect 22060 17020 22094 17060
rect 22060 17008 22066 17020
rect 35434 17008 35440 17060
rect 35492 17048 35498 17060
rect 35529 17051 35587 17057
rect 35529 17048 35541 17051
rect 35492 17020 35541 17048
rect 35492 17008 35498 17020
rect 35529 17017 35541 17020
rect 35575 17017 35587 17051
rect 35529 17011 35587 17017
rect 22094 16980 22100 16992
rect 19628 16952 22100 16980
rect 19153 16943 19211 16949
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 22281 16983 22339 16989
rect 22281 16980 22293 16983
rect 22244 16952 22293 16980
rect 22244 16940 22250 16952
rect 22281 16949 22293 16952
rect 22327 16949 22339 16983
rect 22281 16943 22339 16949
rect 22925 16983 22983 16989
rect 22925 16949 22937 16983
rect 22971 16980 22983 16983
rect 24670 16980 24676 16992
rect 22971 16952 24676 16980
rect 22971 16949 22983 16952
rect 22925 16943 22983 16949
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 29086 16940 29092 16992
rect 29144 16940 29150 16992
rect 33686 16940 33692 16992
rect 33744 16940 33750 16992
rect 1104 16890 43884 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 43884 16890
rect 1104 16816 43884 16838
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 17310 16776 17316 16788
rect 16531 16748 17316 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17586 16736 17592 16788
rect 17644 16736 17650 16788
rect 23566 16736 23572 16788
rect 23624 16736 23630 16788
rect 23934 16736 23940 16788
rect 23992 16776 23998 16788
rect 26326 16776 26332 16788
rect 23992 16748 26332 16776
rect 23992 16736 23998 16748
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 22152 16680 23428 16708
rect 22152 16668 22158 16680
rect 18414 16600 18420 16652
rect 18472 16600 18478 16652
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16640 18567 16643
rect 18598 16640 18604 16652
rect 18555 16612 18604 16640
rect 18555 16609 18567 16612
rect 18509 16603 18567 16609
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 20763 16612 21956 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 16942 16532 16948 16584
rect 17000 16532 17006 16584
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 18782 16532 18788 16584
rect 18840 16532 18846 16584
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16572 20591 16575
rect 20990 16572 20996 16584
rect 20579 16544 20996 16572
rect 20579 16541 20591 16544
rect 20533 16535 20591 16541
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 20806 16464 20812 16516
rect 20864 16464 20870 16516
rect 20898 16464 20904 16516
rect 20956 16464 20962 16516
rect 21928 16504 21956 16612
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16572 22063 16575
rect 22186 16572 22192 16584
rect 22051 16544 22192 16572
rect 22051 16541 22063 16544
rect 22005 16535 22063 16541
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22278 16532 22284 16584
rect 22336 16572 22342 16584
rect 22373 16575 22431 16581
rect 22373 16572 22385 16575
rect 22336 16544 22385 16572
rect 22336 16532 22342 16544
rect 22373 16541 22385 16544
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 22462 16532 22468 16584
rect 22520 16572 22526 16584
rect 23400 16581 23428 16680
rect 24872 16649 24900 16748
rect 26326 16736 26332 16748
rect 26384 16736 26390 16788
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27341 16779 27399 16785
rect 27341 16776 27353 16779
rect 27028 16748 27353 16776
rect 27028 16736 27034 16748
rect 27341 16745 27353 16748
rect 27387 16745 27399 16779
rect 27341 16739 27399 16745
rect 27525 16779 27583 16785
rect 27525 16745 27537 16779
rect 27571 16776 27583 16779
rect 28350 16776 28356 16788
rect 27571 16748 28356 16776
rect 27571 16745 27583 16748
rect 27525 16739 27583 16745
rect 28350 16736 28356 16748
rect 28408 16736 28414 16788
rect 28626 16736 28632 16788
rect 28684 16736 28690 16788
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16609 24915 16643
rect 27614 16640 27620 16652
rect 24857 16603 24915 16609
rect 27448 16612 27620 16640
rect 22649 16575 22707 16581
rect 22649 16572 22661 16575
rect 22520 16544 22661 16572
rect 22520 16532 22526 16544
rect 22649 16541 22661 16544
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23566 16532 23572 16584
rect 23624 16532 23630 16584
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 25113 16575 25171 16581
rect 25113 16572 25125 16575
rect 24728 16544 25125 16572
rect 24728 16532 24734 16544
rect 25113 16541 25125 16544
rect 25159 16541 25171 16575
rect 27448 16572 27476 16612
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 28258 16600 28264 16652
rect 28316 16600 28322 16652
rect 28534 16600 28540 16652
rect 28592 16640 28598 16652
rect 29825 16643 29883 16649
rect 29825 16640 29837 16643
rect 28592 16612 29837 16640
rect 28592 16600 28598 16612
rect 29825 16609 29837 16612
rect 29871 16609 29883 16643
rect 29825 16603 29883 16609
rect 31110 16600 31116 16652
rect 31168 16640 31174 16652
rect 31849 16643 31907 16649
rect 31849 16640 31861 16643
rect 31168 16612 31861 16640
rect 31168 16600 31174 16612
rect 31849 16609 31861 16612
rect 31895 16609 31907 16643
rect 31849 16603 31907 16609
rect 32306 16600 32312 16652
rect 32364 16600 32370 16652
rect 38194 16600 38200 16652
rect 38252 16640 38258 16652
rect 38289 16643 38347 16649
rect 38289 16640 38301 16643
rect 38252 16612 38301 16640
rect 38252 16600 38258 16612
rect 38289 16609 38301 16612
rect 38335 16609 38347 16643
rect 38289 16603 38347 16609
rect 38378 16600 38384 16652
rect 38436 16600 38442 16652
rect 41506 16600 41512 16652
rect 41564 16600 41570 16652
rect 25113 16535 25171 16541
rect 26252 16544 27476 16572
rect 21928 16476 22094 16504
rect 22066 16436 22094 16476
rect 22646 16436 22652 16448
rect 22066 16408 22652 16436
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 26252 16445 26280 16544
rect 27522 16532 27528 16584
rect 27580 16532 27586 16584
rect 30650 16532 30656 16584
rect 30708 16532 30714 16584
rect 31297 16575 31355 16581
rect 31297 16541 31309 16575
rect 31343 16572 31355 16575
rect 31754 16572 31760 16584
rect 31343 16544 31760 16572
rect 31343 16541 31355 16544
rect 31297 16535 31355 16541
rect 31754 16532 31760 16544
rect 31812 16532 31818 16584
rect 32030 16532 32036 16584
rect 32088 16532 32094 16584
rect 32398 16532 32404 16584
rect 32456 16532 32462 16584
rect 34514 16532 34520 16584
rect 34572 16572 34578 16584
rect 35621 16575 35679 16581
rect 35621 16572 35633 16575
rect 34572 16544 35633 16572
rect 34572 16532 34578 16544
rect 35621 16541 35633 16544
rect 35667 16541 35679 16575
rect 35621 16535 35679 16541
rect 35802 16532 35808 16584
rect 35860 16532 35866 16584
rect 35894 16532 35900 16584
rect 35952 16532 35958 16584
rect 35989 16575 36047 16581
rect 35989 16541 36001 16575
rect 36035 16572 36047 16575
rect 36354 16572 36360 16584
rect 36035 16544 36360 16572
rect 36035 16541 36047 16544
rect 35989 16535 36047 16541
rect 36354 16532 36360 16544
rect 36412 16532 36418 16584
rect 27157 16507 27215 16513
rect 27157 16473 27169 16507
rect 27203 16504 27215 16507
rect 27540 16504 27568 16532
rect 27203 16476 27568 16504
rect 28077 16507 28135 16513
rect 27203 16473 27215 16476
rect 27157 16467 27215 16473
rect 28077 16473 28089 16507
rect 28123 16504 28135 16507
rect 29086 16504 29092 16516
rect 28123 16476 29092 16504
rect 28123 16473 28135 16476
rect 28077 16467 28135 16473
rect 29086 16464 29092 16476
rect 29144 16504 29150 16516
rect 30190 16504 30196 16516
rect 29144 16476 30196 16504
rect 29144 16464 29150 16476
rect 30190 16464 30196 16476
rect 30248 16464 30254 16516
rect 31389 16507 31447 16513
rect 31389 16473 31401 16507
rect 31435 16504 31447 16507
rect 31662 16504 31668 16516
rect 31435 16476 31668 16504
rect 31435 16473 31447 16476
rect 31389 16467 31447 16473
rect 31662 16464 31668 16476
rect 31720 16464 31726 16516
rect 38197 16507 38255 16513
rect 38197 16473 38209 16507
rect 38243 16504 38255 16507
rect 38470 16504 38476 16516
rect 38243 16476 38476 16504
rect 38243 16473 38255 16476
rect 38197 16467 38255 16473
rect 38470 16464 38476 16476
rect 38528 16464 38534 16516
rect 40494 16464 40500 16516
rect 40552 16504 40558 16516
rect 41242 16507 41300 16513
rect 41242 16504 41254 16507
rect 40552 16476 41254 16504
rect 40552 16464 40558 16476
rect 41242 16473 41254 16476
rect 41288 16473 41300 16507
rect 41242 16467 41300 16473
rect 26237 16439 26295 16445
rect 26237 16405 26249 16439
rect 26283 16405 26295 16439
rect 26237 16399 26295 16405
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 27357 16439 27415 16445
rect 27357 16436 27369 16439
rect 27120 16408 27369 16436
rect 27120 16396 27126 16408
rect 27357 16405 27369 16408
rect 27403 16405 27415 16439
rect 27357 16399 27415 16405
rect 28166 16396 28172 16448
rect 28224 16396 28230 16448
rect 36265 16439 36323 16445
rect 36265 16405 36277 16439
rect 36311 16436 36323 16439
rect 37458 16436 37464 16448
rect 36311 16408 37464 16436
rect 36311 16405 36323 16408
rect 36265 16399 36323 16405
rect 37458 16396 37464 16408
rect 37516 16396 37522 16448
rect 37734 16396 37740 16448
rect 37792 16436 37798 16448
rect 37829 16439 37887 16445
rect 37829 16436 37841 16439
rect 37792 16408 37841 16436
rect 37792 16396 37798 16408
rect 37829 16405 37841 16408
rect 37875 16405 37887 16439
rect 37829 16399 37887 16405
rect 40126 16396 40132 16448
rect 40184 16396 40190 16448
rect 1104 16346 43884 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 43884 16346
rect 1104 16272 43884 16294
rect 22557 16235 22615 16241
rect 22557 16201 22569 16235
rect 22603 16232 22615 16235
rect 23566 16232 23572 16244
rect 22603 16204 23572 16232
rect 22603 16201 22615 16204
rect 22557 16195 22615 16201
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 27430 16192 27436 16244
rect 27488 16232 27494 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 27488 16204 27629 16232
rect 27488 16192 27494 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 27617 16195 27675 16201
rect 29917 16235 29975 16241
rect 29917 16201 29929 16235
rect 29963 16232 29975 16235
rect 30006 16232 30012 16244
rect 29963 16204 30012 16232
rect 29963 16201 29975 16204
rect 29917 16195 29975 16201
rect 30006 16192 30012 16204
rect 30064 16192 30070 16244
rect 30285 16235 30343 16241
rect 30285 16201 30297 16235
rect 30331 16232 30343 16235
rect 31110 16232 31116 16244
rect 30331 16204 31116 16232
rect 30331 16201 30343 16204
rect 30285 16195 30343 16201
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 31754 16192 31760 16244
rect 31812 16192 31818 16244
rect 37550 16192 37556 16244
rect 37608 16192 37614 16244
rect 38194 16192 38200 16244
rect 38252 16232 38258 16244
rect 40037 16235 40095 16241
rect 40037 16232 40049 16235
rect 38252 16204 40049 16232
rect 38252 16192 38258 16204
rect 40037 16201 40049 16204
rect 40083 16201 40095 16235
rect 40037 16195 40095 16201
rect 40494 16192 40500 16244
rect 40552 16192 40558 16244
rect 22186 16124 22192 16176
rect 22244 16124 22250 16176
rect 22370 16124 22376 16176
rect 22428 16173 22434 16176
rect 22428 16167 22447 16173
rect 22435 16133 22447 16167
rect 22428 16127 22447 16133
rect 22428 16124 22434 16127
rect 22646 16124 22652 16176
rect 22704 16164 22710 16176
rect 23201 16167 23259 16173
rect 23201 16164 23213 16167
rect 22704 16136 23213 16164
rect 22704 16124 22710 16136
rect 23201 16133 23213 16136
rect 23247 16133 23259 16167
rect 23201 16127 23259 16133
rect 23382 16124 23388 16176
rect 23440 16124 23446 16176
rect 25501 16167 25559 16173
rect 25501 16133 25513 16167
rect 25547 16164 25559 16167
rect 29454 16164 29460 16176
rect 25547 16136 29460 16164
rect 25547 16133 25559 16136
rect 25501 16127 25559 16133
rect 29454 16124 29460 16136
rect 29512 16124 29518 16176
rect 30190 16124 30196 16176
rect 30248 16164 30254 16176
rect 35710 16164 35716 16176
rect 30248 16136 31340 16164
rect 30248 16124 30254 16136
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18414 16096 18420 16108
rect 18371 16068 18420 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18506 16056 18512 16108
rect 18564 16056 18570 16108
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20530 16096 20536 16108
rect 20036 16068 20536 16096
rect 20036 16056 20042 16068
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20864 16068 20913 16096
rect 20864 16056 20870 16068
rect 20901 16065 20913 16068
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 27522 16056 27528 16108
rect 27580 16056 27586 16108
rect 30282 16096 30288 16108
rect 27816 16068 30288 16096
rect 23842 15988 23848 16040
rect 23900 15988 23906 16040
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 27816 16037 27844 16068
rect 30282 16056 30288 16068
rect 30340 16096 30346 16108
rect 30340 16068 30512 16096
rect 30340 16056 30346 16068
rect 27801 16031 27859 16037
rect 27801 15997 27813 16031
rect 27847 15997 27859 16031
rect 27801 15991 27859 15997
rect 29914 15988 29920 16040
rect 29972 16028 29978 16040
rect 30484 16037 30512 16068
rect 31110 16056 31116 16108
rect 31168 16056 31174 16108
rect 31312 16105 31340 16136
rect 34992 16136 35716 16164
rect 31297 16099 31355 16105
rect 31297 16065 31309 16099
rect 31343 16065 31355 16099
rect 31297 16059 31355 16065
rect 31386 16056 31392 16108
rect 31444 16056 31450 16108
rect 33318 16105 33324 16108
rect 31481 16099 31539 16105
rect 31481 16065 31493 16099
rect 31527 16065 31539 16099
rect 31481 16059 31539 16065
rect 33312 16059 33324 16105
rect 30377 16031 30435 16037
rect 30377 16028 30389 16031
rect 29972 16000 30389 16028
rect 29972 15988 29978 16000
rect 30377 15997 30389 16000
rect 30423 15997 30435 16031
rect 30377 15991 30435 15997
rect 30469 16031 30527 16037
rect 30469 15997 30481 16031
rect 30515 15997 30527 16031
rect 30469 15991 30527 15997
rect 30098 15920 30104 15972
rect 30156 15960 30162 15972
rect 31496 15960 31524 16059
rect 33318 16056 33324 16059
rect 33376 16056 33382 16108
rect 34992 16105 35020 16136
rect 35710 16124 35716 16136
rect 35768 16124 35774 16176
rect 35250 16105 35256 16108
rect 34977 16099 35035 16105
rect 34977 16065 34989 16099
rect 35023 16065 35035 16099
rect 34977 16059 35035 16065
rect 35244 16059 35256 16105
rect 35250 16056 35256 16059
rect 35308 16056 35314 16108
rect 37458 16056 37464 16108
rect 37516 16056 37522 16108
rect 38286 16056 38292 16108
rect 38344 16056 38350 16108
rect 38933 16099 38991 16105
rect 38933 16065 38945 16099
rect 38979 16096 38991 16099
rect 40126 16096 40132 16108
rect 38979 16068 40132 16096
rect 38979 16065 38991 16068
rect 38933 16059 38991 16065
rect 40126 16056 40132 16068
rect 40184 16056 40190 16108
rect 33042 15988 33048 16040
rect 33100 15988 33106 16040
rect 38470 15988 38476 16040
rect 38528 15988 38534 16040
rect 38654 15988 38660 16040
rect 38712 15988 38718 16040
rect 38838 15988 38844 16040
rect 38896 16028 38902 16040
rect 39853 16031 39911 16037
rect 39853 16028 39865 16031
rect 38896 16000 39865 16028
rect 38896 15988 38902 16000
rect 39853 15997 39865 16000
rect 39899 15997 39911 16031
rect 39853 15991 39911 15997
rect 30156 15932 31524 15960
rect 30156 15920 30162 15932
rect 19981 15895 20039 15901
rect 19981 15861 19993 15895
rect 20027 15892 20039 15895
rect 20898 15892 20904 15904
rect 20027 15864 20904 15892
rect 20027 15861 20039 15864
rect 19981 15855 20039 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21082 15852 21088 15904
rect 21140 15852 21146 15904
rect 22278 15852 22284 15904
rect 22336 15892 22342 15904
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 22336 15864 22385 15892
rect 22336 15852 22342 15864
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 23017 15895 23075 15901
rect 23017 15892 23029 15895
rect 22796 15864 23029 15892
rect 22796 15852 22802 15864
rect 23017 15861 23029 15864
rect 23063 15861 23075 15895
rect 23017 15855 23075 15861
rect 27154 15852 27160 15904
rect 27212 15852 27218 15904
rect 34422 15852 34428 15904
rect 34480 15852 34486 15904
rect 36354 15852 36360 15904
rect 36412 15852 36418 15904
rect 43346 15852 43352 15904
rect 43404 15852 43410 15904
rect 1104 15802 43884 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 43884 15802
rect 1104 15728 43884 15750
rect 22370 15688 22376 15700
rect 20732 15660 22376 15688
rect 20732 15629 20760 15660
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 27522 15648 27528 15700
rect 27580 15688 27586 15700
rect 27617 15691 27675 15697
rect 27617 15688 27629 15691
rect 27580 15660 27629 15688
rect 27580 15648 27586 15660
rect 27617 15657 27629 15660
rect 27663 15657 27675 15691
rect 27617 15651 27675 15657
rect 34333 15691 34391 15697
rect 34333 15657 34345 15691
rect 34379 15688 34391 15691
rect 34514 15688 34520 15700
rect 34379 15660 34520 15688
rect 34379 15657 34391 15660
rect 34333 15651 34391 15657
rect 34514 15648 34520 15660
rect 34572 15648 34578 15700
rect 35342 15648 35348 15700
rect 35400 15688 35406 15700
rect 35437 15691 35495 15697
rect 35437 15688 35449 15691
rect 35400 15660 35449 15688
rect 35400 15648 35406 15660
rect 35437 15657 35449 15660
rect 35483 15657 35495 15691
rect 35437 15651 35495 15657
rect 38470 15648 38476 15700
rect 38528 15688 38534 15700
rect 38841 15691 38899 15697
rect 38841 15688 38853 15691
rect 38528 15660 38853 15688
rect 38528 15648 38534 15660
rect 38841 15657 38853 15660
rect 38887 15657 38899 15691
rect 38841 15651 38899 15657
rect 20717 15623 20775 15629
rect 20717 15589 20729 15623
rect 20763 15589 20775 15623
rect 20717 15583 20775 15589
rect 20898 15580 20904 15632
rect 20956 15620 20962 15632
rect 24118 15620 24124 15632
rect 20956 15592 24124 15620
rect 20956 15580 20962 15592
rect 24118 15580 24124 15592
rect 24176 15580 24182 15632
rect 18049 15555 18107 15561
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 22833 15555 22891 15561
rect 18095 15524 18644 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 18616 15496 18644 15524
rect 22833 15521 22845 15555
rect 22879 15552 22891 15555
rect 23661 15555 23719 15561
rect 23661 15552 23673 15555
rect 22879 15524 23673 15552
rect 22879 15521 22891 15524
rect 22833 15515 22891 15521
rect 23661 15521 23673 15524
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 29914 15552 29920 15564
rect 29052 15524 29920 15552
rect 29052 15512 29058 15524
rect 29914 15512 29920 15524
rect 29972 15552 29978 15564
rect 30193 15555 30251 15561
rect 30193 15552 30205 15555
rect 29972 15524 30205 15552
rect 29972 15512 29978 15524
rect 30193 15521 30205 15524
rect 30239 15521 30251 15555
rect 30193 15515 30251 15521
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15552 30343 15555
rect 30466 15552 30472 15564
rect 30331 15524 30472 15552
rect 30331 15521 30343 15524
rect 30285 15515 30343 15521
rect 30466 15512 30472 15524
rect 30524 15512 30530 15564
rect 35342 15552 35348 15564
rect 31726 15524 35348 15552
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 18506 15484 18512 15496
rect 18371 15456 18512 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 18598 15444 18604 15496
rect 18656 15444 18662 15496
rect 18782 15444 18788 15496
rect 18840 15444 18846 15496
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20404 15456 20545 15484
rect 20404 15444 20410 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20898 15444 20904 15496
rect 20956 15444 20962 15496
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 22554 15444 22560 15496
rect 22612 15444 22618 15496
rect 22738 15444 22744 15496
rect 22796 15444 22802 15496
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 23569 15487 23627 15493
rect 23569 15484 23581 15487
rect 23440 15456 23581 15484
rect 23440 15444 23446 15456
rect 23569 15453 23581 15456
rect 23615 15453 23627 15487
rect 23569 15447 23627 15453
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15484 26295 15487
rect 26326 15484 26332 15496
rect 26283 15456 26332 15484
rect 26283 15453 26295 15456
rect 26237 15447 26295 15453
rect 26326 15444 26332 15456
rect 26384 15484 26390 15496
rect 28718 15484 28724 15496
rect 26384 15456 28724 15484
rect 26384 15444 26390 15456
rect 28718 15444 28724 15456
rect 28776 15444 28782 15496
rect 30098 15444 30104 15496
rect 30156 15444 30162 15496
rect 22094 15376 22100 15428
rect 22152 15376 22158 15428
rect 24302 15376 24308 15428
rect 24360 15416 24366 15428
rect 25314 15416 25320 15428
rect 24360 15388 25320 15416
rect 24360 15376 24366 15388
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 26504 15419 26562 15425
rect 26504 15385 26516 15419
rect 26550 15416 26562 15419
rect 27154 15416 27160 15428
rect 26550 15388 27160 15416
rect 26550 15385 26562 15388
rect 26504 15379 26562 15385
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 31386 15416 31392 15428
rect 29656 15388 31392 15416
rect 18785 15351 18843 15357
rect 18785 15317 18797 15351
rect 18831 15348 18843 15351
rect 19426 15348 19432 15360
rect 18831 15320 19432 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 25332 15348 25360 15376
rect 29656 15348 29684 15388
rect 31386 15376 31392 15388
rect 31444 15416 31450 15428
rect 31726 15416 31754 15524
rect 32600 15493 32628 15524
rect 35342 15512 35348 15524
rect 35400 15512 35406 15564
rect 35710 15512 35716 15564
rect 35768 15552 35774 15564
rect 35989 15555 36047 15561
rect 35989 15552 36001 15555
rect 35768 15524 36001 15552
rect 35768 15512 35774 15524
rect 35989 15521 36001 15524
rect 36035 15521 36047 15555
rect 35989 15515 36047 15521
rect 32585 15487 32643 15493
rect 32585 15453 32597 15487
rect 32631 15453 32643 15487
rect 32585 15447 32643 15453
rect 32950 15444 32956 15496
rect 33008 15444 33014 15496
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15484 34207 15487
rect 34422 15484 34428 15496
rect 34195 15456 34428 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 34422 15444 34428 15456
rect 34480 15444 34486 15496
rect 35526 15444 35532 15496
rect 35584 15484 35590 15496
rect 37734 15493 37740 15496
rect 37461 15487 37519 15493
rect 37461 15484 37473 15487
rect 35584 15456 37473 15484
rect 35584 15444 35590 15456
rect 37461 15453 37473 15456
rect 37507 15453 37519 15487
rect 37728 15484 37740 15493
rect 37695 15456 37740 15484
rect 37461 15447 37519 15453
rect 37728 15447 37740 15456
rect 37734 15444 37740 15447
rect 37792 15444 37798 15496
rect 31444 15388 31754 15416
rect 31444 15376 31450 15388
rect 33962 15376 33968 15428
rect 34020 15376 34026 15428
rect 35805 15419 35863 15425
rect 35805 15385 35817 15419
rect 35851 15416 35863 15419
rect 36354 15416 36360 15428
rect 35851 15388 36360 15416
rect 35851 15385 35863 15388
rect 35805 15379 35863 15385
rect 36354 15376 36360 15388
rect 36412 15376 36418 15428
rect 25332 15320 29684 15348
rect 29730 15308 29736 15360
rect 29788 15308 29794 15360
rect 32030 15308 32036 15360
rect 32088 15308 32094 15360
rect 33134 15308 33140 15360
rect 33192 15348 33198 15360
rect 35897 15351 35955 15357
rect 35897 15348 35909 15351
rect 33192 15320 35909 15348
rect 33192 15308 33198 15320
rect 35897 15317 35909 15320
rect 35943 15348 35955 15351
rect 38194 15348 38200 15360
rect 35943 15320 38200 15348
rect 35943 15317 35955 15320
rect 35897 15311 35955 15317
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 43884 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 43884 15258
rect 1104 15184 43884 15206
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18104 15116 18245 15144
rect 18104 15104 18110 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 22097 15147 22155 15153
rect 22097 15113 22109 15147
rect 22143 15144 22155 15147
rect 22278 15144 22284 15156
rect 22143 15116 22284 15144
rect 22143 15113 22155 15116
rect 22097 15107 22155 15113
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 29917 15147 29975 15153
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 30098 15144 30104 15156
rect 29963 15116 30104 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 30098 15104 30104 15116
rect 30156 15104 30162 15156
rect 30745 15147 30803 15153
rect 30745 15113 30757 15147
rect 30791 15144 30803 15147
rect 31110 15144 31116 15156
rect 30791 15116 31116 15144
rect 30791 15113 30803 15116
rect 30745 15107 30803 15113
rect 31110 15104 31116 15116
rect 31168 15104 31174 15156
rect 33042 15104 33048 15156
rect 33100 15144 33106 15156
rect 35526 15144 35532 15156
rect 33100 15116 35532 15144
rect 33100 15104 33106 15116
rect 35526 15104 35532 15116
rect 35584 15104 35590 15156
rect 41141 15147 41199 15153
rect 41141 15113 41153 15147
rect 41187 15113 41199 15147
rect 41141 15107 41199 15113
rect 19168 15048 22094 15076
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 19168 15017 19196 15048
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 14977 19027 15011
rect 18969 14971 19027 14977
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 18414 14940 18420 14952
rect 17175 14912 18420 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18984 14872 19012 14971
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20364 15017 20392 15048
rect 22066 15020 22094 15048
rect 23290 15036 23296 15088
rect 23348 15076 23354 15088
rect 23658 15076 23664 15088
rect 23348 15048 23664 15076
rect 23348 15036 23354 15048
rect 23658 15036 23664 15048
rect 23716 15076 23722 15088
rect 28804 15079 28862 15085
rect 23716 15048 24072 15076
rect 23716 15036 23722 15048
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 15008 20683 15011
rect 20714 15008 20720 15020
rect 20671 14980 20720 15008
rect 20671 14977 20683 14980
rect 20625 14971 20683 14977
rect 20714 14968 20720 14980
rect 20772 15008 20778 15020
rect 21082 15008 21088 15020
rect 20772 14980 21088 15008
rect 20772 14968 20778 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 22066 14980 22100 15020
rect 22094 14968 22100 14980
rect 22152 15008 22158 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22152 14980 22293 15008
rect 22152 14968 22158 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 20441 14943 20499 14949
rect 20441 14940 20453 14943
rect 19484 14912 20453 14940
rect 19484 14900 19490 14912
rect 20441 14909 20453 14912
rect 20487 14909 20499 14943
rect 22388 14940 22416 14971
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22612 14980 22661 15008
rect 22612 14968 22618 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 23106 14968 23112 15020
rect 23164 15008 23170 15020
rect 24044 15017 24072 15048
rect 28804 15045 28816 15079
rect 28850 15076 28862 15079
rect 29730 15076 29736 15088
rect 28850 15048 29736 15076
rect 28850 15045 28862 15048
rect 28804 15039 28862 15045
rect 29730 15036 29736 15048
rect 29788 15036 29794 15088
rect 33689 15079 33747 15085
rect 33689 15045 33701 15079
rect 33735 15076 33747 15079
rect 34422 15076 34428 15088
rect 33735 15048 34428 15076
rect 33735 15045 33747 15048
rect 33689 15039 33747 15045
rect 34422 15036 34428 15048
rect 34480 15036 34486 15088
rect 39114 15076 39120 15088
rect 38948 15048 39120 15076
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23164 14980 23857 15008
rect 23164 14968 23170 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 28534 14968 28540 15020
rect 28592 14968 28598 15020
rect 30377 15011 30435 15017
rect 30377 14977 30389 15011
rect 30423 14977 30435 15011
rect 30377 14971 30435 14977
rect 20441 14903 20499 14909
rect 22066 14912 22416 14940
rect 18984 14844 20208 14872
rect 20180 14816 20208 14844
rect 20346 14832 20352 14884
rect 20404 14832 20410 14884
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 18969 14807 19027 14813
rect 18969 14804 18981 14807
rect 18932 14776 18981 14804
rect 18932 14764 18938 14776
rect 18969 14773 18981 14776
rect 19015 14773 19027 14807
rect 18969 14767 19027 14773
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 22066 14804 22094 14912
rect 29730 14900 29736 14952
rect 29788 14940 29794 14952
rect 30392 14940 30420 14971
rect 30558 14968 30564 15020
rect 30616 14968 30622 15020
rect 31662 14968 31668 15020
rect 31720 15008 31726 15020
rect 32401 15011 32459 15017
rect 32401 15008 32413 15011
rect 31720 14980 32413 15008
rect 31720 14968 31726 14980
rect 32401 14977 32413 14980
rect 32447 14977 32459 15011
rect 32401 14971 32459 14977
rect 33134 14968 33140 15020
rect 33192 15008 33198 15020
rect 33781 15011 33839 15017
rect 33781 15008 33793 15011
rect 33192 14980 33793 15008
rect 33192 14968 33198 14980
rect 33781 14977 33793 14980
rect 33827 14977 33839 15011
rect 33781 14971 33839 14977
rect 34514 14968 34520 15020
rect 34572 15008 34578 15020
rect 35621 15011 35679 15017
rect 35621 15008 35633 15011
rect 34572 14980 35633 15008
rect 34572 14968 34578 14980
rect 35621 14977 35633 14980
rect 35667 14977 35679 15011
rect 35621 14971 35679 14977
rect 35802 14968 35808 15020
rect 35860 14968 35866 15020
rect 35894 14968 35900 15020
rect 35952 14968 35958 15020
rect 35989 15011 36047 15017
rect 35989 14977 36001 15011
rect 36035 14977 36047 15011
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 35989 14971 36047 14977
rect 36280 14980 37473 15008
rect 29788 14912 30420 14940
rect 29788 14900 29794 14912
rect 32306 14900 32312 14952
rect 32364 14900 32370 14952
rect 33873 14943 33931 14949
rect 33873 14909 33885 14943
rect 33919 14909 33931 14943
rect 36004 14940 36032 14971
rect 36280 14949 36308 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 38010 14968 38016 15020
rect 38068 14968 38074 15020
rect 38286 15008 38292 15020
rect 38120 14980 38292 15008
rect 33873 14903 33931 14909
rect 35912 14912 36032 14940
rect 36265 14943 36323 14949
rect 22557 14875 22615 14881
rect 22557 14841 22569 14875
rect 22603 14872 22615 14875
rect 23382 14872 23388 14884
rect 22603 14844 23388 14872
rect 22603 14841 22615 14844
rect 22557 14835 22615 14841
rect 23382 14832 23388 14844
rect 23440 14832 23446 14884
rect 32030 14832 32036 14884
rect 32088 14872 32094 14884
rect 32088 14844 33272 14872
rect 32088 14832 32094 14844
rect 20220 14776 22094 14804
rect 20220 14764 20226 14776
rect 23934 14764 23940 14816
rect 23992 14764 23998 14816
rect 28810 14764 28816 14816
rect 28868 14804 28874 14816
rect 31202 14804 31208 14816
rect 28868 14776 31208 14804
rect 28868 14764 28874 14776
rect 31202 14764 31208 14776
rect 31260 14804 31266 14816
rect 32585 14807 32643 14813
rect 32585 14804 32597 14807
rect 31260 14776 32597 14804
rect 31260 14764 31266 14776
rect 32585 14773 32597 14776
rect 32631 14804 32643 14807
rect 33134 14804 33140 14816
rect 32631 14776 33140 14804
rect 32631 14773 32643 14776
rect 32585 14767 32643 14773
rect 33134 14764 33140 14776
rect 33192 14764 33198 14816
rect 33244 14804 33272 14844
rect 33318 14832 33324 14884
rect 33376 14832 33382 14884
rect 33410 14832 33416 14884
rect 33468 14872 33474 14884
rect 33888 14872 33916 14903
rect 35912 14884 35940 14912
rect 36265 14909 36277 14943
rect 36311 14909 36323 14943
rect 36265 14903 36323 14909
rect 33468 14844 33916 14872
rect 33468 14832 33474 14844
rect 35894 14832 35900 14884
rect 35952 14832 35958 14884
rect 38120 14804 38148 14980
rect 38286 14968 38292 14980
rect 38344 14968 38350 15020
rect 38654 14968 38660 15020
rect 38712 14968 38718 15020
rect 38948 15017 38976 15048
rect 39114 15036 39120 15048
rect 39172 15076 39178 15088
rect 41156 15076 41184 15107
rect 39172 15048 41184 15076
rect 39172 15036 39178 15048
rect 38933 15011 38991 15017
rect 38933 14977 38945 15011
rect 38979 14977 38991 15011
rect 38933 14971 38991 14977
rect 39482 14968 39488 15020
rect 39540 15008 39546 15020
rect 40017 15011 40075 15017
rect 40017 15008 40029 15011
rect 39540 14980 40029 15008
rect 39540 14968 39546 14980
rect 40017 14977 40029 14980
rect 40063 14977 40075 15011
rect 40017 14971 40075 14977
rect 38470 14900 38476 14952
rect 38528 14900 38534 14952
rect 39758 14900 39764 14952
rect 39816 14900 39822 14952
rect 33244 14776 38148 14804
rect 1104 14714 43884 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 43884 14714
rect 1104 14640 43884 14662
rect 18414 14560 18420 14612
rect 18472 14560 18478 14612
rect 23569 14603 23627 14609
rect 23569 14569 23581 14603
rect 23615 14600 23627 14603
rect 27798 14600 27804 14612
rect 23615 14572 27804 14600
rect 23615 14569 23627 14572
rect 23569 14563 23627 14569
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 31573 14603 31631 14609
rect 31573 14569 31585 14603
rect 31619 14600 31631 14603
rect 33318 14600 33324 14612
rect 31619 14572 33324 14600
rect 31619 14569 31631 14572
rect 31573 14563 31631 14569
rect 18601 14535 18659 14541
rect 18601 14501 18613 14535
rect 18647 14532 18659 14535
rect 20346 14532 20352 14544
rect 18647 14504 20352 14532
rect 18647 14501 18659 14504
rect 18601 14495 18659 14501
rect 20346 14492 20352 14504
rect 20404 14492 20410 14544
rect 27062 14492 27068 14544
rect 27120 14492 27126 14544
rect 27338 14492 27344 14544
rect 27396 14532 27402 14544
rect 31588 14532 31616 14563
rect 33318 14560 33324 14572
rect 33376 14560 33382 14612
rect 33689 14603 33747 14609
rect 33689 14569 33701 14603
rect 33735 14600 33747 14603
rect 33778 14600 33784 14612
rect 33735 14572 33784 14600
rect 33735 14569 33747 14572
rect 33689 14563 33747 14569
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 39482 14560 39488 14612
rect 39540 14560 39546 14612
rect 27396 14504 31616 14532
rect 33520 14504 38884 14532
rect 27396 14492 27402 14504
rect 18874 14424 18880 14476
rect 18932 14424 18938 14476
rect 22002 14424 22008 14476
rect 22060 14424 22066 14476
rect 25590 14424 25596 14476
rect 25648 14464 25654 14476
rect 27080 14464 27108 14492
rect 28552 14473 28580 14504
rect 28537 14467 28595 14473
rect 25648 14436 27384 14464
rect 25648 14424 25654 14436
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19484 14368 19717 14396
rect 19484 14356 19490 14368
rect 19705 14365 19717 14368
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14396 20591 14399
rect 20714 14396 20720 14408
rect 20579 14368 20720 14396
rect 20579 14365 20591 14368
rect 20533 14359 20591 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 22281 14399 22339 14405
rect 22281 14396 22293 14399
rect 22066 14368 22293 14396
rect 21266 14328 21272 14340
rect 21206 14300 21272 14328
rect 21266 14288 21272 14300
rect 21324 14328 21330 14340
rect 22066 14328 22094 14368
rect 22281 14365 22293 14368
rect 22327 14365 22339 14399
rect 22281 14359 22339 14365
rect 23842 14356 23848 14408
rect 23900 14396 23906 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 23900 14368 24593 14396
rect 23900 14356 23906 14368
rect 24581 14365 24593 14368
rect 24627 14396 24639 14399
rect 26142 14396 26148 14408
rect 24627 14368 26148 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 27062 14356 27068 14408
rect 27120 14356 27126 14408
rect 27356 14405 27384 14436
rect 28537 14433 28549 14467
rect 28583 14433 28595 14467
rect 30558 14464 30564 14476
rect 28537 14427 28595 14433
rect 28828 14436 30564 14464
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14396 27399 14399
rect 27798 14396 27804 14408
rect 27387 14368 27804 14396
rect 27387 14365 27399 14368
rect 27341 14359 27399 14365
rect 27798 14356 27804 14368
rect 27856 14356 27862 14408
rect 28828 14405 28856 14436
rect 30558 14424 30564 14436
rect 30616 14424 30622 14476
rect 31128 14436 31340 14464
rect 28813 14399 28871 14405
rect 28813 14365 28825 14399
rect 28859 14365 28871 14399
rect 28813 14359 28871 14365
rect 29730 14356 29736 14408
rect 29788 14356 29794 14408
rect 30009 14399 30067 14405
rect 30009 14396 30021 14399
rect 29840 14368 30021 14396
rect 21324 14300 22094 14328
rect 24848 14331 24906 14337
rect 21324 14288 21330 14300
rect 24848 14297 24860 14331
rect 24894 14328 24906 14331
rect 25130 14328 25136 14340
rect 24894 14300 25136 14328
rect 24894 14297 24906 14300
rect 24848 14291 24906 14297
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 26970 14328 26976 14340
rect 25424 14300 26976 14328
rect 23658 14220 23664 14272
rect 23716 14260 23722 14272
rect 25424 14260 25452 14300
rect 26970 14288 26976 14300
rect 27028 14328 27034 14340
rect 27249 14331 27307 14337
rect 27249 14328 27261 14331
rect 27028 14300 27261 14328
rect 27028 14288 27034 14300
rect 27249 14297 27261 14300
rect 27295 14297 27307 14331
rect 27249 14291 27307 14297
rect 28721 14331 28779 14337
rect 28721 14297 28733 14331
rect 28767 14328 28779 14331
rect 28994 14328 29000 14340
rect 28767 14300 29000 14328
rect 28767 14297 28779 14300
rect 28721 14291 28779 14297
rect 28994 14288 29000 14300
rect 29052 14288 29058 14340
rect 29840 14328 29868 14368
rect 30009 14365 30021 14368
rect 30055 14396 30067 14399
rect 31128 14396 31156 14436
rect 30055 14368 31156 14396
rect 31205 14399 31263 14405
rect 30055 14365 30067 14368
rect 30009 14359 30067 14365
rect 31205 14365 31217 14399
rect 31251 14365 31263 14399
rect 31312 14396 31340 14436
rect 31409 14399 31467 14405
rect 31409 14396 31421 14399
rect 31312 14368 31421 14396
rect 31205 14359 31263 14365
rect 31409 14365 31421 14368
rect 31455 14396 31467 14399
rect 31662 14396 31668 14408
rect 31455 14368 31668 14396
rect 31455 14365 31467 14368
rect 31409 14359 31467 14365
rect 29104 14300 29868 14328
rect 23716 14232 25452 14260
rect 23716 14220 23722 14232
rect 25498 14220 25504 14272
rect 25556 14260 25562 14272
rect 25961 14263 26019 14269
rect 25961 14260 25973 14263
rect 25556 14232 25973 14260
rect 25556 14220 25562 14232
rect 25961 14229 25973 14232
rect 26007 14229 26019 14263
rect 25961 14223 26019 14229
rect 26602 14220 26608 14272
rect 26660 14260 26666 14272
rect 26881 14263 26939 14269
rect 26881 14260 26893 14263
rect 26660 14232 26893 14260
rect 26660 14220 26666 14232
rect 26881 14229 26893 14232
rect 26927 14229 26939 14263
rect 26881 14223 26939 14229
rect 27982 14220 27988 14272
rect 28040 14260 28046 14272
rect 29104 14260 29132 14300
rect 29914 14288 29920 14340
rect 29972 14328 29978 14340
rect 30190 14328 30196 14340
rect 29972 14300 30196 14328
rect 29972 14288 29978 14300
rect 30190 14288 30196 14300
rect 30248 14288 30254 14340
rect 30466 14288 30472 14340
rect 30524 14288 30530 14340
rect 28040 14232 29132 14260
rect 28040 14220 28046 14232
rect 29178 14220 29184 14272
rect 29236 14220 29242 14272
rect 31220 14260 31248 14359
rect 31662 14356 31668 14368
rect 31720 14356 31726 14408
rect 32309 14399 32367 14405
rect 32309 14365 32321 14399
rect 32355 14396 32367 14399
rect 33042 14396 33048 14408
rect 32355 14368 33048 14396
rect 32355 14365 32367 14368
rect 32309 14359 32367 14365
rect 33042 14356 33048 14368
rect 33100 14356 33106 14408
rect 33134 14356 33140 14408
rect 33192 14396 33198 14408
rect 33520 14396 33548 14504
rect 38856 14476 38884 14504
rect 35710 14424 35716 14476
rect 35768 14464 35774 14476
rect 36081 14467 36139 14473
rect 36081 14464 36093 14467
rect 35768 14436 36093 14464
rect 35768 14424 35774 14436
rect 36081 14433 36093 14436
rect 36127 14433 36139 14467
rect 36081 14427 36139 14433
rect 38838 14424 38844 14476
rect 38896 14424 38902 14476
rect 35986 14396 35992 14408
rect 33192 14368 33548 14396
rect 33704 14368 35992 14396
rect 33192 14356 33198 14368
rect 31297 14331 31355 14337
rect 31297 14297 31309 14331
rect 31343 14328 31355 14331
rect 31570 14328 31576 14340
rect 31343 14300 31576 14328
rect 31343 14297 31355 14300
rect 31297 14291 31355 14297
rect 31570 14288 31576 14300
rect 31628 14288 31634 14340
rect 32576 14331 32634 14337
rect 31726 14300 32536 14328
rect 31386 14260 31392 14272
rect 31220 14232 31392 14260
rect 31386 14220 31392 14232
rect 31444 14260 31450 14272
rect 31726 14260 31754 14300
rect 31444 14232 31754 14260
rect 32508 14260 32536 14300
rect 32576 14297 32588 14331
rect 32622 14328 32634 14331
rect 32766 14328 32772 14340
rect 32622 14300 32772 14328
rect 32622 14297 32634 14300
rect 32576 14291 32634 14297
rect 32766 14288 32772 14300
rect 32824 14288 32830 14340
rect 33704 14260 33732 14368
rect 35986 14356 35992 14368
rect 36044 14356 36050 14408
rect 39114 14356 39120 14408
rect 39172 14356 39178 14408
rect 39758 14356 39764 14408
rect 39816 14396 39822 14408
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 39816 14368 40049 14396
rect 39816 14356 39822 14368
rect 40037 14365 40049 14368
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 43346 14356 43352 14408
rect 43404 14356 43410 14408
rect 34422 14288 34428 14340
rect 34480 14328 34486 14340
rect 39025 14331 39083 14337
rect 39025 14328 39037 14331
rect 34480 14300 39037 14328
rect 34480 14288 34486 14300
rect 32508 14232 33732 14260
rect 31444 14220 31450 14232
rect 35434 14220 35440 14272
rect 35492 14260 35498 14272
rect 35529 14263 35587 14269
rect 35529 14260 35541 14263
rect 35492 14232 35541 14260
rect 35492 14220 35498 14232
rect 35529 14229 35541 14232
rect 35575 14229 35587 14263
rect 35529 14223 35587 14229
rect 35894 14220 35900 14272
rect 35952 14220 35958 14272
rect 36004 14269 36032 14300
rect 39025 14297 39037 14300
rect 39071 14328 39083 14331
rect 39942 14328 39948 14340
rect 39071 14300 39948 14328
rect 39071 14297 39083 14300
rect 39025 14291 39083 14297
rect 39942 14288 39948 14300
rect 40000 14288 40006 14340
rect 40304 14331 40362 14337
rect 40304 14297 40316 14331
rect 40350 14328 40362 14331
rect 40402 14328 40408 14340
rect 40350 14300 40408 14328
rect 40350 14297 40362 14300
rect 40304 14291 40362 14297
rect 40402 14288 40408 14300
rect 40460 14288 40466 14340
rect 35989 14263 36047 14269
rect 35989 14229 36001 14263
rect 36035 14229 36047 14263
rect 35989 14223 36047 14229
rect 41414 14220 41420 14272
rect 41472 14220 41478 14272
rect 1104 14170 43884 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 43884 14170
rect 1104 14096 43884 14118
rect 19705 14059 19763 14065
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 20162 14056 20168 14068
rect 19751 14028 20168 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 25498 14016 25504 14068
rect 25556 14016 25562 14068
rect 27062 14016 27068 14068
rect 27120 14056 27126 14068
rect 27522 14056 27528 14068
rect 27120 14028 27528 14056
rect 27120 14016 27126 14028
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 30101 14059 30159 14065
rect 30101 14025 30113 14059
rect 30147 14056 30159 14059
rect 30558 14056 30564 14068
rect 30147 14028 30564 14056
rect 30147 14025 30159 14028
rect 30101 14019 30159 14025
rect 30558 14016 30564 14028
rect 30616 14016 30622 14068
rect 32766 14016 32772 14068
rect 32824 14016 32830 14068
rect 33226 14016 33232 14068
rect 33284 14056 33290 14068
rect 34422 14056 34428 14068
rect 33284 14028 34428 14056
rect 33284 14016 33290 14028
rect 34422 14016 34428 14028
rect 34480 14016 34486 14068
rect 34514 14016 34520 14068
rect 34572 14016 34578 14068
rect 34716 14028 35664 14056
rect 23382 13948 23388 14000
rect 23440 13988 23446 14000
rect 23661 13991 23719 13997
rect 23661 13988 23673 13991
rect 23440 13960 23673 13988
rect 23440 13948 23446 13960
rect 23661 13957 23673 13960
rect 23707 13957 23719 13991
rect 23661 13951 23719 13957
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 19978 13920 19984 13932
rect 19935 13892 19984 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20714 13920 20720 13932
rect 20119 13892 20720 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 23474 13880 23480 13932
rect 23532 13880 23538 13932
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13920 23811 13923
rect 24762 13920 24768 13932
rect 23799 13892 24768 13920
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 24762 13880 24768 13892
rect 24820 13880 24826 13932
rect 25516 13920 25544 14016
rect 25593 13991 25651 13997
rect 25593 13957 25605 13991
rect 25639 13988 25651 13991
rect 26605 13991 26663 13997
rect 25639 13960 26556 13988
rect 25639 13957 25651 13960
rect 25593 13951 25651 13957
rect 26329 13923 26387 13929
rect 26329 13920 26341 13923
rect 25516 13892 26341 13920
rect 26329 13889 26341 13892
rect 26375 13889 26387 13923
rect 26528 13920 26556 13960
rect 26605 13957 26617 13991
rect 26651 13988 26663 13991
rect 28166 13988 28172 14000
rect 26651 13960 28172 13988
rect 26651 13957 26663 13960
rect 26605 13951 26663 13957
rect 28166 13948 28172 13960
rect 28224 13948 28230 14000
rect 28988 13991 29046 13997
rect 28988 13957 29000 13991
rect 29034 13988 29046 13991
rect 29178 13988 29184 14000
rect 29034 13960 29184 13988
rect 29034 13957 29046 13960
rect 28988 13951 29046 13957
rect 29178 13948 29184 13960
rect 29236 13948 29242 14000
rect 30282 13948 30288 14000
rect 30340 13988 30346 14000
rect 31205 13991 31263 13997
rect 31205 13988 31217 13991
rect 30340 13960 31217 13988
rect 30340 13948 30346 13960
rect 31205 13957 31217 13960
rect 31251 13957 31263 13991
rect 31205 13951 31263 13957
rect 33137 13991 33195 13997
rect 33137 13957 33149 13991
rect 33183 13988 33195 13991
rect 33778 13988 33784 14000
rect 33183 13960 33784 13988
rect 33183 13957 33195 13960
rect 33137 13951 33195 13957
rect 27430 13920 27436 13932
rect 26528 13892 27436 13920
rect 26329 13883 26387 13889
rect 27430 13880 27436 13892
rect 27488 13920 27494 13932
rect 27617 13923 27675 13929
rect 27617 13920 27629 13923
rect 27488 13892 27629 13920
rect 27488 13880 27494 13892
rect 27617 13889 27629 13892
rect 27663 13889 27675 13923
rect 27617 13883 27675 13889
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 19484 13824 20177 13852
rect 19484 13812 19490 13824
rect 20165 13821 20177 13824
rect 20211 13821 20223 13855
rect 20165 13815 20223 13821
rect 25685 13855 25743 13861
rect 25685 13821 25697 13855
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 25130 13744 25136 13796
rect 25188 13784 25194 13796
rect 25700 13784 25728 13815
rect 26602 13812 26608 13864
rect 26660 13812 26666 13864
rect 27338 13812 27344 13864
rect 27396 13852 27402 13864
rect 27709 13855 27767 13861
rect 27709 13852 27721 13855
rect 27396 13824 27721 13852
rect 27396 13812 27402 13824
rect 27709 13821 27721 13824
rect 27755 13821 27767 13855
rect 27709 13815 27767 13821
rect 28718 13812 28724 13864
rect 28776 13812 28782 13864
rect 31220 13852 31248 13951
rect 33778 13948 33784 13960
rect 33836 13988 33842 14000
rect 34333 13991 34391 13997
rect 34333 13988 34345 13991
rect 33836 13960 34345 13988
rect 33836 13948 33842 13960
rect 34333 13957 34345 13960
rect 34379 13957 34391 13991
rect 34333 13951 34391 13957
rect 31662 13880 31668 13932
rect 31720 13880 31726 13932
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13920 31815 13923
rect 32030 13920 32036 13932
rect 31803 13892 32036 13920
rect 31803 13889 31815 13892
rect 31757 13883 31815 13889
rect 32030 13880 32036 13892
rect 32088 13880 32094 13932
rect 33152 13892 33456 13920
rect 33152 13852 33180 13892
rect 31220 13824 33180 13852
rect 33318 13812 33324 13864
rect 33376 13812 33382 13864
rect 33428 13852 33456 13892
rect 33962 13880 33968 13932
rect 34020 13920 34026 13932
rect 34149 13923 34207 13929
rect 34149 13920 34161 13923
rect 34020 13892 34161 13920
rect 34020 13880 34026 13892
rect 34149 13889 34161 13892
rect 34195 13889 34207 13923
rect 34149 13883 34207 13889
rect 34716 13852 34744 14028
rect 35526 13988 35532 14000
rect 35176 13960 35532 13988
rect 34790 13880 34796 13932
rect 34848 13920 34854 13932
rect 35176 13929 35204 13960
rect 35526 13948 35532 13960
rect 35584 13948 35590 14000
rect 35636 13988 35664 14028
rect 35894 14016 35900 14068
rect 35952 14056 35958 14068
rect 36541 14059 36599 14065
rect 36541 14056 36553 14059
rect 35952 14028 36553 14056
rect 35952 14016 35958 14028
rect 36541 14025 36553 14028
rect 36587 14025 36599 14059
rect 36541 14019 36599 14025
rect 38470 14016 38476 14068
rect 38528 14056 38534 14068
rect 40037 14059 40095 14065
rect 40037 14056 40049 14059
rect 38528 14028 40049 14056
rect 38528 14016 38534 14028
rect 40037 14025 40049 14028
rect 40083 14025 40095 14059
rect 40037 14019 40095 14025
rect 38378 13988 38384 14000
rect 35636 13960 38384 13988
rect 38378 13948 38384 13960
rect 38436 13948 38442 14000
rect 39942 13948 39948 14000
rect 40000 13948 40006 14000
rect 40052 13988 40080 14019
rect 40402 14016 40408 14068
rect 40460 14016 40466 14068
rect 41414 13988 41420 14000
rect 40052 13960 41420 13988
rect 41414 13948 41420 13960
rect 41472 13948 41478 14000
rect 35434 13929 35440 13932
rect 35161 13923 35219 13929
rect 35161 13920 35173 13923
rect 34848 13892 35173 13920
rect 34848 13880 34854 13892
rect 35161 13889 35173 13892
rect 35207 13889 35219 13923
rect 35428 13920 35440 13929
rect 35395 13892 35440 13920
rect 35161 13883 35219 13889
rect 35428 13883 35440 13892
rect 35434 13880 35440 13883
rect 35492 13880 35498 13932
rect 33428 13824 34744 13852
rect 39853 13855 39911 13861
rect 39853 13821 39865 13855
rect 39899 13821 39911 13855
rect 39853 13815 39911 13821
rect 25188 13756 25728 13784
rect 25188 13744 25194 13756
rect 26418 13744 26424 13796
rect 26476 13784 26482 13796
rect 27246 13784 27252 13796
rect 26476 13756 27252 13784
rect 26476 13744 26482 13756
rect 27246 13744 27252 13756
rect 27304 13744 27310 13796
rect 39868 13784 39896 13815
rect 40218 13784 40224 13796
rect 39868 13756 40224 13784
rect 40218 13744 40224 13756
rect 40276 13744 40282 13796
rect 23477 13719 23535 13725
rect 23477 13685 23489 13719
rect 23523 13716 23535 13719
rect 24670 13716 24676 13728
rect 23523 13688 24676 13716
rect 23523 13685 23535 13688
rect 23477 13679 23535 13685
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 27154 13676 27160 13728
rect 27212 13676 27218 13728
rect 28534 13676 28540 13728
rect 28592 13716 28598 13728
rect 28994 13716 29000 13728
rect 28592 13688 29000 13716
rect 28592 13676 28598 13688
rect 28994 13676 29000 13688
rect 29052 13676 29058 13728
rect 1104 13626 43884 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 43884 13626
rect 1104 13552 43884 13574
rect 23385 13515 23443 13521
rect 23385 13481 23397 13515
rect 23431 13481 23443 13515
rect 23385 13475 23443 13481
rect 23400 13444 23428 13475
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 23569 13515 23627 13521
rect 23569 13512 23581 13515
rect 23532 13484 23581 13512
rect 23532 13472 23538 13484
rect 23569 13481 23581 13484
rect 23615 13481 23627 13515
rect 23569 13475 23627 13481
rect 27522 13472 27528 13524
rect 27580 13472 27586 13524
rect 23658 13444 23664 13456
rect 23400 13416 23664 13444
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 32306 13404 32312 13456
rect 32364 13444 32370 13456
rect 38654 13444 38660 13456
rect 32364 13416 38660 13444
rect 32364 13404 32370 13416
rect 38654 13404 38660 13416
rect 38712 13444 38718 13456
rect 38712 13416 38792 13444
rect 38712 13404 38718 13416
rect 25314 13336 25320 13388
rect 25372 13336 25378 13388
rect 33962 13376 33968 13388
rect 32600 13348 33968 13376
rect 23934 13268 23940 13320
rect 23992 13308 23998 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 23992 13280 24593 13308
rect 23992 13268 23998 13280
rect 24581 13277 24593 13280
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 26142 13268 26148 13320
rect 26200 13308 26206 13320
rect 28534 13308 28540 13320
rect 26200 13280 28540 13308
rect 26200 13268 26206 13280
rect 28534 13268 28540 13280
rect 28592 13268 28598 13320
rect 29730 13268 29736 13320
rect 29788 13308 29794 13320
rect 32600 13317 32628 13348
rect 33962 13336 33968 13348
rect 34020 13336 34026 13388
rect 37274 13336 37280 13388
rect 37332 13376 37338 13388
rect 38764 13385 38792 13416
rect 38838 13404 38844 13456
rect 38896 13444 38902 13456
rect 38896 13416 40632 13444
rect 38896 13404 38902 13416
rect 40604 13385 40632 13416
rect 37461 13379 37519 13385
rect 37461 13376 37473 13379
rect 37332 13348 37473 13376
rect 37332 13336 37338 13348
rect 37461 13345 37473 13348
rect 37507 13345 37519 13379
rect 37461 13339 37519 13345
rect 38381 13379 38439 13385
rect 38381 13345 38393 13379
rect 38427 13345 38439 13379
rect 38381 13339 38439 13345
rect 38749 13379 38807 13385
rect 38749 13345 38761 13379
rect 38795 13345 38807 13379
rect 40589 13379 40647 13385
rect 38749 13339 38807 13345
rect 38856 13348 40448 13376
rect 32585 13311 32643 13317
rect 32585 13308 32597 13311
rect 29788 13280 32597 13308
rect 29788 13268 29794 13280
rect 32585 13277 32597 13280
rect 32631 13277 32643 13311
rect 32585 13271 32643 13277
rect 32950 13268 32956 13320
rect 33008 13308 33014 13320
rect 33045 13311 33103 13317
rect 33045 13308 33057 13311
rect 33008 13280 33057 13308
rect 33008 13268 33014 13280
rect 33045 13277 33057 13280
rect 33091 13277 33103 13311
rect 33045 13271 33103 13277
rect 23198 13200 23204 13252
rect 23256 13200 23262 13252
rect 26412 13243 26470 13249
rect 26412 13209 26424 13243
rect 26458 13240 26470 13243
rect 27154 13240 27160 13252
rect 26458 13212 27160 13240
rect 26458 13209 26470 13212
rect 26412 13203 26470 13209
rect 27154 13200 27160 13212
rect 27212 13200 27218 13252
rect 29914 13200 29920 13252
rect 29972 13240 29978 13252
rect 33060 13240 33088 13271
rect 34698 13268 34704 13320
rect 34756 13308 34762 13320
rect 35621 13311 35679 13317
rect 35621 13308 35633 13311
rect 34756 13280 35633 13308
rect 34756 13268 34762 13280
rect 35621 13277 35633 13280
rect 35667 13277 35679 13311
rect 35621 13271 35679 13277
rect 35802 13268 35808 13320
rect 35860 13268 35866 13320
rect 35894 13268 35900 13320
rect 35952 13268 35958 13320
rect 35989 13311 36047 13317
rect 35989 13277 36001 13311
rect 36035 13308 36047 13311
rect 36078 13308 36084 13320
rect 36035 13280 36084 13308
rect 36035 13277 36047 13280
rect 35989 13271 36047 13277
rect 36078 13268 36084 13280
rect 36136 13268 36142 13320
rect 37369 13311 37427 13317
rect 37369 13277 37381 13311
rect 37415 13277 37427 13311
rect 37369 13271 37427 13277
rect 35820 13240 35848 13268
rect 29972 13212 35848 13240
rect 36265 13243 36323 13249
rect 29972 13200 29978 13212
rect 36265 13209 36277 13243
rect 36311 13240 36323 13243
rect 37384 13240 37412 13271
rect 38286 13268 38292 13320
rect 38344 13268 38350 13320
rect 36311 13212 37412 13240
rect 38396 13240 38424 13339
rect 38856 13317 38884 13348
rect 40420 13317 40448 13348
rect 40589 13345 40601 13379
rect 40635 13345 40647 13379
rect 40589 13339 40647 13345
rect 38841 13311 38899 13317
rect 38841 13277 38853 13311
rect 38887 13277 38899 13311
rect 38841 13271 38899 13277
rect 40405 13311 40463 13317
rect 40405 13277 40417 13311
rect 40451 13308 40463 13311
rect 41138 13308 41144 13320
rect 40451 13280 41144 13308
rect 40451 13277 40463 13280
rect 40405 13271 40463 13277
rect 41138 13268 41144 13280
rect 41196 13268 41202 13320
rect 39942 13240 39948 13252
rect 38396 13212 39948 13240
rect 36311 13209 36323 13212
rect 36265 13203 36323 13209
rect 39942 13200 39948 13212
rect 40000 13200 40006 13252
rect 40126 13200 40132 13252
rect 40184 13240 40190 13252
rect 40497 13243 40555 13249
rect 40497 13240 40509 13243
rect 40184 13212 40509 13240
rect 40184 13200 40190 13212
rect 40497 13209 40509 13212
rect 40543 13209 40555 13243
rect 40497 13203 40555 13209
rect 23106 13132 23112 13184
rect 23164 13172 23170 13184
rect 23401 13175 23459 13181
rect 23401 13172 23413 13175
rect 23164 13144 23413 13172
rect 23164 13132 23170 13144
rect 23401 13141 23413 13144
rect 23447 13172 23459 13175
rect 25590 13172 25596 13184
rect 23447 13144 25596 13172
rect 23447 13141 23459 13144
rect 23401 13135 23459 13141
rect 25590 13132 25596 13144
rect 25648 13132 25654 13184
rect 32217 13175 32275 13181
rect 32217 13141 32229 13175
rect 32263 13172 32275 13175
rect 32306 13172 32312 13184
rect 32263 13144 32312 13172
rect 32263 13141 32275 13144
rect 32217 13135 32275 13141
rect 32306 13132 32312 13144
rect 32364 13132 32370 13184
rect 40034 13132 40040 13184
rect 40092 13132 40098 13184
rect 1104 13082 43884 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 43884 13082
rect 1104 13008 43884 13030
rect 23382 12928 23388 12980
rect 23440 12928 23446 12980
rect 29914 12968 29920 12980
rect 24964 12940 29920 12968
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 22272 12835 22330 12841
rect 22272 12801 22284 12835
rect 22318 12832 22330 12835
rect 22646 12832 22652 12844
rect 22318 12804 22652 12832
rect 22318 12801 22330 12804
rect 22272 12795 22330 12801
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 24670 12792 24676 12844
rect 24728 12792 24734 12844
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12832 24823 12835
rect 24854 12832 24860 12844
rect 24811 12804 24860 12832
rect 24811 12801 24823 12804
rect 24765 12795 24823 12801
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 24964 12841 24992 12940
rect 29914 12928 29920 12940
rect 29972 12928 29978 12980
rect 34698 12928 34704 12980
rect 34756 12928 34762 12980
rect 35618 12928 35624 12980
rect 35676 12928 35682 12980
rect 36446 12928 36452 12980
rect 36504 12968 36510 12980
rect 37553 12971 37611 12977
rect 37553 12968 37565 12971
rect 36504 12940 37565 12968
rect 36504 12928 36510 12940
rect 37553 12937 37565 12940
rect 37599 12937 37611 12971
rect 37553 12931 37611 12937
rect 41138 12928 41144 12980
rect 41196 12928 41202 12980
rect 25409 12903 25467 12909
rect 25409 12869 25421 12903
rect 25455 12900 25467 12903
rect 28261 12903 28319 12909
rect 25455 12872 27936 12900
rect 25455 12869 25467 12872
rect 25409 12863 25467 12869
rect 24949 12835 25007 12841
rect 24949 12801 24961 12835
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 26970 12792 26976 12844
rect 27028 12832 27034 12844
rect 27709 12835 27767 12841
rect 27709 12832 27721 12835
rect 27028 12804 27721 12832
rect 27028 12792 27034 12804
rect 27709 12801 27721 12804
rect 27755 12801 27767 12835
rect 27709 12795 27767 12801
rect 27798 12792 27804 12844
rect 27856 12792 27862 12844
rect 27908 12832 27936 12872
rect 28261 12869 28273 12903
rect 28307 12900 28319 12903
rect 29730 12900 29736 12912
rect 28307 12872 29736 12900
rect 28307 12869 28319 12872
rect 28261 12863 28319 12869
rect 29730 12860 29736 12872
rect 29788 12860 29794 12912
rect 31297 12903 31355 12909
rect 31297 12869 31309 12903
rect 31343 12900 31355 12903
rect 31478 12900 31484 12912
rect 31343 12872 31484 12900
rect 31343 12869 31355 12872
rect 31297 12863 31355 12869
rect 31478 12860 31484 12872
rect 31536 12860 31542 12912
rect 33042 12900 33048 12912
rect 32508 12872 33048 12900
rect 29546 12832 29552 12844
rect 27908 12804 29552 12832
rect 29546 12792 29552 12804
rect 29604 12792 29610 12844
rect 30650 12792 30656 12844
rect 30708 12792 30714 12844
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12832 30895 12835
rect 31570 12832 31576 12844
rect 30883 12804 31576 12832
rect 30883 12801 30895 12804
rect 30837 12795 30895 12801
rect 31570 12792 31576 12804
rect 31628 12792 31634 12844
rect 32398 12792 32404 12844
rect 32456 12832 32462 12844
rect 32508 12841 32536 12872
rect 33042 12860 33048 12872
rect 33100 12860 33106 12912
rect 35342 12860 35348 12912
rect 35400 12900 35406 12912
rect 35636 12900 35664 12928
rect 40034 12909 40040 12912
rect 40028 12900 40040 12909
rect 35400 12872 35572 12900
rect 35636 12872 39068 12900
rect 39995 12872 40040 12900
rect 35400 12860 35406 12872
rect 32766 12841 32772 12844
rect 32493 12835 32551 12841
rect 32493 12832 32505 12835
rect 32456 12804 32505 12832
rect 32456 12792 32462 12804
rect 32493 12801 32505 12804
rect 32539 12801 32551 12835
rect 32493 12795 32551 12801
rect 32760 12795 32772 12841
rect 32766 12792 32772 12795
rect 32824 12792 32830 12844
rect 33962 12792 33968 12844
rect 34020 12832 34026 12844
rect 34146 12832 34152 12844
rect 34020 12804 34152 12832
rect 34020 12792 34026 12804
rect 34146 12792 34152 12804
rect 34204 12832 34210 12844
rect 34333 12835 34391 12841
rect 34333 12832 34345 12835
rect 34204 12804 34345 12832
rect 34204 12792 34210 12804
rect 34333 12801 34345 12804
rect 34379 12801 34391 12835
rect 34333 12795 34391 12801
rect 34517 12835 34575 12841
rect 34517 12801 34529 12835
rect 34563 12801 34575 12835
rect 34517 12795 34575 12801
rect 30558 12724 30564 12776
rect 30616 12724 30622 12776
rect 34532 12764 34560 12795
rect 34698 12792 34704 12844
rect 34756 12832 34762 12844
rect 35544 12841 35572 12872
rect 35253 12835 35311 12841
rect 35253 12832 35265 12835
rect 34756 12804 35265 12832
rect 34756 12792 34762 12804
rect 35253 12801 35265 12804
rect 35299 12801 35311 12835
rect 35253 12795 35311 12801
rect 35437 12835 35495 12841
rect 35437 12801 35449 12835
rect 35483 12801 35495 12835
rect 35437 12795 35495 12801
rect 35529 12835 35587 12841
rect 35529 12801 35541 12835
rect 35575 12801 35587 12835
rect 35529 12795 35587 12801
rect 33888 12736 34560 12764
rect 35452 12764 35480 12795
rect 35618 12792 35624 12844
rect 35676 12792 35682 12844
rect 37461 12835 37519 12841
rect 37461 12832 37473 12835
rect 35912 12804 37473 12832
rect 35802 12764 35808 12776
rect 35452 12736 35808 12764
rect 23658 12656 23664 12708
rect 23716 12696 23722 12708
rect 25682 12696 25688 12708
rect 23716 12668 25688 12696
rect 23716 12656 23722 12668
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 33888 12640 33916 12736
rect 35802 12724 35808 12736
rect 35860 12724 35866 12776
rect 35912 12773 35940 12804
rect 37461 12801 37473 12804
rect 37507 12801 37519 12835
rect 37461 12795 37519 12801
rect 38286 12792 38292 12844
rect 38344 12792 38350 12844
rect 38654 12792 38660 12844
rect 38712 12792 38718 12844
rect 38930 12792 38936 12844
rect 38988 12792 38994 12844
rect 39040 12832 39068 12872
rect 40028 12863 40040 12872
rect 40034 12860 40040 12863
rect 40092 12860 40098 12912
rect 42889 12835 42947 12841
rect 42889 12832 42901 12835
rect 39040 12804 42901 12832
rect 42889 12801 42901 12804
rect 42935 12801 42947 12835
rect 42889 12795 42947 12801
rect 35897 12767 35955 12773
rect 35897 12733 35909 12767
rect 35943 12733 35955 12767
rect 35897 12727 35955 12733
rect 38470 12724 38476 12776
rect 38528 12724 38534 12776
rect 39758 12724 39764 12776
rect 39816 12724 39822 12776
rect 43162 12724 43168 12776
rect 43220 12724 43226 12776
rect 25130 12588 25136 12640
rect 25188 12628 25194 12640
rect 30466 12628 30472 12640
rect 25188 12600 30472 12628
rect 25188 12588 25194 12600
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 33870 12588 33876 12640
rect 33928 12588 33934 12640
rect 1104 12538 43884 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 43884 12538
rect 1104 12464 43884 12486
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 26605 12427 26663 12433
rect 26605 12424 26617 12427
rect 24912 12396 26617 12424
rect 24912 12384 24918 12396
rect 26605 12393 26617 12396
rect 26651 12393 26663 12427
rect 26605 12387 26663 12393
rect 29181 12427 29239 12433
rect 29181 12393 29193 12427
rect 29227 12424 29239 12427
rect 30558 12424 30564 12436
rect 29227 12396 30564 12424
rect 29227 12393 29239 12396
rect 29181 12387 29239 12393
rect 30558 12384 30564 12396
rect 30616 12384 30622 12436
rect 30650 12384 30656 12436
rect 30708 12424 30714 12436
rect 30837 12427 30895 12433
rect 30837 12424 30849 12427
rect 30708 12396 30849 12424
rect 30708 12384 30714 12396
rect 30837 12393 30849 12396
rect 30883 12393 30895 12427
rect 30837 12387 30895 12393
rect 32766 12384 32772 12436
rect 32824 12424 32830 12436
rect 32953 12427 33011 12433
rect 32953 12424 32965 12427
rect 32824 12396 32965 12424
rect 32824 12384 32830 12396
rect 32953 12393 32965 12396
rect 32999 12393 33011 12427
rect 32953 12387 33011 12393
rect 39942 12384 39948 12436
rect 40000 12424 40006 12436
rect 41417 12427 41475 12433
rect 41417 12424 41429 12427
rect 40000 12396 41429 12424
rect 40000 12384 40006 12396
rect 41417 12393 41429 12396
rect 41463 12393 41475 12427
rect 41417 12387 41475 12393
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 26418 12356 26424 12368
rect 24820 12328 26424 12356
rect 24820 12316 24826 12328
rect 26418 12316 26424 12328
rect 26476 12356 26482 12368
rect 26476 12328 26740 12356
rect 26476 12316 26482 12328
rect 26712 12297 26740 12328
rect 33318 12316 33324 12368
rect 33376 12356 33382 12368
rect 33376 12328 33548 12356
rect 33376 12316 33382 12328
rect 23293 12291 23351 12297
rect 23293 12257 23305 12291
rect 23339 12288 23351 12291
rect 26053 12291 26111 12297
rect 23339 12260 24900 12288
rect 23339 12257 23351 12260
rect 23293 12251 23351 12257
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12220 23075 12223
rect 23382 12220 23388 12232
rect 23063 12192 23388 12220
rect 23063 12189 23075 12192
rect 23017 12183 23075 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 24762 12180 24768 12232
rect 24820 12180 24826 12232
rect 24872 12152 24900 12260
rect 26053 12257 26065 12291
rect 26099 12288 26111 12291
rect 26513 12291 26571 12297
rect 26513 12288 26525 12291
rect 26099 12260 26525 12288
rect 26099 12257 26111 12260
rect 26053 12251 26111 12257
rect 26513 12257 26525 12260
rect 26559 12257 26571 12291
rect 26513 12251 26571 12257
rect 26697 12291 26755 12297
rect 26697 12257 26709 12291
rect 26743 12288 26755 12291
rect 28629 12291 28687 12297
rect 28629 12288 28641 12291
rect 26743 12260 28641 12288
rect 26743 12257 26755 12260
rect 26697 12251 26755 12257
rect 28629 12257 28641 12260
rect 28675 12288 28687 12291
rect 31294 12288 31300 12300
rect 28675 12260 31300 12288
rect 28675 12257 28687 12260
rect 28629 12251 28687 12257
rect 31294 12248 31300 12260
rect 31352 12288 31358 12300
rect 31389 12291 31447 12297
rect 31389 12288 31401 12291
rect 31352 12260 31401 12288
rect 31352 12248 31358 12260
rect 31389 12257 31401 12260
rect 31435 12257 31447 12291
rect 31389 12251 31447 12257
rect 32582 12248 32588 12300
rect 32640 12288 32646 12300
rect 33520 12297 33548 12328
rect 33413 12291 33471 12297
rect 33413 12288 33425 12291
rect 32640 12260 33425 12288
rect 32640 12248 32646 12260
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25314 12220 25320 12232
rect 25087 12192 25320 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 25314 12180 25320 12192
rect 25372 12180 25378 12232
rect 25590 12180 25596 12232
rect 25648 12180 25654 12232
rect 25682 12180 25688 12232
rect 25740 12180 25746 12232
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 26602 12220 26608 12232
rect 25915 12192 26608 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 26786 12180 26792 12232
rect 26844 12180 26850 12232
rect 28810 12220 28816 12232
rect 28644 12192 28816 12220
rect 28644 12164 28672 12192
rect 28810 12180 28816 12192
rect 28868 12180 28874 12232
rect 28626 12152 28632 12164
rect 24872 12124 28632 12152
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 28721 12155 28779 12161
rect 28721 12121 28733 12155
rect 28767 12152 28779 12155
rect 28902 12152 28908 12164
rect 28767 12124 28908 12152
rect 28767 12121 28779 12124
rect 28721 12115 28779 12121
rect 28902 12112 28908 12124
rect 28960 12112 28966 12164
rect 33244 12152 33272 12260
rect 33413 12257 33425 12260
rect 33459 12257 33471 12291
rect 33413 12251 33471 12257
rect 33505 12291 33563 12297
rect 33505 12257 33517 12291
rect 33551 12257 33563 12291
rect 33505 12251 33563 12257
rect 35710 12248 35716 12300
rect 35768 12288 35774 12300
rect 36081 12291 36139 12297
rect 36081 12288 36093 12291
rect 35768 12260 36093 12288
rect 35768 12248 35774 12260
rect 36081 12257 36093 12260
rect 36127 12257 36139 12291
rect 36081 12251 36139 12257
rect 33321 12223 33379 12229
rect 33321 12189 33333 12223
rect 33367 12220 33379 12223
rect 33870 12220 33876 12232
rect 33367 12192 33876 12220
rect 33367 12189 33379 12192
rect 33321 12183 33379 12189
rect 33870 12180 33876 12192
rect 33928 12180 33934 12232
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 39758 12220 39764 12232
rect 37608 12192 39764 12220
rect 37608 12180 37614 12192
rect 39758 12180 39764 12192
rect 39816 12220 39822 12232
rect 40037 12223 40095 12229
rect 40037 12220 40049 12223
rect 39816 12192 40049 12220
rect 39816 12180 39822 12192
rect 40037 12189 40049 12192
rect 40083 12189 40095 12223
rect 40037 12183 40095 12189
rect 35989 12155 36047 12161
rect 35989 12152 36001 12155
rect 33244 12124 36001 12152
rect 35989 12121 36001 12124
rect 36035 12152 36047 12155
rect 40126 12152 40132 12164
rect 36035 12124 40132 12152
rect 36035 12121 36047 12124
rect 35989 12115 36047 12121
rect 40126 12112 40132 12124
rect 40184 12112 40190 12164
rect 40304 12155 40362 12161
rect 40304 12121 40316 12155
rect 40350 12152 40362 12155
rect 40586 12152 40592 12164
rect 40350 12124 40592 12152
rect 40350 12121 40362 12124
rect 40304 12115 40362 12121
rect 40586 12112 40592 12124
rect 40644 12112 40650 12164
rect 23106 12044 23112 12096
rect 23164 12044 23170 12096
rect 28810 12044 28816 12096
rect 28868 12044 28874 12096
rect 31202 12044 31208 12096
rect 31260 12044 31266 12096
rect 31294 12044 31300 12096
rect 31352 12044 31358 12096
rect 35526 12044 35532 12096
rect 35584 12044 35590 12096
rect 35897 12087 35955 12093
rect 35897 12053 35909 12087
rect 35943 12084 35955 12087
rect 36078 12084 36084 12096
rect 35943 12056 36084 12084
rect 35943 12053 35955 12056
rect 35897 12047 35955 12053
rect 36078 12044 36084 12056
rect 36136 12084 36142 12096
rect 36538 12084 36544 12096
rect 36136 12056 36544 12084
rect 36136 12044 36142 12056
rect 36538 12044 36544 12056
rect 36596 12044 36602 12096
rect 1104 11994 43884 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 43884 11994
rect 1104 11920 43884 11942
rect 23109 11883 23167 11889
rect 23109 11849 23121 11883
rect 23155 11880 23167 11883
rect 23198 11880 23204 11892
rect 23155 11852 23204 11880
rect 23155 11849 23167 11852
rect 23109 11843 23167 11849
rect 23198 11840 23204 11852
rect 23256 11840 23262 11892
rect 24949 11883 25007 11889
rect 24949 11880 24961 11883
rect 24412 11852 24961 11880
rect 23106 11704 23112 11756
rect 23164 11744 23170 11756
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 23164 11716 23213 11744
rect 23164 11704 23170 11716
rect 23201 11713 23213 11716
rect 23247 11744 23259 11747
rect 24412 11744 24440 11852
rect 24949 11849 24961 11852
rect 24995 11880 25007 11883
rect 26329 11883 26387 11889
rect 26329 11880 26341 11883
rect 24995 11852 26341 11880
rect 24995 11849 25007 11852
rect 24949 11843 25007 11849
rect 26329 11849 26341 11852
rect 26375 11880 26387 11883
rect 27890 11880 27896 11892
rect 26375 11852 27896 11880
rect 26375 11849 26387 11852
rect 26329 11843 26387 11849
rect 27890 11840 27896 11852
rect 27948 11840 27954 11892
rect 28445 11883 28503 11889
rect 28445 11849 28457 11883
rect 28491 11880 28503 11883
rect 28810 11880 28816 11892
rect 28491 11852 28816 11880
rect 28491 11849 28503 11852
rect 28445 11843 28503 11849
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 29822 11840 29828 11892
rect 29880 11880 29886 11892
rect 30926 11880 30932 11892
rect 29880 11852 30932 11880
rect 29880 11840 29886 11852
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 34149 11883 34207 11889
rect 34149 11849 34161 11883
rect 34195 11880 34207 11883
rect 34698 11880 34704 11892
rect 34195 11852 34704 11880
rect 34195 11849 34207 11852
rect 34149 11843 34207 11849
rect 34698 11840 34704 11852
rect 34756 11840 34762 11892
rect 36538 11840 36544 11892
rect 36596 11840 36602 11892
rect 36814 11840 36820 11892
rect 36872 11880 36878 11892
rect 36872 11852 39712 11880
rect 36872 11840 36878 11852
rect 24857 11815 24915 11821
rect 24857 11781 24869 11815
rect 24903 11812 24915 11815
rect 26786 11812 26792 11824
rect 24903 11784 26792 11812
rect 24903 11781 24915 11784
rect 24857 11775 24915 11781
rect 26786 11772 26792 11784
rect 26844 11772 26850 11824
rect 28534 11772 28540 11824
rect 28592 11812 28598 11824
rect 29840 11812 29868 11840
rect 28592 11784 29868 11812
rect 33781 11815 33839 11821
rect 28592 11772 28598 11784
rect 33781 11781 33793 11815
rect 33827 11812 33839 11815
rect 34054 11812 34060 11824
rect 33827 11784 34060 11812
rect 33827 11781 33839 11784
rect 33781 11775 33839 11781
rect 34054 11772 34060 11784
rect 34112 11772 34118 11824
rect 35428 11815 35486 11821
rect 35428 11781 35440 11815
rect 35474 11812 35486 11815
rect 35526 11812 35532 11824
rect 35474 11784 35532 11812
rect 35474 11781 35486 11784
rect 35428 11775 35486 11781
rect 35526 11772 35532 11784
rect 35584 11772 35590 11824
rect 38197 11815 38255 11821
rect 38197 11781 38209 11815
rect 38243 11812 38255 11815
rect 38286 11812 38292 11824
rect 38243 11784 38292 11812
rect 38243 11781 38255 11784
rect 38197 11775 38255 11781
rect 38286 11772 38292 11784
rect 38344 11772 38350 11824
rect 23247 11716 24440 11744
rect 26237 11747 26295 11753
rect 23247 11713 23259 11716
rect 23201 11707 23259 11713
rect 26237 11713 26249 11747
rect 26283 11744 26295 11747
rect 26602 11744 26608 11756
rect 26283 11716 26608 11744
rect 26283 11713 26295 11716
rect 26237 11707 26295 11713
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 30837 11747 30895 11753
rect 27356 11716 30788 11744
rect 27356 11688 27384 11716
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 23400 11608 23428 11639
rect 25130 11636 25136 11688
rect 25188 11636 25194 11688
rect 26513 11679 26571 11685
rect 26513 11645 26525 11679
rect 26559 11676 26571 11679
rect 27338 11676 27344 11688
rect 26559 11648 27344 11676
rect 26559 11645 26571 11648
rect 26513 11639 26571 11645
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 28721 11679 28779 11685
rect 28721 11645 28733 11679
rect 28767 11676 28779 11679
rect 30282 11676 30288 11688
rect 28767 11648 30288 11676
rect 28767 11645 28779 11648
rect 28721 11639 28779 11645
rect 28736 11608 28764 11639
rect 30282 11636 30288 11648
rect 30340 11636 30346 11688
rect 30760 11676 30788 11716
rect 30837 11713 30849 11747
rect 30883 11744 30895 11747
rect 31294 11744 31300 11756
rect 30883 11716 31300 11744
rect 30883 11713 30895 11716
rect 30837 11707 30895 11713
rect 31294 11704 31300 11716
rect 31352 11704 31358 11756
rect 33962 11704 33968 11756
rect 34020 11704 34026 11756
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 35161 11747 35219 11753
rect 35161 11744 35173 11747
rect 34848 11716 35173 11744
rect 34848 11704 34854 11716
rect 35161 11713 35173 11716
rect 35207 11713 35219 11747
rect 35161 11707 35219 11713
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11744 38163 11747
rect 38470 11744 38476 11756
rect 38151 11716 38476 11744
rect 38151 11713 38163 11716
rect 38105 11707 38163 11713
rect 38470 11704 38476 11716
rect 38528 11704 38534 11756
rect 39684 11744 39712 11852
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 40221 11883 40279 11889
rect 40221 11880 40233 11883
rect 40000 11852 40233 11880
rect 40000 11840 40006 11852
rect 40221 11849 40233 11852
rect 40267 11849 40279 11883
rect 40221 11843 40279 11849
rect 40586 11840 40592 11892
rect 40644 11840 40650 11892
rect 40126 11772 40132 11824
rect 40184 11772 40190 11824
rect 42889 11747 42947 11753
rect 42889 11744 42901 11747
rect 39684 11716 42901 11744
rect 42889 11713 42901 11716
rect 42935 11713 42947 11747
rect 42889 11707 42947 11713
rect 31021 11679 31079 11685
rect 31021 11676 31033 11679
rect 30760 11648 31033 11676
rect 31021 11645 31033 11648
rect 31067 11645 31079 11679
rect 31021 11639 31079 11645
rect 38378 11636 38384 11688
rect 38436 11676 38442 11688
rect 39945 11679 40003 11685
rect 39945 11676 39957 11679
rect 38436 11648 39957 11676
rect 38436 11636 38442 11648
rect 39945 11645 39957 11648
rect 39991 11676 40003 11679
rect 40218 11676 40224 11688
rect 39991 11648 40224 11676
rect 39991 11645 40003 11648
rect 39945 11639 40003 11645
rect 40218 11636 40224 11648
rect 40276 11636 40282 11688
rect 43162 11636 43168 11688
rect 43220 11636 43226 11688
rect 23400 11580 28764 11608
rect 22738 11500 22744 11552
rect 22796 11500 22802 11552
rect 24489 11543 24547 11549
rect 24489 11509 24501 11543
rect 24535 11540 24547 11543
rect 24670 11540 24676 11552
rect 24535 11512 24676 11540
rect 24535 11509 24547 11512
rect 24489 11503 24547 11509
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 25866 11500 25872 11552
rect 25924 11500 25930 11552
rect 28074 11500 28080 11552
rect 28132 11500 28138 11552
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30469 11543 30527 11549
rect 30469 11540 30481 11543
rect 30432 11512 30481 11540
rect 30432 11500 30438 11512
rect 30469 11509 30481 11512
rect 30515 11509 30527 11543
rect 30469 11503 30527 11509
rect 37737 11543 37795 11549
rect 37737 11509 37749 11543
rect 37783 11540 37795 11543
rect 37826 11540 37832 11552
rect 37783 11512 37832 11540
rect 37783 11509 37795 11512
rect 37737 11503 37795 11509
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 1104 11450 43884 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 43884 11450
rect 1104 11376 43884 11398
rect 23198 11296 23204 11348
rect 23256 11296 23262 11348
rect 25961 11339 26019 11345
rect 25961 11305 25973 11339
rect 26007 11336 26019 11339
rect 26786 11336 26792 11348
rect 26007 11308 26792 11336
rect 26007 11305 26019 11308
rect 25961 11299 26019 11305
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 28721 11339 28779 11345
rect 28721 11305 28733 11339
rect 28767 11336 28779 11339
rect 28810 11336 28816 11348
rect 28767 11308 28816 11336
rect 28767 11305 28779 11308
rect 28721 11299 28779 11305
rect 28810 11296 28816 11308
rect 28868 11296 28874 11348
rect 31294 11296 31300 11348
rect 31352 11336 31358 11348
rect 31481 11339 31539 11345
rect 31481 11336 31493 11339
rect 31352 11308 31493 11336
rect 31352 11296 31358 11308
rect 31481 11305 31493 11308
rect 31527 11305 31539 11339
rect 31481 11299 31539 11305
rect 33781 11339 33839 11345
rect 33781 11305 33793 11339
rect 33827 11336 33839 11339
rect 33962 11336 33968 11348
rect 33827 11308 33968 11336
rect 33827 11305 33839 11308
rect 33781 11299 33839 11305
rect 33962 11296 33968 11308
rect 34020 11296 34026 11348
rect 35618 11296 35624 11348
rect 35676 11336 35682 11348
rect 36265 11339 36323 11345
rect 36265 11336 36277 11339
rect 35676 11308 36277 11336
rect 35676 11296 35682 11308
rect 36265 11305 36277 11308
rect 36311 11305 36323 11339
rect 36265 11299 36323 11305
rect 38470 11296 38476 11348
rect 38528 11336 38534 11348
rect 38933 11339 38991 11345
rect 38933 11336 38945 11339
rect 38528 11308 38945 11336
rect 38528 11296 38534 11308
rect 38933 11305 38945 11308
rect 38979 11305 38991 11339
rect 38933 11299 38991 11305
rect 26142 11160 26148 11212
rect 26200 11200 26206 11212
rect 27341 11203 27399 11209
rect 27341 11200 27353 11203
rect 26200 11172 27353 11200
rect 26200 11160 26206 11172
rect 27341 11169 27353 11172
rect 27387 11169 27399 11203
rect 27341 11163 27399 11169
rect 28994 11160 29000 11212
rect 29052 11200 29058 11212
rect 30098 11200 30104 11212
rect 29052 11172 30104 11200
rect 29052 11160 29058 11172
rect 30098 11160 30104 11172
rect 30156 11160 30162 11212
rect 32398 11160 32404 11212
rect 32456 11160 32462 11212
rect 34790 11160 34796 11212
rect 34848 11200 34854 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34848 11172 34897 11200
rect 34848 11160 34854 11172
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 34885 11163 34943 11169
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11132 21879 11135
rect 21910 11132 21916 11144
rect 21867 11104 21916 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 21910 11092 21916 11104
rect 21968 11132 21974 11144
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 21968 11104 24593 11132
rect 21968 11092 21974 11104
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24670 11092 24676 11144
rect 24728 11132 24734 11144
rect 24837 11135 24895 11141
rect 24837 11132 24849 11135
rect 24728 11104 24849 11132
rect 24728 11092 24734 11104
rect 24837 11101 24849 11104
rect 24883 11101 24895 11135
rect 24837 11095 24895 11101
rect 27608 11135 27666 11141
rect 27608 11101 27620 11135
rect 27654 11132 27666 11135
rect 28074 11132 28080 11144
rect 27654 11104 28080 11132
rect 27654 11101 27666 11104
rect 27608 11095 27666 11101
rect 28074 11092 28080 11104
rect 28132 11092 28138 11144
rect 30374 11141 30380 11144
rect 30368 11132 30380 11141
rect 30335 11104 30380 11132
rect 30368 11095 30380 11104
rect 30374 11092 30380 11095
rect 30432 11092 30438 11144
rect 34900 11132 34928 11163
rect 37550 11132 37556 11144
rect 34900 11104 37556 11132
rect 37550 11092 37556 11104
rect 37608 11092 37614 11144
rect 37826 11141 37832 11144
rect 37820 11132 37832 11141
rect 37787 11104 37832 11132
rect 37820 11095 37832 11104
rect 37826 11092 37832 11095
rect 37884 11092 37890 11144
rect 22088 11067 22146 11073
rect 22088 11033 22100 11067
rect 22134 11064 22146 11067
rect 22738 11064 22744 11076
rect 22134 11036 22744 11064
rect 22134 11033 22146 11036
rect 22088 11027 22146 11033
rect 22738 11024 22744 11036
rect 22796 11024 22802 11076
rect 32668 11067 32726 11073
rect 32668 11033 32680 11067
rect 32714 11064 32726 11067
rect 32858 11064 32864 11076
rect 32714 11036 32864 11064
rect 32714 11033 32726 11036
rect 32668 11027 32726 11033
rect 32858 11024 32864 11036
rect 32916 11024 32922 11076
rect 35158 11073 35164 11076
rect 35152 11027 35164 11073
rect 35158 11024 35164 11027
rect 35216 11024 35222 11076
rect 1104 10906 43884 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 43884 10906
rect 1104 10832 43884 10854
rect 26602 10752 26608 10804
rect 26660 10752 26666 10804
rect 28902 10752 28908 10804
rect 28960 10792 28966 10804
rect 28997 10795 29055 10801
rect 28997 10792 29009 10795
rect 28960 10764 29009 10792
rect 28960 10752 28966 10764
rect 28997 10761 29009 10764
rect 29043 10761 29055 10795
rect 28997 10755 29055 10761
rect 31202 10752 31208 10804
rect 31260 10792 31266 10804
rect 31481 10795 31539 10801
rect 31481 10792 31493 10795
rect 31260 10764 31493 10792
rect 31260 10752 31266 10764
rect 31481 10761 31493 10764
rect 31527 10761 31539 10795
rect 31481 10755 31539 10761
rect 32858 10752 32864 10804
rect 32916 10752 32922 10804
rect 33229 10795 33287 10801
rect 33229 10761 33241 10795
rect 33275 10792 33287 10795
rect 33962 10792 33968 10804
rect 33275 10764 33968 10792
rect 33275 10761 33287 10764
rect 33229 10755 33287 10761
rect 33962 10752 33968 10764
rect 34020 10752 34026 10804
rect 35069 10795 35127 10801
rect 35069 10761 35081 10795
rect 35115 10792 35127 10795
rect 35158 10792 35164 10804
rect 35115 10764 35164 10792
rect 35115 10761 35127 10764
rect 35069 10755 35127 10761
rect 35158 10752 35164 10764
rect 35216 10752 35222 10804
rect 35437 10795 35495 10801
rect 35437 10761 35449 10795
rect 35483 10792 35495 10795
rect 35618 10792 35624 10804
rect 35483 10764 35624 10792
rect 35483 10761 35495 10764
rect 35437 10755 35495 10761
rect 35618 10752 35624 10764
rect 35676 10752 35682 10804
rect 38930 10752 38936 10804
rect 38988 10752 38994 10804
rect 26142 10724 26148 10736
rect 25240 10696 26148 10724
rect 25240 10665 25268 10696
rect 26142 10684 26148 10696
rect 26200 10684 26206 10736
rect 28718 10724 28724 10736
rect 27632 10696 28724 10724
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 25492 10659 25550 10665
rect 25492 10625 25504 10659
rect 25538 10656 25550 10659
rect 25866 10656 25872 10668
rect 25538 10628 25872 10656
rect 25538 10625 25550 10628
rect 25492 10619 25550 10625
rect 25866 10616 25872 10628
rect 25924 10616 25930 10668
rect 27632 10665 27660 10696
rect 28718 10684 28724 10696
rect 28776 10684 28782 10736
rect 31018 10684 31024 10736
rect 31076 10724 31082 10736
rect 33321 10727 33379 10733
rect 33321 10724 33333 10727
rect 31076 10696 33333 10724
rect 31076 10684 31082 10696
rect 33321 10693 33333 10696
rect 33367 10724 33379 10727
rect 35529 10727 35587 10733
rect 35529 10724 35541 10727
rect 33367 10696 35541 10724
rect 33367 10693 33379 10696
rect 33321 10687 33379 10693
rect 35529 10693 35541 10696
rect 35575 10724 35587 10727
rect 38286 10724 38292 10736
rect 35575 10696 38292 10724
rect 35575 10693 35587 10696
rect 35529 10687 35587 10693
rect 38286 10684 38292 10696
rect 38344 10684 38350 10736
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 27884 10659 27942 10665
rect 27884 10625 27896 10659
rect 27930 10656 27942 10659
rect 28258 10656 28264 10668
rect 27930 10628 28264 10656
rect 27930 10625 27942 10628
rect 27884 10619 27942 10625
rect 28258 10616 28264 10628
rect 28316 10616 28322 10668
rect 30098 10616 30104 10668
rect 30156 10616 30162 10668
rect 30374 10665 30380 10668
rect 30368 10619 30380 10665
rect 30374 10616 30380 10619
rect 30432 10616 30438 10668
rect 37550 10616 37556 10668
rect 37608 10616 37614 10668
rect 37826 10665 37832 10668
rect 37820 10619 37832 10665
rect 37826 10616 37832 10619
rect 37884 10616 37890 10668
rect 33318 10548 33324 10600
rect 33376 10588 33382 10600
rect 33413 10591 33471 10597
rect 33413 10588 33425 10591
rect 33376 10560 33425 10588
rect 33376 10548 33382 10560
rect 33413 10557 33425 10560
rect 33459 10557 33471 10591
rect 33413 10551 33471 10557
rect 35618 10548 35624 10600
rect 35676 10548 35682 10600
rect 1104 10362 43884 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 43884 10362
rect 1104 10288 43884 10310
rect 28258 10208 28264 10260
rect 28316 10208 28322 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 30469 10251 30527 10257
rect 30469 10248 30481 10251
rect 30432 10220 30481 10248
rect 30432 10208 30438 10220
rect 30469 10217 30481 10220
rect 30515 10217 30527 10251
rect 30469 10211 30527 10217
rect 37826 10208 37832 10260
rect 37884 10208 37890 10260
rect 28626 10140 28632 10192
rect 28684 10180 28690 10192
rect 28684 10152 28856 10180
rect 28684 10140 28690 10152
rect 28534 10072 28540 10124
rect 28592 10112 28598 10124
rect 28828 10121 28856 10152
rect 30558 10140 30564 10192
rect 30616 10180 30622 10192
rect 35618 10180 35624 10192
rect 30616 10152 35624 10180
rect 30616 10140 30622 10152
rect 28721 10115 28779 10121
rect 28721 10112 28733 10115
rect 28592 10084 28733 10112
rect 28592 10072 28598 10084
rect 28721 10081 28733 10084
rect 28767 10081 28779 10115
rect 28721 10075 28779 10081
rect 28813 10115 28871 10121
rect 28813 10081 28825 10115
rect 28859 10081 28871 10115
rect 28813 10075 28871 10081
rect 30926 10072 30932 10124
rect 30984 10072 30990 10124
rect 31036 10121 31064 10152
rect 35618 10140 35624 10152
rect 35676 10140 35682 10192
rect 36906 10140 36912 10192
rect 36964 10180 36970 10192
rect 36964 10152 42932 10180
rect 36964 10140 36970 10152
rect 31021 10115 31079 10121
rect 31021 10081 31033 10115
rect 31067 10081 31079 10115
rect 31021 10075 31079 10081
rect 38286 10072 38292 10124
rect 38344 10072 38350 10124
rect 38473 10115 38531 10121
rect 38473 10081 38485 10115
rect 38519 10112 38531 10115
rect 38838 10112 38844 10124
rect 38519 10084 38844 10112
rect 38519 10081 38531 10084
rect 38473 10075 38531 10081
rect 38838 10072 38844 10084
rect 38896 10072 38902 10124
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10044 28687 10047
rect 28902 10044 28908 10056
rect 28675 10016 28908 10044
rect 28675 10013 28687 10016
rect 28629 10007 28687 10013
rect 28902 10004 28908 10016
rect 28960 10004 28966 10056
rect 30837 10047 30895 10053
rect 30837 10013 30849 10047
rect 30883 10044 30895 10047
rect 31202 10044 31208 10056
rect 30883 10016 31208 10044
rect 30883 10013 30895 10016
rect 30837 10007 30895 10013
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 38197 10047 38255 10053
rect 38197 10013 38209 10047
rect 38243 10044 38255 10047
rect 38930 10044 38936 10056
rect 38243 10016 38936 10044
rect 38243 10013 38255 10016
rect 38197 10007 38255 10013
rect 38930 10004 38936 10016
rect 38988 10004 38994 10056
rect 42904 10053 42932 10152
rect 42889 10047 42947 10053
rect 42889 10013 42901 10047
rect 42935 10013 42947 10047
rect 42889 10007 42947 10013
rect 43162 9936 43168 9988
rect 43220 9936 43226 9988
rect 1104 9818 43884 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 43884 9818
rect 1104 9744 43884 9766
rect 1104 9274 43884 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 43884 9274
rect 1104 9200 43884 9222
rect 1104 8730 43884 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 43884 8730
rect 1104 8656 43884 8678
rect 33778 8440 33784 8492
rect 33836 8480 33842 8492
rect 42889 8483 42947 8489
rect 42889 8480 42901 8483
rect 33836 8452 42901 8480
rect 33836 8440 33842 8452
rect 42889 8449 42901 8452
rect 42935 8449 42947 8483
rect 42889 8443 42947 8449
rect 43165 8415 43223 8421
rect 43165 8381 43177 8415
rect 43211 8412 43223 8415
rect 43990 8412 43996 8424
rect 43211 8384 43996 8412
rect 43211 8381 43223 8384
rect 43165 8375 43223 8381
rect 43990 8372 43996 8384
rect 44048 8372 44054 8424
rect 1104 8186 43884 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 43884 8186
rect 1104 8112 43884 8134
rect 1104 7642 43884 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 43884 7642
rect 1104 7568 43884 7590
rect 1104 7098 43884 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 43884 7098
rect 1104 7024 43884 7046
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 42889 6783 42947 6789
rect 42889 6780 42901 6783
rect 33744 6752 42901 6780
rect 33744 6740 33750 6752
rect 42889 6749 42901 6752
rect 42935 6749 42947 6783
rect 42889 6743 42947 6749
rect 43162 6672 43168 6724
rect 43220 6672 43226 6724
rect 1104 6554 43884 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 43884 6554
rect 1104 6480 43884 6502
rect 1104 6010 43884 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 43884 6010
rect 1104 5936 43884 5958
rect 42794 5652 42800 5704
rect 42852 5692 42858 5704
rect 42889 5695 42947 5701
rect 42889 5692 42901 5695
rect 42852 5664 42901 5692
rect 42852 5652 42858 5664
rect 42889 5661 42901 5664
rect 42935 5661 42947 5695
rect 42889 5655 42947 5661
rect 43165 5627 43223 5633
rect 43165 5593 43177 5627
rect 43211 5624 43223 5627
rect 43990 5624 43996 5636
rect 43211 5596 43996 5624
rect 43211 5593 43223 5596
rect 43165 5587 43223 5593
rect 43990 5584 43996 5596
rect 44048 5584 44054 5636
rect 1104 5466 43884 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 43884 5466
rect 1104 5392 43884 5414
rect 1104 4922 43884 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 43884 4922
rect 1104 4848 43884 4870
rect 1104 4378 43884 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 43884 4378
rect 1104 4304 43884 4326
rect 36998 4088 37004 4140
rect 37056 4128 37062 4140
rect 42889 4131 42947 4137
rect 42889 4128 42901 4131
rect 37056 4100 42901 4128
rect 37056 4088 37062 4100
rect 42889 4097 42901 4100
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 43162 4020 43168 4072
rect 43220 4020 43226 4072
rect 1104 3834 43884 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 43884 3834
rect 1104 3760 43884 3782
rect 1104 3290 43884 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 43884 3290
rect 1104 3216 43884 3238
rect 1104 2746 43884 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 43884 2746
rect 1104 2672 43884 2694
rect 34698 2388 34704 2440
rect 34756 2428 34762 2440
rect 42889 2431 42947 2437
rect 42889 2428 42901 2431
rect 34756 2400 42901 2428
rect 34756 2388 34762 2400
rect 42889 2397 42901 2400
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43162 2320 43168 2372
rect 43220 2320 43226 2372
rect 1104 2202 43884 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 43884 2202
rect 1104 2128 43884 2150
<< via1 >>
rect 16948 44072 17000 44124
rect 18144 44072 18196 44124
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 23388 42304 23440 42356
rect 7196 42236 7248 42288
rect 14372 42236 14424 42288
rect 28356 42236 28408 42288
rect 2228 42168 2280 42220
rect 5908 42211 5960 42220
rect 5908 42177 5917 42211
rect 5917 42177 5951 42211
rect 5951 42177 5960 42211
rect 5908 42168 5960 42177
rect 9680 42168 9732 42220
rect 13268 42168 13320 42220
rect 13728 42168 13780 42220
rect 14556 42168 14608 42220
rect 15108 42168 15160 42220
rect 17224 42211 17276 42220
rect 17224 42177 17233 42211
rect 17233 42177 17267 42211
rect 17267 42177 17276 42211
rect 17224 42168 17276 42177
rect 5632 42143 5684 42152
rect 5632 42109 5641 42143
rect 5641 42109 5675 42143
rect 5675 42109 5684 42143
rect 5632 42100 5684 42109
rect 7012 42143 7064 42152
rect 7012 42109 7021 42143
rect 7021 42109 7055 42143
rect 7055 42109 7064 42143
rect 7012 42100 7064 42109
rect 9220 42100 9272 42152
rect 10324 42143 10376 42152
rect 10324 42109 10333 42143
rect 10333 42109 10367 42143
rect 10367 42109 10376 42143
rect 10324 42100 10376 42109
rect 13636 42143 13688 42152
rect 13636 42109 13645 42143
rect 13645 42109 13679 42143
rect 13679 42109 13688 42143
rect 13636 42100 13688 42109
rect 14556 42032 14608 42084
rect 17316 42143 17368 42152
rect 17316 42109 17325 42143
rect 17325 42109 17359 42143
rect 17359 42109 17368 42143
rect 17316 42100 17368 42109
rect 17776 42100 17828 42152
rect 18144 42211 18196 42220
rect 18144 42177 18153 42211
rect 18153 42177 18187 42211
rect 18187 42177 18196 42211
rect 18144 42168 18196 42177
rect 20720 42168 20772 42220
rect 24308 42168 24360 42220
rect 27252 42211 27304 42220
rect 27252 42177 27261 42211
rect 27261 42177 27295 42211
rect 27295 42177 27304 42211
rect 27252 42168 27304 42177
rect 27988 42168 28040 42220
rect 30564 42211 30616 42220
rect 30564 42177 30573 42211
rect 30573 42177 30607 42211
rect 30607 42177 30616 42211
rect 30564 42168 30616 42177
rect 31760 42236 31812 42288
rect 35348 42236 35400 42288
rect 43996 42236 44048 42288
rect 34152 42168 34204 42220
rect 18696 42143 18748 42152
rect 18696 42109 18705 42143
rect 18705 42109 18739 42143
rect 18739 42109 18748 42143
rect 18696 42100 18748 42109
rect 24952 42143 25004 42152
rect 24952 42109 24961 42143
rect 24961 42109 24995 42143
rect 24995 42109 25004 42143
rect 24952 42100 25004 42109
rect 30012 42032 30064 42084
rect 31576 42032 31628 42084
rect 32588 42075 32640 42084
rect 32588 42041 32597 42075
rect 32597 42041 32631 42075
rect 32631 42041 32640 42075
rect 32588 42032 32640 42041
rect 41604 42211 41656 42220
rect 41604 42177 41613 42211
rect 41613 42177 41647 42211
rect 41647 42177 41656 42211
rect 41604 42168 41656 42177
rect 42708 42211 42760 42220
rect 42708 42177 42717 42211
rect 42717 42177 42751 42211
rect 42751 42177 42760 42211
rect 42708 42168 42760 42177
rect 6552 42007 6604 42016
rect 6552 41973 6561 42007
rect 6561 41973 6595 42007
rect 6595 41973 6604 42007
rect 6552 41964 6604 41973
rect 12992 42007 13044 42016
rect 12992 41973 13001 42007
rect 13001 41973 13035 42007
rect 13035 41973 13044 42007
rect 12992 41964 13044 41973
rect 14280 42007 14332 42016
rect 14280 41973 14289 42007
rect 14289 41973 14323 42007
rect 14323 41973 14332 42007
rect 14280 41964 14332 41973
rect 16580 41964 16632 42016
rect 27528 42007 27580 42016
rect 27528 41973 27537 42007
rect 27537 41973 27571 42007
rect 27571 41973 27580 42007
rect 27528 41964 27580 41973
rect 31668 42007 31720 42016
rect 31668 41973 31677 42007
rect 31677 41973 31711 42007
rect 31711 41973 31720 42007
rect 31668 41964 31720 41973
rect 35624 42007 35676 42016
rect 35624 41973 35633 42007
rect 35633 41973 35667 42007
rect 35667 41973 35676 42007
rect 35624 41964 35676 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 7012 41760 7064 41812
rect 27252 41760 27304 41812
rect 5540 41599 5592 41608
rect 5540 41565 5549 41599
rect 5549 41565 5583 41599
rect 5583 41565 5592 41599
rect 5540 41556 5592 41565
rect 6552 41556 6604 41608
rect 9128 41599 9180 41608
rect 9128 41565 9137 41599
rect 9137 41565 9171 41599
rect 9171 41565 9180 41599
rect 9128 41556 9180 41565
rect 12072 41556 12124 41608
rect 12992 41556 13044 41608
rect 16580 41556 16632 41608
rect 17132 41599 17184 41608
rect 17132 41565 17141 41599
rect 17141 41565 17175 41599
rect 17175 41565 17184 41599
rect 17132 41556 17184 41565
rect 20260 41556 20312 41608
rect 21088 41556 21140 41608
rect 27344 41624 27396 41676
rect 27528 41624 27580 41676
rect 30472 41624 30524 41676
rect 34612 41624 34664 41676
rect 22836 41556 22888 41608
rect 23388 41556 23440 41608
rect 9588 41488 9640 41540
rect 17408 41531 17460 41540
rect 17408 41497 17417 41531
rect 17417 41497 17451 41531
rect 17451 41497 17460 41531
rect 17408 41488 17460 41497
rect 21180 41488 21232 41540
rect 22284 41488 22336 41540
rect 24032 41488 24084 41540
rect 10048 41420 10100 41472
rect 13728 41463 13780 41472
rect 13728 41429 13737 41463
rect 13737 41429 13771 41463
rect 13771 41429 13780 41463
rect 13728 41420 13780 41429
rect 17316 41420 17368 41472
rect 17592 41420 17644 41472
rect 22560 41420 22612 41472
rect 23848 41420 23900 41472
rect 26976 41488 27028 41540
rect 28540 41556 28592 41608
rect 28908 41556 28960 41608
rect 29920 41488 29972 41540
rect 31668 41488 31720 41540
rect 27896 41420 27948 41472
rect 30840 41420 30892 41472
rect 31116 41420 31168 41472
rect 33968 41599 34020 41608
rect 33968 41565 34007 41599
rect 34007 41565 34020 41599
rect 33968 41556 34020 41565
rect 34244 41556 34296 41608
rect 41604 41624 41656 41676
rect 35532 41556 35584 41608
rect 41880 41556 41932 41608
rect 32496 41488 32548 41540
rect 35348 41488 35400 41540
rect 38016 41488 38068 41540
rect 40132 41488 40184 41540
rect 43996 41488 44048 41540
rect 33876 41420 33928 41472
rect 35900 41420 35952 41472
rect 39304 41463 39356 41472
rect 39304 41429 39313 41463
rect 39313 41429 39347 41463
rect 39347 41429 39356 41463
rect 39304 41420 39356 41429
rect 41420 41463 41472 41472
rect 41420 41429 41429 41463
rect 41429 41429 41463 41463
rect 41463 41429 41472 41463
rect 41420 41420 41472 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 6828 41216 6880 41268
rect 5540 41148 5592 41200
rect 9128 41148 9180 41200
rect 9588 41259 9640 41268
rect 9588 41225 9597 41259
rect 9597 41225 9631 41259
rect 9631 41225 9640 41259
rect 9588 41216 9640 41225
rect 12164 41259 12216 41268
rect 12164 41225 12173 41259
rect 12173 41225 12207 41259
rect 12207 41225 12216 41259
rect 12164 41216 12216 41225
rect 14280 41148 14332 41200
rect 14556 41148 14608 41200
rect 8392 41080 8444 41132
rect 10324 41080 10376 41132
rect 11980 41080 12032 41132
rect 10048 41055 10100 41064
rect 10048 41021 10057 41055
rect 10057 41021 10091 41055
rect 10091 41021 10100 41055
rect 10048 41012 10100 41021
rect 9220 40944 9272 40996
rect 13636 41012 13688 41064
rect 12072 40944 12124 40996
rect 15016 40944 15068 40996
rect 15844 41123 15896 41132
rect 15844 41089 15853 41123
rect 15853 41089 15887 41123
rect 15887 41089 15896 41123
rect 15844 41080 15896 41089
rect 17224 41191 17276 41200
rect 17224 41157 17233 41191
rect 17233 41157 17267 41191
rect 17267 41157 17276 41191
rect 17224 41148 17276 41157
rect 17592 41216 17644 41268
rect 19984 41148 20036 41200
rect 20352 41148 20404 41200
rect 22284 41216 22336 41268
rect 24400 41216 24452 41268
rect 17960 41080 18012 41132
rect 18052 41123 18104 41132
rect 18052 41089 18061 41123
rect 18061 41089 18095 41123
rect 18095 41089 18104 41123
rect 18052 41080 18104 41089
rect 22284 41123 22336 41132
rect 22284 41089 22293 41123
rect 22293 41089 22327 41123
rect 22327 41089 22336 41123
rect 22284 41080 22336 41089
rect 22836 41080 22888 41132
rect 16488 41012 16540 41064
rect 18420 41012 18472 41064
rect 23848 41080 23900 41132
rect 24124 41123 24176 41132
rect 24124 41089 24133 41123
rect 24133 41089 24167 41123
rect 24167 41089 24176 41123
rect 24124 41080 24176 41089
rect 25228 41123 25280 41132
rect 25228 41089 25237 41123
rect 25237 41089 25271 41123
rect 25271 41089 25280 41123
rect 25228 41080 25280 41089
rect 25964 41080 26016 41132
rect 9036 40919 9088 40928
rect 9036 40885 9045 40919
rect 9045 40885 9079 40919
rect 9079 40885 9088 40919
rect 9036 40876 9088 40885
rect 11704 40919 11756 40928
rect 11704 40885 11713 40919
rect 11713 40885 11747 40919
rect 11747 40885 11756 40919
rect 11704 40876 11756 40885
rect 14648 40876 14700 40928
rect 15108 40876 15160 40928
rect 17132 40944 17184 40996
rect 24676 41055 24728 41064
rect 24676 41021 24685 41055
rect 24685 41021 24719 41055
rect 24719 41021 24728 41055
rect 26240 41055 26292 41064
rect 24676 41012 24728 41021
rect 26240 41021 26249 41055
rect 26249 41021 26283 41055
rect 26283 41021 26292 41055
rect 26240 41012 26292 41021
rect 27252 41123 27304 41132
rect 27252 41089 27261 41123
rect 27261 41089 27295 41123
rect 27295 41089 27304 41123
rect 27252 41080 27304 41089
rect 28632 41216 28684 41268
rect 28816 41216 28868 41268
rect 29000 41216 29052 41268
rect 29092 41216 29144 41268
rect 28908 41148 28960 41200
rect 30840 41216 30892 41268
rect 28080 41012 28132 41064
rect 28448 41012 28500 41064
rect 30104 41080 30156 41132
rect 30196 41080 30248 41132
rect 31024 41080 31076 41132
rect 31116 41123 31168 41132
rect 31116 41089 31125 41123
rect 31125 41089 31159 41123
rect 31159 41089 31168 41123
rect 31116 41080 31168 41089
rect 18696 40876 18748 40928
rect 28540 40944 28592 40996
rect 21088 40876 21140 40928
rect 23480 40919 23532 40928
rect 23480 40885 23489 40919
rect 23489 40885 23523 40919
rect 23523 40885 23532 40919
rect 23480 40876 23532 40885
rect 23848 40876 23900 40928
rect 24952 40876 25004 40928
rect 27068 40876 27120 40928
rect 28448 40876 28500 40928
rect 28816 41012 28868 41064
rect 31668 41123 31720 41132
rect 31668 41089 31677 41123
rect 31677 41089 31711 41123
rect 31711 41089 31720 41123
rect 31668 41080 31720 41089
rect 32496 41123 32548 41132
rect 32496 41089 32502 41123
rect 32502 41089 32548 41123
rect 32496 41080 32548 41089
rect 28724 40944 28776 40996
rect 32036 41012 32088 41064
rect 38016 41259 38068 41268
rect 38016 41225 38025 41259
rect 38025 41225 38059 41259
rect 38059 41225 38068 41259
rect 38016 41216 38068 41225
rect 40132 41216 40184 41268
rect 34244 41148 34296 41200
rect 35624 41148 35676 41200
rect 38384 41148 38436 41200
rect 33692 41123 33744 41132
rect 33692 41089 33701 41123
rect 33701 41089 33735 41123
rect 33735 41089 33744 41123
rect 33692 41080 33744 41089
rect 33968 41080 34020 41132
rect 35532 41123 35584 41132
rect 35532 41089 35541 41123
rect 35541 41089 35575 41123
rect 35575 41089 35584 41123
rect 35532 41080 35584 41089
rect 38568 41080 38620 41132
rect 40684 41080 40736 41132
rect 43076 41080 43128 41132
rect 35440 41012 35492 41064
rect 37556 41055 37608 41064
rect 37556 41021 37565 41055
rect 37565 41021 37599 41055
rect 37599 41021 37608 41055
rect 37556 41012 37608 41021
rect 38476 41012 38528 41064
rect 40040 41012 40092 41064
rect 43996 41012 44048 41064
rect 29920 40987 29972 40996
rect 29920 40953 29929 40987
rect 29929 40953 29963 40987
rect 29963 40953 29972 40987
rect 29920 40944 29972 40953
rect 32588 40987 32640 40996
rect 32588 40953 32597 40987
rect 32597 40953 32631 40987
rect 32631 40953 32640 40987
rect 32588 40944 32640 40953
rect 34244 40944 34296 40996
rect 28816 40876 28868 40928
rect 30104 40876 30156 40928
rect 31852 40876 31904 40928
rect 33508 40919 33560 40928
rect 33508 40885 33517 40919
rect 33517 40885 33551 40919
rect 33551 40885 33560 40919
rect 33508 40876 33560 40885
rect 36912 40919 36964 40928
rect 36912 40885 36921 40919
rect 36921 40885 36955 40919
rect 36955 40885 36964 40919
rect 36912 40876 36964 40885
rect 41512 40876 41564 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 12164 40672 12216 40724
rect 15200 40672 15252 40724
rect 15844 40672 15896 40724
rect 8944 40604 8996 40656
rect 9220 40604 9272 40656
rect 15108 40647 15160 40656
rect 15108 40613 15117 40647
rect 15117 40613 15151 40647
rect 15151 40613 15160 40647
rect 15108 40604 15160 40613
rect 7104 40579 7156 40588
rect 7104 40545 7113 40579
rect 7113 40545 7147 40579
rect 7147 40545 7156 40579
rect 7104 40536 7156 40545
rect 9128 40536 9180 40588
rect 5632 40511 5684 40520
rect 5632 40477 5641 40511
rect 5641 40477 5675 40511
rect 5675 40477 5684 40511
rect 5632 40468 5684 40477
rect 6828 40468 6880 40520
rect 9588 40511 9640 40520
rect 9588 40477 9597 40511
rect 9597 40477 9631 40511
rect 9631 40477 9640 40511
rect 9588 40468 9640 40477
rect 7012 40400 7064 40452
rect 8760 40400 8812 40452
rect 5264 40375 5316 40384
rect 5264 40341 5273 40375
rect 5273 40341 5307 40375
rect 5307 40341 5316 40375
rect 5264 40332 5316 40341
rect 6000 40332 6052 40384
rect 6644 40332 6696 40384
rect 7196 40332 7248 40384
rect 9036 40332 9088 40384
rect 12072 40468 12124 40520
rect 17960 40604 18012 40656
rect 20352 40715 20404 40724
rect 20352 40681 20361 40715
rect 20361 40681 20395 40715
rect 20395 40681 20404 40715
rect 20352 40672 20404 40681
rect 22468 40672 22520 40724
rect 25228 40672 25280 40724
rect 23388 40604 23440 40656
rect 24860 40604 24912 40656
rect 27620 40672 27672 40724
rect 28908 40672 28960 40724
rect 32496 40672 32548 40724
rect 35348 40672 35400 40724
rect 36912 40672 36964 40724
rect 38476 40715 38528 40724
rect 38476 40681 38485 40715
rect 38485 40681 38519 40715
rect 38519 40681 38528 40715
rect 38476 40672 38528 40681
rect 40684 40672 40736 40724
rect 17224 40536 17276 40588
rect 21088 40536 21140 40588
rect 11704 40400 11756 40452
rect 9864 40332 9916 40384
rect 14280 40400 14332 40452
rect 14556 40443 14608 40452
rect 14556 40409 14565 40443
rect 14565 40409 14599 40443
rect 14599 40409 14608 40443
rect 14556 40400 14608 40409
rect 14648 40443 14700 40452
rect 14648 40409 14657 40443
rect 14657 40409 14691 40443
rect 14691 40409 14700 40443
rect 14648 40400 14700 40409
rect 14740 40400 14792 40452
rect 14924 40400 14976 40452
rect 17132 40511 17184 40520
rect 17132 40477 17141 40511
rect 17141 40477 17175 40511
rect 17175 40477 17184 40511
rect 17132 40468 17184 40477
rect 20260 40511 20312 40520
rect 20260 40477 20269 40511
rect 20269 40477 20303 40511
rect 20303 40477 20312 40511
rect 22284 40536 22336 40588
rect 22560 40536 22612 40588
rect 20260 40468 20312 40477
rect 21548 40511 21600 40520
rect 21548 40477 21557 40511
rect 21557 40477 21591 40511
rect 21591 40477 21600 40511
rect 21548 40468 21600 40477
rect 23388 40468 23440 40520
rect 22284 40400 22336 40452
rect 23480 40400 23532 40452
rect 24860 40511 24912 40520
rect 24860 40477 24869 40511
rect 24869 40477 24903 40511
rect 24903 40477 24912 40511
rect 24860 40468 24912 40477
rect 26240 40536 26292 40588
rect 28724 40604 28776 40656
rect 26516 40536 26568 40588
rect 30564 40604 30616 40656
rect 32588 40604 32640 40656
rect 25964 40511 26016 40520
rect 25964 40477 25973 40511
rect 25973 40477 26007 40511
rect 26007 40477 26016 40511
rect 25964 40468 26016 40477
rect 26976 40511 27028 40520
rect 26976 40477 26985 40511
rect 26985 40477 27019 40511
rect 27019 40477 27028 40511
rect 26976 40468 27028 40477
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27068 40468 27120 40477
rect 27896 40511 27948 40520
rect 27896 40477 27905 40511
rect 27905 40477 27939 40511
rect 27939 40477 27948 40511
rect 27896 40468 27948 40477
rect 28080 40511 28132 40520
rect 28080 40477 28089 40511
rect 28089 40477 28123 40511
rect 28123 40477 28132 40511
rect 28080 40468 28132 40477
rect 24768 40400 24820 40452
rect 26148 40443 26200 40452
rect 26148 40409 26182 40443
rect 26182 40409 26200 40443
rect 26148 40400 26200 40409
rect 23848 40332 23900 40384
rect 24124 40332 24176 40384
rect 24216 40332 24268 40384
rect 25964 40332 26016 40384
rect 26792 40375 26844 40384
rect 26792 40341 26801 40375
rect 26801 40341 26835 40375
rect 26835 40341 26844 40375
rect 26792 40332 26844 40341
rect 27160 40443 27212 40452
rect 27160 40409 27169 40443
rect 27169 40409 27203 40443
rect 27203 40409 27212 40443
rect 27160 40400 27212 40409
rect 27252 40400 27304 40452
rect 28908 40536 28960 40588
rect 30288 40536 30340 40588
rect 31116 40536 31168 40588
rect 31668 40536 31720 40588
rect 28724 40511 28776 40520
rect 28724 40477 28733 40511
rect 28733 40477 28767 40511
rect 28767 40477 28776 40511
rect 28724 40468 28776 40477
rect 28816 40511 28868 40520
rect 28816 40477 28825 40511
rect 28825 40477 28859 40511
rect 28859 40477 28868 40511
rect 28816 40468 28868 40477
rect 29920 40468 29972 40520
rect 30656 40511 30708 40520
rect 30656 40477 30665 40511
rect 30665 40477 30699 40511
rect 30699 40477 30708 40511
rect 30656 40468 30708 40477
rect 31852 40468 31904 40520
rect 29092 40443 29144 40452
rect 29092 40409 29101 40443
rect 29101 40409 29135 40443
rect 29135 40409 29144 40443
rect 29092 40400 29144 40409
rect 29184 40443 29236 40452
rect 29184 40409 29193 40443
rect 29193 40409 29227 40443
rect 29227 40409 29236 40443
rect 29184 40400 29236 40409
rect 28540 40375 28592 40384
rect 28540 40341 28549 40375
rect 28549 40341 28583 40375
rect 28583 40341 28592 40375
rect 28540 40332 28592 40341
rect 29828 40375 29880 40384
rect 29828 40341 29837 40375
rect 29837 40341 29871 40375
rect 29871 40341 29880 40375
rect 29828 40332 29880 40341
rect 30656 40332 30708 40384
rect 31484 40332 31536 40384
rect 32036 40511 32088 40520
rect 32036 40477 32045 40511
rect 32045 40477 32079 40511
rect 32079 40477 32088 40511
rect 32036 40468 32088 40477
rect 33048 40468 33100 40520
rect 33600 40468 33652 40520
rect 34796 40468 34848 40520
rect 34980 40511 35032 40520
rect 34980 40477 34989 40511
rect 34989 40477 35023 40511
rect 35023 40477 35032 40511
rect 34980 40468 35032 40477
rect 40132 40579 40184 40588
rect 40132 40545 40141 40579
rect 40141 40545 40175 40579
rect 40175 40545 40184 40579
rect 40132 40536 40184 40545
rect 35900 40511 35952 40520
rect 35900 40477 35909 40511
rect 35909 40477 35943 40511
rect 35943 40477 35952 40511
rect 35900 40468 35952 40477
rect 32128 40332 32180 40384
rect 33784 40400 33836 40452
rect 35624 40400 35676 40452
rect 38384 40511 38436 40520
rect 38384 40477 38393 40511
rect 38393 40477 38427 40511
rect 38427 40477 38436 40511
rect 38384 40468 38436 40477
rect 38568 40511 38620 40520
rect 38568 40477 38577 40511
rect 38577 40477 38611 40511
rect 38611 40477 38620 40511
rect 38568 40468 38620 40477
rect 38844 40468 38896 40520
rect 41880 40511 41932 40520
rect 41880 40477 41889 40511
rect 41889 40477 41923 40511
rect 41923 40477 41932 40511
rect 41880 40468 41932 40477
rect 42616 40400 42668 40452
rect 42892 40332 42944 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 6000 40171 6052 40180
rect 6000 40137 6009 40171
rect 6009 40137 6043 40171
rect 6043 40137 6052 40171
rect 6000 40128 6052 40137
rect 8392 40171 8444 40180
rect 8392 40137 8401 40171
rect 8401 40137 8435 40171
rect 8435 40137 8444 40171
rect 8392 40128 8444 40137
rect 9036 40128 9088 40180
rect 11980 40128 12032 40180
rect 12164 40171 12216 40180
rect 12164 40137 12173 40171
rect 12173 40137 12207 40171
rect 12207 40137 12216 40171
rect 12164 40128 12216 40137
rect 14372 40128 14424 40180
rect 5264 40060 5316 40112
rect 6828 40060 6880 40112
rect 9864 40060 9916 40112
rect 10048 40060 10100 40112
rect 9680 39992 9732 40044
rect 7104 39967 7156 39976
rect 7104 39933 7113 39967
rect 7113 39933 7147 39967
rect 7147 39933 7156 39967
rect 7104 39924 7156 39933
rect 8944 39967 8996 39976
rect 8944 39933 8953 39967
rect 8953 39933 8987 39967
rect 8987 39933 8996 39967
rect 8944 39924 8996 39933
rect 9956 39967 10008 39976
rect 9956 39933 9965 39967
rect 9965 39933 9999 39967
rect 9999 39933 10008 39967
rect 9956 39924 10008 39933
rect 13728 39992 13780 40044
rect 10692 39967 10744 39976
rect 10692 39933 10701 39967
rect 10701 39933 10735 39967
rect 10735 39933 10744 39967
rect 10692 39924 10744 39933
rect 12440 39924 12492 39976
rect 14280 39924 14332 39976
rect 17132 39856 17184 39908
rect 17776 40035 17828 40044
rect 17776 40001 17785 40035
rect 17785 40001 17819 40035
rect 17819 40001 17828 40035
rect 17776 39992 17828 40001
rect 18236 40060 18288 40112
rect 23848 40128 23900 40180
rect 24124 40128 24176 40180
rect 24952 40128 25004 40180
rect 26240 40128 26292 40180
rect 27068 40128 27120 40180
rect 27436 40128 27488 40180
rect 28080 40128 28132 40180
rect 33692 40128 33744 40180
rect 34704 40128 34756 40180
rect 42616 40171 42668 40180
rect 42616 40137 42625 40171
rect 42625 40137 42659 40171
rect 42659 40137 42668 40171
rect 42616 40128 42668 40137
rect 20260 40060 20312 40112
rect 22284 40035 22336 40044
rect 22284 40001 22293 40035
rect 22293 40001 22327 40035
rect 22327 40001 22336 40035
rect 22284 39992 22336 40001
rect 22376 40035 22428 40044
rect 22376 40001 22385 40035
rect 22385 40001 22419 40035
rect 22419 40001 22428 40035
rect 22376 39992 22428 40001
rect 22836 39992 22888 40044
rect 23388 40035 23440 40044
rect 23388 40001 23397 40035
rect 23397 40001 23431 40035
rect 23431 40001 23440 40035
rect 23388 39992 23440 40001
rect 24216 39992 24268 40044
rect 24676 39992 24728 40044
rect 24768 39992 24820 40044
rect 26148 39992 26200 40044
rect 27252 40060 27304 40112
rect 18328 39924 18380 39976
rect 23940 39967 23992 39976
rect 23940 39933 23949 39967
rect 23949 39933 23983 39967
rect 23983 39933 23992 39967
rect 23940 39924 23992 39933
rect 25044 39924 25096 39976
rect 18236 39856 18288 39908
rect 4620 39788 4672 39840
rect 5540 39788 5592 39840
rect 6552 39831 6604 39840
rect 6552 39797 6561 39831
rect 6561 39797 6595 39831
rect 6595 39797 6604 39831
rect 6552 39788 6604 39797
rect 11796 39788 11848 39840
rect 18880 39788 18932 39840
rect 24584 39856 24636 39908
rect 25320 39788 25372 39840
rect 27160 39992 27212 40044
rect 27068 39924 27120 39976
rect 29000 40060 29052 40112
rect 29828 40060 29880 40112
rect 30288 40060 30340 40112
rect 27620 40035 27672 40044
rect 27620 40001 27629 40035
rect 27629 40001 27663 40035
rect 27663 40001 27672 40035
rect 27620 39992 27672 40001
rect 29184 39992 29236 40044
rect 30196 40035 30248 40044
rect 30196 40001 30205 40035
rect 30205 40001 30239 40035
rect 30239 40001 30248 40035
rect 30196 39992 30248 40001
rect 31024 40035 31076 40044
rect 31024 40001 31033 40035
rect 31033 40001 31067 40035
rect 31067 40001 31076 40035
rect 31024 39992 31076 40001
rect 31484 40035 31536 40044
rect 31484 40001 31493 40035
rect 31493 40001 31527 40035
rect 31527 40001 31536 40035
rect 31484 39992 31536 40001
rect 33508 40060 33560 40112
rect 34612 40060 34664 40112
rect 38660 40060 38712 40112
rect 38844 40060 38896 40112
rect 42892 40060 42944 40112
rect 34520 40035 34572 40044
rect 34520 40001 34554 40035
rect 34554 40001 34572 40035
rect 34520 39992 34572 40001
rect 28172 39924 28224 39976
rect 28816 39924 28868 39976
rect 32772 39924 32824 39976
rect 32864 39967 32916 39976
rect 32864 39933 32873 39967
rect 32873 39933 32907 39967
rect 32907 39933 32916 39967
rect 32864 39924 32916 39933
rect 43076 39967 43128 39976
rect 43076 39933 43085 39967
rect 43085 39933 43119 39967
rect 43119 39933 43128 39967
rect 43076 39924 43128 39933
rect 43168 39967 43220 39976
rect 43168 39933 43177 39967
rect 43177 39933 43211 39967
rect 43211 39933 43220 39967
rect 43168 39924 43220 39933
rect 27252 39856 27304 39908
rect 26608 39788 26660 39840
rect 31760 39788 31812 39840
rect 36452 39856 36504 39908
rect 39304 39856 39356 39908
rect 40408 39856 40460 39908
rect 34428 39788 34480 39840
rect 34612 39788 34664 39840
rect 34980 39788 35032 39840
rect 38568 39831 38620 39840
rect 38568 39797 38577 39831
rect 38577 39797 38611 39831
rect 38611 39797 38620 39831
rect 38568 39788 38620 39797
rect 38936 39788 38988 39840
rect 40132 39788 40184 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 18328 39627 18380 39636
rect 18328 39593 18337 39627
rect 18337 39593 18371 39627
rect 18371 39593 18380 39627
rect 18328 39584 18380 39593
rect 6736 39448 6788 39500
rect 9956 39448 10008 39500
rect 6644 39423 6696 39432
rect 6644 39389 6653 39423
rect 6653 39389 6687 39423
rect 6687 39389 6696 39423
rect 6644 39380 6696 39389
rect 7380 39380 7432 39432
rect 10416 39423 10468 39432
rect 10416 39389 10425 39423
rect 10425 39389 10459 39423
rect 10459 39389 10468 39423
rect 10416 39380 10468 39389
rect 16856 39448 16908 39500
rect 17684 39448 17736 39500
rect 20168 39516 20220 39568
rect 21180 39627 21232 39636
rect 21180 39593 21189 39627
rect 21189 39593 21223 39627
rect 21223 39593 21232 39627
rect 21180 39584 21232 39593
rect 24032 39627 24084 39636
rect 24032 39593 24041 39627
rect 24041 39593 24075 39627
rect 24075 39593 24084 39627
rect 24032 39584 24084 39593
rect 27620 39627 27672 39636
rect 27620 39593 27629 39627
rect 27629 39593 27663 39627
rect 27663 39593 27672 39627
rect 27620 39584 27672 39593
rect 31668 39584 31720 39636
rect 33048 39627 33100 39636
rect 11336 39380 11388 39432
rect 15752 39380 15804 39432
rect 7104 39355 7156 39364
rect 7104 39321 7113 39355
rect 7113 39321 7147 39355
rect 7147 39321 7156 39355
rect 7104 39312 7156 39321
rect 10232 39312 10284 39364
rect 11888 39355 11940 39364
rect 11888 39321 11897 39355
rect 11897 39321 11931 39355
rect 11931 39321 11940 39355
rect 11888 39312 11940 39321
rect 14740 39312 14792 39364
rect 16488 39380 16540 39432
rect 17960 39380 18012 39432
rect 18420 39423 18472 39432
rect 18420 39389 18429 39423
rect 18429 39389 18463 39423
rect 18463 39389 18472 39423
rect 18420 39380 18472 39389
rect 20076 39380 20128 39432
rect 20812 39423 20864 39432
rect 20812 39389 20821 39423
rect 20821 39389 20855 39423
rect 20855 39389 20864 39423
rect 20812 39380 20864 39389
rect 28540 39516 28592 39568
rect 33048 39593 33057 39627
rect 33057 39593 33091 39627
rect 33091 39593 33100 39627
rect 33048 39584 33100 39593
rect 34520 39584 34572 39636
rect 34888 39584 34940 39636
rect 27160 39448 27212 39500
rect 27344 39448 27396 39500
rect 29092 39448 29144 39500
rect 21088 39380 21140 39432
rect 22928 39423 22980 39432
rect 22928 39389 22937 39423
rect 22937 39389 22971 39423
rect 22971 39389 22980 39423
rect 22928 39380 22980 39389
rect 23112 39423 23164 39432
rect 23112 39389 23121 39423
rect 23121 39389 23155 39423
rect 23155 39389 23164 39423
rect 23112 39380 23164 39389
rect 23756 39423 23808 39432
rect 23756 39389 23765 39423
rect 23765 39389 23799 39423
rect 23799 39389 23808 39423
rect 23756 39380 23808 39389
rect 11980 39244 12032 39296
rect 16304 39287 16356 39296
rect 16304 39253 16313 39287
rect 16313 39253 16347 39287
rect 16347 39253 16356 39287
rect 16304 39244 16356 39253
rect 16948 39312 17000 39364
rect 18052 39244 18104 39296
rect 20260 39287 20312 39296
rect 20260 39253 20269 39287
rect 20269 39253 20303 39287
rect 20303 39253 20312 39287
rect 20260 39244 20312 39253
rect 27896 39380 27948 39432
rect 30104 39423 30156 39432
rect 30104 39389 30113 39423
rect 30113 39389 30147 39423
rect 30147 39389 30156 39423
rect 30104 39380 30156 39389
rect 31300 39448 31352 39500
rect 31944 39491 31996 39500
rect 31944 39457 31953 39491
rect 31953 39457 31987 39491
rect 31987 39457 31996 39491
rect 31944 39448 31996 39457
rect 33784 39516 33836 39568
rect 38384 39584 38436 39636
rect 39212 39584 39264 39636
rect 40960 39584 41012 39636
rect 41420 39584 41472 39636
rect 23020 39287 23072 39296
rect 23020 39253 23029 39287
rect 23029 39253 23063 39287
rect 23063 39253 23072 39287
rect 24952 39312 25004 39364
rect 28264 39312 28316 39364
rect 31576 39380 31628 39432
rect 32036 39423 32088 39432
rect 32036 39389 32045 39423
rect 32045 39389 32079 39423
rect 32079 39389 32088 39423
rect 32036 39380 32088 39389
rect 34060 39380 34112 39432
rect 34152 39423 34204 39432
rect 34152 39389 34161 39423
rect 34161 39389 34195 39423
rect 34195 39389 34204 39423
rect 34152 39380 34204 39389
rect 34428 39380 34480 39432
rect 34888 39380 34940 39432
rect 36636 39448 36688 39500
rect 37004 39448 37056 39500
rect 31760 39355 31812 39364
rect 31760 39321 31769 39355
rect 31769 39321 31803 39355
rect 31803 39321 31812 39355
rect 31760 39312 31812 39321
rect 32864 39312 32916 39364
rect 36084 39312 36136 39364
rect 37096 39423 37148 39432
rect 37096 39389 37105 39423
rect 37105 39389 37139 39423
rect 37139 39389 37148 39423
rect 37096 39380 37148 39389
rect 37188 39423 37240 39432
rect 37188 39389 37198 39423
rect 37198 39389 37232 39423
rect 37232 39389 37240 39423
rect 37188 39380 37240 39389
rect 39672 39516 39724 39568
rect 37740 39448 37792 39500
rect 37924 39380 37976 39432
rect 38936 39423 38988 39432
rect 38936 39389 38945 39423
rect 38945 39389 38979 39423
rect 38979 39389 38988 39423
rect 38936 39380 38988 39389
rect 38660 39355 38712 39364
rect 38660 39321 38669 39355
rect 38669 39321 38703 39355
rect 38703 39321 38712 39355
rect 38660 39312 38712 39321
rect 38844 39355 38896 39364
rect 38844 39321 38853 39355
rect 38853 39321 38887 39355
rect 38887 39321 38896 39355
rect 38844 39312 38896 39321
rect 23020 39244 23072 39253
rect 30564 39287 30616 39296
rect 30564 39253 30573 39287
rect 30573 39253 30607 39287
rect 30607 39253 30616 39287
rect 30564 39244 30616 39253
rect 34704 39244 34756 39296
rect 37280 39244 37332 39296
rect 41788 39380 41840 39432
rect 42708 39380 42760 39432
rect 39120 39312 39172 39364
rect 43996 39312 44048 39364
rect 41328 39244 41380 39296
rect 41420 39287 41472 39296
rect 41420 39253 41429 39287
rect 41429 39253 41463 39287
rect 41463 39253 41472 39287
rect 41420 39244 41472 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 6736 38972 6788 39024
rect 5816 38947 5868 38956
rect 5816 38913 5825 38947
rect 5825 38913 5859 38947
rect 5859 38913 5868 38947
rect 5816 38904 5868 38913
rect 5908 38904 5960 38956
rect 6552 38904 6604 38956
rect 7380 38947 7432 38956
rect 7380 38913 7389 38947
rect 7389 38913 7423 38947
rect 7423 38913 7432 38947
rect 7380 38904 7432 38913
rect 8760 39015 8812 39024
rect 8760 38981 8769 39015
rect 8769 38981 8803 39015
rect 8803 38981 8812 39015
rect 8760 38972 8812 38981
rect 12992 38972 13044 39024
rect 9956 38947 10008 38956
rect 9956 38913 9965 38947
rect 9965 38913 9999 38947
rect 9999 38913 10008 38947
rect 9956 38904 10008 38913
rect 10416 38904 10468 38956
rect 11796 38904 11848 38956
rect 6736 38836 6788 38888
rect 12808 38904 12860 38956
rect 16948 39083 17000 39092
rect 16948 39049 16957 39083
rect 16957 39049 16991 39083
rect 16991 39049 17000 39083
rect 16948 39040 17000 39049
rect 17408 39040 17460 39092
rect 20076 39083 20128 39092
rect 20076 39049 20085 39083
rect 20085 39049 20119 39083
rect 20119 39049 20128 39083
rect 20076 39040 20128 39049
rect 21088 39040 21140 39092
rect 21548 39040 21600 39092
rect 20996 38972 21048 39024
rect 26516 39083 26568 39092
rect 26516 39049 26525 39083
rect 26525 39049 26559 39083
rect 26559 39049 26568 39083
rect 26516 39040 26568 39049
rect 27160 39083 27212 39092
rect 27160 39049 27169 39083
rect 27169 39049 27203 39083
rect 27203 39049 27212 39083
rect 27160 39040 27212 39049
rect 11428 38768 11480 38820
rect 13084 38836 13136 38888
rect 14004 38904 14056 38956
rect 15108 38904 15160 38956
rect 12440 38768 12492 38820
rect 14740 38768 14792 38820
rect 16856 38947 16908 38956
rect 16856 38913 16865 38947
rect 16865 38913 16899 38947
rect 16899 38913 16908 38947
rect 16856 38904 16908 38913
rect 16580 38836 16632 38888
rect 18788 38947 18840 38956
rect 18788 38913 18797 38947
rect 18797 38913 18831 38947
rect 18831 38913 18840 38947
rect 18788 38904 18840 38913
rect 18880 38947 18932 38956
rect 18880 38913 18889 38947
rect 18889 38913 18923 38947
rect 18923 38913 18932 38947
rect 18880 38904 18932 38913
rect 19432 38947 19484 38956
rect 19432 38913 19441 38947
rect 19441 38913 19475 38947
rect 19475 38913 19484 38947
rect 19432 38904 19484 38913
rect 19524 38904 19576 38956
rect 19984 38904 20036 38956
rect 21180 38904 21232 38956
rect 23480 38904 23532 38956
rect 24492 38947 24544 38956
rect 24492 38913 24501 38947
rect 24501 38913 24535 38947
rect 24535 38913 24544 38947
rect 24492 38904 24544 38913
rect 24952 38947 25004 38956
rect 24952 38913 24961 38947
rect 24961 38913 24995 38947
rect 24995 38913 25004 38947
rect 24952 38904 25004 38913
rect 26056 38904 26108 38956
rect 16304 38768 16356 38820
rect 20904 38836 20956 38888
rect 7012 38700 7064 38752
rect 7288 38700 7340 38752
rect 9036 38700 9088 38752
rect 14188 38700 14240 38752
rect 14832 38700 14884 38752
rect 21180 38768 21232 38820
rect 23204 38768 23256 38820
rect 23388 38879 23440 38888
rect 23388 38845 23397 38879
rect 23397 38845 23431 38879
rect 23431 38845 23440 38879
rect 23388 38836 23440 38845
rect 26424 38836 26476 38888
rect 25044 38768 25096 38820
rect 26056 38768 26108 38820
rect 26976 38904 27028 38956
rect 27988 38972 28040 39024
rect 28816 38972 28868 39024
rect 27804 38904 27856 38956
rect 28540 38904 28592 38956
rect 32128 39040 32180 39092
rect 32772 39040 32824 39092
rect 31300 38972 31352 39024
rect 33968 38972 34020 39024
rect 36544 39015 36596 39024
rect 36544 38981 36553 39015
rect 36553 38981 36587 39015
rect 36587 38981 36596 39015
rect 36544 38972 36596 38981
rect 36728 39040 36780 39092
rect 37556 39040 37608 39092
rect 37924 39040 37976 39092
rect 38936 39040 38988 39092
rect 39120 39083 39172 39092
rect 39120 39049 39129 39083
rect 39129 39049 39163 39083
rect 39163 39049 39172 39083
rect 39120 39040 39172 39049
rect 29644 38879 29696 38888
rect 29644 38845 29653 38879
rect 29653 38845 29687 38879
rect 29687 38845 29696 38879
rect 29644 38836 29696 38845
rect 30472 38904 30524 38956
rect 31760 38904 31812 38956
rect 32312 38904 32364 38956
rect 33784 38904 33836 38956
rect 33876 38947 33928 38956
rect 33876 38913 33885 38947
rect 33885 38913 33919 38947
rect 33919 38913 33928 38947
rect 33876 38904 33928 38913
rect 34796 38947 34848 38956
rect 34796 38913 34805 38947
rect 34805 38913 34839 38947
rect 34839 38913 34848 38947
rect 34796 38904 34848 38913
rect 36268 38947 36320 38956
rect 36268 38913 36277 38947
rect 36277 38913 36311 38947
rect 36311 38913 36320 38947
rect 36268 38904 36320 38913
rect 36452 38947 36504 38956
rect 36452 38913 36459 38947
rect 36459 38913 36504 38947
rect 36452 38904 36504 38913
rect 37740 39015 37792 39024
rect 37740 38981 37749 39015
rect 37749 38981 37783 39015
rect 37783 38981 37792 39015
rect 37740 38972 37792 38981
rect 37372 38904 37424 38956
rect 37648 38947 37700 38956
rect 37648 38913 37655 38947
rect 37655 38913 37700 38947
rect 37648 38904 37700 38913
rect 20260 38700 20312 38752
rect 24216 38700 24268 38752
rect 24584 38743 24636 38752
rect 24584 38709 24593 38743
rect 24593 38709 24627 38743
rect 24627 38709 24636 38743
rect 24584 38700 24636 38709
rect 26148 38743 26200 38752
rect 26148 38709 26157 38743
rect 26157 38709 26191 38743
rect 26191 38709 26200 38743
rect 26148 38700 26200 38709
rect 27712 38768 27764 38820
rect 28080 38768 28132 38820
rect 28724 38768 28776 38820
rect 30104 38768 30156 38820
rect 31668 38836 31720 38888
rect 32680 38768 32732 38820
rect 36084 38836 36136 38888
rect 36912 38836 36964 38888
rect 37924 38947 37976 38956
rect 37924 38913 37938 38947
rect 37938 38913 37972 38947
rect 37972 38913 37976 38947
rect 37924 38904 37976 38913
rect 38568 38904 38620 38956
rect 39212 38947 39264 38956
rect 39212 38913 39221 38947
rect 39221 38913 39255 38947
rect 39255 38913 39264 38947
rect 39212 38904 39264 38913
rect 42984 38947 43036 38956
rect 42984 38913 42993 38947
rect 42993 38913 43027 38947
rect 43027 38913 43036 38947
rect 42984 38904 43036 38913
rect 39764 38836 39816 38888
rect 42708 38836 42760 38888
rect 43168 38879 43220 38888
rect 43168 38845 43177 38879
rect 43177 38845 43211 38879
rect 43211 38845 43220 38879
rect 43168 38836 43220 38845
rect 34704 38768 34756 38820
rect 36728 38768 36780 38820
rect 39212 38768 39264 38820
rect 29000 38743 29052 38752
rect 29000 38709 29009 38743
rect 29009 38709 29043 38743
rect 29043 38709 29052 38743
rect 29000 38700 29052 38709
rect 31300 38700 31352 38752
rect 33048 38700 33100 38752
rect 35532 38700 35584 38752
rect 37188 38700 37240 38752
rect 40960 38700 41012 38752
rect 42616 38743 42668 38752
rect 42616 38709 42625 38743
rect 42625 38709 42659 38743
rect 42659 38709 42668 38743
rect 42616 38700 42668 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 12348 38496 12400 38548
rect 5816 38335 5868 38344
rect 5816 38301 5825 38335
rect 5825 38301 5859 38335
rect 5859 38301 5868 38335
rect 5816 38292 5868 38301
rect 5908 38335 5960 38344
rect 5908 38301 5917 38335
rect 5917 38301 5951 38335
rect 5951 38301 5960 38335
rect 5908 38292 5960 38301
rect 7012 38335 7064 38344
rect 7012 38301 7021 38335
rect 7021 38301 7055 38335
rect 7055 38301 7064 38335
rect 7012 38292 7064 38301
rect 7196 38292 7248 38344
rect 10140 38403 10192 38412
rect 10140 38369 10149 38403
rect 10149 38369 10183 38403
rect 10183 38369 10192 38403
rect 10140 38360 10192 38369
rect 14280 38428 14332 38480
rect 17960 38496 18012 38548
rect 19524 38496 19576 38548
rect 19892 38496 19944 38548
rect 19984 38496 20036 38548
rect 20812 38496 20864 38548
rect 21180 38539 21232 38548
rect 21180 38505 21189 38539
rect 21189 38505 21223 38539
rect 21223 38505 21232 38539
rect 21180 38496 21232 38505
rect 21364 38539 21416 38548
rect 21364 38505 21373 38539
rect 21373 38505 21407 38539
rect 21407 38505 21416 38539
rect 21364 38496 21416 38505
rect 23940 38539 23992 38548
rect 23940 38505 23949 38539
rect 23949 38505 23983 38539
rect 23983 38505 23992 38539
rect 23940 38496 23992 38505
rect 24860 38539 24912 38548
rect 24860 38505 24869 38539
rect 24869 38505 24903 38539
rect 24903 38505 24912 38539
rect 24860 38496 24912 38505
rect 7932 38335 7984 38344
rect 7932 38301 7941 38335
rect 7941 38301 7975 38335
rect 7975 38301 7984 38335
rect 7932 38292 7984 38301
rect 8116 38335 8168 38344
rect 8116 38301 8125 38335
rect 8125 38301 8159 38335
rect 8159 38301 8168 38335
rect 8116 38292 8168 38301
rect 8760 38292 8812 38344
rect 6184 38224 6236 38276
rect 11152 38292 11204 38344
rect 8208 38156 8260 38208
rect 11980 38224 12032 38276
rect 12624 38224 12676 38276
rect 14096 38360 14148 38412
rect 15108 38360 15160 38412
rect 13452 38335 13504 38344
rect 13452 38301 13461 38335
rect 13461 38301 13495 38335
rect 13495 38301 13504 38335
rect 13452 38292 13504 38301
rect 12900 38224 12952 38276
rect 14740 38335 14792 38344
rect 14740 38301 14749 38335
rect 14749 38301 14783 38335
rect 14783 38301 14792 38335
rect 14740 38292 14792 38301
rect 16856 38360 16908 38412
rect 17132 38360 17184 38412
rect 16396 38335 16448 38344
rect 16396 38301 16405 38335
rect 16405 38301 16439 38335
rect 16439 38301 16448 38335
rect 16396 38292 16448 38301
rect 16488 38335 16540 38344
rect 16488 38301 16497 38335
rect 16497 38301 16531 38335
rect 16531 38301 16540 38335
rect 16488 38292 16540 38301
rect 17684 38335 17736 38344
rect 17684 38301 17693 38335
rect 17693 38301 17727 38335
rect 17727 38301 17736 38335
rect 17684 38292 17736 38301
rect 18696 38335 18748 38344
rect 18696 38301 18705 38335
rect 18705 38301 18739 38335
rect 18739 38301 18748 38335
rect 18696 38292 18748 38301
rect 18880 38335 18932 38344
rect 18880 38301 18889 38335
rect 18889 38301 18923 38335
rect 18923 38301 18932 38335
rect 18880 38292 18932 38301
rect 16856 38224 16908 38276
rect 13084 38156 13136 38208
rect 13268 38199 13320 38208
rect 13268 38165 13277 38199
rect 13277 38165 13311 38199
rect 13311 38165 13320 38199
rect 13268 38156 13320 38165
rect 13360 38199 13412 38208
rect 13360 38165 13369 38199
rect 13369 38165 13403 38199
rect 13403 38165 13412 38199
rect 13360 38156 13412 38165
rect 13820 38156 13872 38208
rect 16672 38199 16724 38208
rect 16672 38165 16681 38199
rect 16681 38165 16715 38199
rect 16715 38165 16724 38199
rect 16672 38156 16724 38165
rect 19340 38156 19392 38208
rect 19800 38335 19852 38344
rect 19800 38301 19809 38335
rect 19809 38301 19843 38335
rect 19843 38301 19852 38335
rect 19800 38292 19852 38301
rect 19892 38224 19944 38276
rect 20076 38224 20128 38276
rect 20352 38360 20404 38412
rect 20260 38335 20312 38344
rect 20260 38301 20269 38335
rect 20269 38301 20303 38335
rect 20303 38301 20312 38335
rect 20260 38292 20312 38301
rect 20628 38292 20680 38344
rect 23020 38360 23072 38412
rect 25872 38428 25924 38480
rect 29000 38428 29052 38480
rect 31024 38428 31076 38480
rect 31944 38428 31996 38480
rect 20628 38156 20680 38208
rect 22928 38292 22980 38344
rect 24308 38292 24360 38344
rect 25964 38292 26016 38344
rect 25136 38156 25188 38208
rect 25228 38199 25280 38208
rect 25228 38165 25237 38199
rect 25237 38165 25271 38199
rect 25271 38165 25280 38199
rect 25228 38156 25280 38165
rect 28540 38360 28592 38412
rect 28908 38360 28960 38412
rect 30012 38360 30064 38412
rect 37096 38496 37148 38548
rect 38660 38496 38712 38548
rect 43076 38496 43128 38548
rect 36176 38360 36228 38412
rect 27068 38335 27120 38344
rect 27068 38301 27077 38335
rect 27077 38301 27111 38335
rect 27111 38301 27120 38335
rect 27068 38292 27120 38301
rect 27160 38335 27212 38344
rect 27160 38301 27169 38335
rect 27169 38301 27203 38335
rect 27203 38301 27212 38335
rect 27160 38292 27212 38301
rect 28172 38292 28224 38344
rect 28448 38292 28500 38344
rect 30104 38292 30156 38344
rect 30472 38335 30524 38344
rect 30472 38301 30481 38335
rect 30481 38301 30515 38335
rect 30515 38301 30524 38335
rect 30472 38292 30524 38301
rect 31392 38292 31444 38344
rect 31576 38292 31628 38344
rect 31760 38335 31812 38344
rect 31760 38301 31769 38335
rect 31769 38301 31803 38335
rect 31803 38301 31812 38335
rect 31760 38292 31812 38301
rect 32680 38335 32732 38344
rect 32680 38301 32689 38335
rect 32689 38301 32723 38335
rect 32723 38301 32732 38335
rect 32680 38292 32732 38301
rect 32772 38335 32824 38344
rect 32772 38301 32781 38335
rect 32781 38301 32815 38335
rect 32815 38301 32824 38335
rect 32772 38292 32824 38301
rect 27528 38224 27580 38276
rect 28264 38156 28316 38208
rect 31668 38267 31720 38276
rect 31668 38233 31677 38267
rect 31677 38233 31711 38267
rect 31711 38233 31720 38267
rect 31668 38224 31720 38233
rect 33048 38335 33100 38344
rect 33048 38301 33057 38335
rect 33057 38301 33091 38335
rect 33091 38301 33100 38335
rect 33048 38292 33100 38301
rect 34244 38335 34296 38344
rect 34244 38301 34253 38335
rect 34253 38301 34287 38335
rect 34287 38301 34296 38335
rect 34244 38292 34296 38301
rect 34428 38292 34480 38344
rect 35072 38335 35124 38344
rect 35072 38301 35081 38335
rect 35081 38301 35115 38335
rect 35115 38301 35124 38335
rect 35072 38292 35124 38301
rect 36084 38292 36136 38344
rect 36360 38335 36412 38344
rect 36360 38301 36370 38335
rect 36370 38301 36404 38335
rect 36404 38301 36412 38335
rect 36360 38292 36412 38301
rect 36728 38335 36780 38344
rect 36728 38301 36742 38335
rect 36742 38301 36776 38335
rect 36776 38301 36780 38335
rect 36728 38292 36780 38301
rect 37464 38335 37516 38344
rect 37464 38301 37473 38335
rect 37473 38301 37507 38335
rect 37507 38301 37516 38335
rect 37464 38292 37516 38301
rect 37648 38335 37700 38344
rect 37648 38301 37655 38335
rect 37655 38301 37700 38335
rect 37648 38292 37700 38301
rect 32404 38199 32456 38208
rect 32404 38165 32413 38199
rect 32413 38165 32447 38199
rect 32447 38165 32456 38199
rect 32404 38156 32456 38165
rect 33600 38224 33652 38276
rect 33784 38267 33836 38276
rect 33784 38233 33793 38267
rect 33793 38233 33827 38267
rect 33827 38233 33836 38267
rect 33784 38224 33836 38233
rect 34520 38224 34572 38276
rect 32864 38156 32916 38208
rect 34796 38156 34848 38208
rect 35992 38156 36044 38208
rect 36820 38224 36872 38276
rect 37004 38224 37056 38276
rect 37740 38267 37792 38276
rect 37740 38233 37749 38267
rect 37749 38233 37783 38267
rect 37783 38233 37792 38267
rect 37740 38224 37792 38233
rect 37924 38335 37976 38344
rect 37924 38301 37938 38335
rect 37938 38301 37972 38335
rect 37972 38301 37976 38335
rect 37924 38292 37976 38301
rect 38660 38224 38712 38276
rect 36912 38156 36964 38208
rect 39212 38335 39264 38344
rect 39212 38301 39221 38335
rect 39221 38301 39255 38335
rect 39255 38301 39264 38335
rect 39212 38292 39264 38301
rect 39304 38335 39356 38344
rect 39304 38301 39313 38335
rect 39313 38301 39347 38335
rect 39347 38301 39356 38335
rect 39304 38292 39356 38301
rect 39120 38267 39172 38276
rect 39120 38233 39129 38267
rect 39129 38233 39163 38267
rect 39163 38233 39172 38267
rect 39120 38224 39172 38233
rect 40408 38335 40460 38344
rect 40408 38301 40417 38335
rect 40417 38301 40451 38335
rect 40451 38301 40460 38335
rect 40408 38292 40460 38301
rect 41144 38292 41196 38344
rect 41788 38403 41840 38412
rect 41788 38369 41797 38403
rect 41797 38369 41831 38403
rect 41831 38369 41840 38403
rect 41788 38360 41840 38369
rect 42616 38292 42668 38344
rect 39212 38156 39264 38208
rect 42892 38224 42944 38276
rect 40408 38156 40460 38208
rect 43076 38156 43128 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4620 37884 4672 37936
rect 7012 37884 7064 37936
rect 4896 37816 4948 37868
rect 7196 37816 7248 37868
rect 7840 37816 7892 37868
rect 9588 37952 9640 38004
rect 12624 37952 12676 38004
rect 14004 37952 14056 38004
rect 18696 37952 18748 38004
rect 19340 37952 19392 38004
rect 23480 37952 23532 38004
rect 24860 37952 24912 38004
rect 8116 37859 8168 37868
rect 8116 37825 8125 37859
rect 8125 37825 8159 37859
rect 8159 37825 8168 37859
rect 8116 37816 8168 37825
rect 9864 37884 9916 37936
rect 10232 37884 10284 37936
rect 9036 37859 9088 37868
rect 9036 37825 9045 37859
rect 9045 37825 9079 37859
rect 9079 37825 9088 37859
rect 9036 37816 9088 37825
rect 10416 37816 10468 37868
rect 10508 37816 10560 37868
rect 9496 37748 9548 37800
rect 9680 37680 9732 37732
rect 5540 37612 5592 37664
rect 7380 37612 7432 37664
rect 10508 37680 10560 37732
rect 10692 37791 10744 37800
rect 10692 37757 10701 37791
rect 10701 37757 10735 37791
rect 10735 37757 10744 37791
rect 10692 37748 10744 37757
rect 11060 37816 11112 37868
rect 11428 37748 11480 37800
rect 9864 37612 9916 37664
rect 10692 37612 10744 37664
rect 11520 37612 11572 37664
rect 11612 37612 11664 37664
rect 12348 37816 12400 37868
rect 12808 37816 12860 37868
rect 13084 37816 13136 37868
rect 13820 37859 13872 37868
rect 13820 37825 13829 37859
rect 13829 37825 13863 37859
rect 13863 37825 13872 37859
rect 13820 37816 13872 37825
rect 14004 37859 14056 37868
rect 14004 37825 14013 37859
rect 14013 37825 14047 37859
rect 14047 37825 14056 37859
rect 14004 37816 14056 37825
rect 14096 37859 14148 37868
rect 14096 37825 14105 37859
rect 14105 37825 14139 37859
rect 14139 37825 14148 37859
rect 14096 37816 14148 37825
rect 16672 37884 16724 37936
rect 14832 37816 14884 37868
rect 15936 37859 15988 37868
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 16580 37816 16632 37868
rect 14188 37791 14240 37800
rect 14188 37757 14197 37791
rect 14197 37757 14231 37791
rect 14231 37757 14240 37791
rect 14188 37748 14240 37757
rect 12716 37680 12768 37732
rect 15108 37680 15160 37732
rect 15752 37723 15804 37732
rect 15752 37689 15761 37723
rect 15761 37689 15795 37723
rect 15795 37689 15804 37723
rect 15752 37680 15804 37689
rect 16488 37748 16540 37800
rect 16948 37816 17000 37868
rect 17960 37859 18012 37868
rect 17960 37825 17969 37859
rect 17969 37825 18003 37859
rect 18003 37825 18012 37859
rect 17960 37816 18012 37825
rect 18052 37859 18104 37868
rect 18052 37825 18061 37859
rect 18061 37825 18095 37859
rect 18095 37825 18104 37859
rect 18052 37816 18104 37825
rect 19432 37884 19484 37936
rect 20260 37884 20312 37936
rect 25412 37952 25464 38004
rect 25228 37884 25280 37936
rect 30380 37952 30432 38004
rect 33600 37952 33652 38004
rect 34336 37952 34388 38004
rect 36084 37952 36136 38004
rect 36176 37952 36228 38004
rect 36268 37952 36320 38004
rect 19892 37859 19944 37868
rect 19892 37825 19901 37859
rect 19901 37825 19935 37859
rect 19935 37825 19944 37859
rect 19892 37816 19944 37825
rect 20168 37816 20220 37868
rect 20720 37816 20772 37868
rect 21088 37748 21140 37800
rect 22560 37859 22612 37868
rect 22560 37825 22569 37859
rect 22569 37825 22603 37859
rect 22603 37825 22612 37859
rect 22560 37816 22612 37825
rect 22744 37859 22796 37868
rect 22744 37825 22753 37859
rect 22753 37825 22787 37859
rect 22787 37825 22796 37859
rect 22744 37816 22796 37825
rect 23388 37859 23440 37868
rect 23388 37825 23397 37859
rect 23397 37825 23431 37859
rect 23431 37825 23440 37859
rect 23388 37816 23440 37825
rect 23480 37816 23532 37868
rect 24492 37816 24544 37868
rect 22376 37791 22428 37800
rect 22376 37757 22385 37791
rect 22385 37757 22419 37791
rect 22419 37757 22428 37791
rect 22376 37748 22428 37757
rect 22468 37791 22520 37800
rect 22468 37757 22477 37791
rect 22477 37757 22511 37791
rect 22511 37757 22520 37791
rect 22468 37748 22520 37757
rect 12256 37612 12308 37664
rect 12992 37612 13044 37664
rect 14372 37612 14424 37664
rect 16304 37655 16356 37664
rect 16304 37621 16313 37655
rect 16313 37621 16347 37655
rect 16347 37621 16356 37655
rect 16304 37612 16356 37621
rect 16764 37612 16816 37664
rect 21272 37612 21324 37664
rect 22192 37680 22244 37732
rect 24768 37791 24820 37800
rect 24768 37757 24777 37791
rect 24777 37757 24811 37791
rect 24811 37757 24820 37791
rect 24768 37748 24820 37757
rect 25136 37816 25188 37868
rect 25872 37859 25924 37868
rect 25872 37825 25881 37859
rect 25881 37825 25915 37859
rect 25915 37825 25924 37859
rect 25872 37816 25924 37825
rect 26700 37816 26752 37868
rect 27068 37816 27120 37868
rect 27528 37816 27580 37868
rect 28080 37816 28132 37868
rect 28632 37816 28684 37868
rect 25780 37748 25832 37800
rect 26240 37748 26292 37800
rect 25872 37680 25924 37732
rect 30196 37859 30248 37868
rect 30196 37825 30205 37859
rect 30205 37825 30239 37859
rect 30239 37825 30248 37859
rect 30196 37816 30248 37825
rect 30380 37859 30432 37868
rect 30380 37825 30389 37859
rect 30389 37825 30423 37859
rect 30423 37825 30432 37859
rect 30380 37816 30432 37825
rect 31668 37884 31720 37936
rect 32312 37859 32364 37868
rect 32312 37825 32321 37859
rect 32321 37825 32355 37859
rect 32355 37825 32364 37859
rect 32312 37816 32364 37825
rect 34428 37884 34480 37936
rect 33784 37859 33836 37868
rect 33784 37825 33793 37859
rect 33793 37825 33827 37859
rect 33827 37825 33836 37859
rect 33784 37816 33836 37825
rect 33968 37816 34020 37868
rect 29460 37791 29512 37800
rect 29460 37757 29469 37791
rect 29469 37757 29503 37791
rect 29503 37757 29512 37791
rect 29460 37748 29512 37757
rect 30012 37748 30064 37800
rect 33600 37748 33652 37800
rect 34428 37680 34480 37732
rect 24492 37612 24544 37664
rect 25228 37612 25280 37664
rect 25688 37655 25740 37664
rect 25688 37621 25697 37655
rect 25697 37621 25731 37655
rect 25731 37621 25740 37655
rect 25688 37612 25740 37621
rect 26148 37655 26200 37664
rect 26148 37621 26157 37655
rect 26157 37621 26191 37655
rect 26191 37621 26200 37655
rect 26148 37612 26200 37621
rect 27712 37612 27764 37664
rect 28632 37612 28684 37664
rect 28724 37655 28776 37664
rect 28724 37621 28733 37655
rect 28733 37621 28767 37655
rect 28767 37621 28776 37655
rect 28724 37612 28776 37621
rect 29552 37655 29604 37664
rect 29552 37621 29561 37655
rect 29561 37621 29595 37655
rect 29595 37621 29604 37655
rect 29552 37612 29604 37621
rect 30288 37612 30340 37664
rect 32036 37612 32088 37664
rect 32404 37612 32456 37664
rect 35072 37816 35124 37868
rect 35900 37859 35952 37868
rect 35900 37825 35910 37859
rect 35910 37825 35944 37859
rect 35944 37825 35952 37859
rect 35900 37816 35952 37825
rect 35992 37748 36044 37800
rect 36452 37816 36504 37868
rect 36728 37816 36780 37868
rect 37280 37816 37332 37868
rect 38292 37748 38344 37800
rect 36360 37680 36412 37732
rect 39304 37816 39356 37868
rect 40960 37927 41012 37936
rect 40960 37893 40969 37927
rect 40969 37893 41003 37927
rect 41003 37893 41012 37927
rect 40960 37884 41012 37893
rect 42708 37952 42760 38004
rect 43076 37884 43128 37936
rect 39120 37680 39172 37732
rect 39212 37612 39264 37664
rect 40408 37748 40460 37800
rect 41144 37816 41196 37868
rect 42984 37816 43036 37868
rect 43996 37748 44048 37800
rect 39672 37612 39724 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 4896 37451 4948 37460
rect 4896 37417 4905 37451
rect 4905 37417 4939 37451
rect 4939 37417 4948 37451
rect 4896 37408 4948 37417
rect 11704 37408 11756 37460
rect 11980 37408 12032 37460
rect 13268 37408 13320 37460
rect 14096 37408 14148 37460
rect 14740 37408 14792 37460
rect 20444 37451 20496 37460
rect 20444 37417 20453 37451
rect 20453 37417 20487 37451
rect 20487 37417 20496 37451
rect 20444 37408 20496 37417
rect 22376 37408 22428 37460
rect 26056 37408 26108 37460
rect 27620 37408 27672 37460
rect 11152 37340 11204 37392
rect 11520 37383 11572 37392
rect 11520 37349 11529 37383
rect 11529 37349 11563 37383
rect 11563 37349 11572 37383
rect 11520 37340 11572 37349
rect 12716 37340 12768 37392
rect 13360 37340 13412 37392
rect 22468 37340 22520 37392
rect 24768 37340 24820 37392
rect 25596 37383 25648 37392
rect 25596 37349 25605 37383
rect 25605 37349 25639 37383
rect 25639 37349 25648 37383
rect 25596 37340 25648 37349
rect 5356 37272 5408 37324
rect 6184 37272 6236 37324
rect 7932 37272 7984 37324
rect 12256 37272 12308 37324
rect 13084 37272 13136 37324
rect 13728 37272 13780 37324
rect 15936 37272 15988 37324
rect 17132 37315 17184 37324
rect 17132 37281 17141 37315
rect 17141 37281 17175 37315
rect 17175 37281 17184 37315
rect 17132 37272 17184 37281
rect 5540 37136 5592 37188
rect 7012 37204 7064 37256
rect 6920 37136 6972 37188
rect 8208 37247 8260 37256
rect 8208 37213 8217 37247
rect 8217 37213 8251 37247
rect 8251 37213 8260 37247
rect 8208 37204 8260 37213
rect 9680 37204 9732 37256
rect 10048 37247 10100 37256
rect 10048 37213 10057 37247
rect 10057 37213 10091 37247
rect 10091 37213 10100 37247
rect 10048 37204 10100 37213
rect 10324 37247 10376 37256
rect 10324 37213 10333 37247
rect 10333 37213 10367 37247
rect 10367 37213 10376 37247
rect 10324 37204 10376 37213
rect 11612 37204 11664 37256
rect 7840 37136 7892 37188
rect 8116 37136 8168 37188
rect 11336 37136 11388 37188
rect 11888 37204 11940 37256
rect 12164 37204 12216 37256
rect 14464 37247 14516 37256
rect 14464 37213 14473 37247
rect 14473 37213 14507 37247
rect 14507 37213 14516 37247
rect 14464 37204 14516 37213
rect 16764 37247 16816 37256
rect 16764 37213 16773 37247
rect 16773 37213 16807 37247
rect 16807 37213 16816 37247
rect 16764 37204 16816 37213
rect 17684 37204 17736 37256
rect 12532 37136 12584 37188
rect 14188 37136 14240 37188
rect 15568 37136 15620 37188
rect 17040 37179 17092 37188
rect 17040 37145 17049 37179
rect 17049 37145 17083 37179
rect 17083 37145 17092 37179
rect 17040 37136 17092 37145
rect 6828 37068 6880 37120
rect 7380 37111 7432 37120
rect 7380 37077 7389 37111
rect 7389 37077 7423 37111
rect 7423 37077 7432 37111
rect 7380 37068 7432 37077
rect 10692 37068 10744 37120
rect 11796 37068 11848 37120
rect 15752 37068 15804 37120
rect 25688 37272 25740 37324
rect 26516 37272 26568 37324
rect 27620 37272 27672 37324
rect 28448 37272 28500 37324
rect 20536 37136 20588 37188
rect 23388 37204 23440 37256
rect 21364 37136 21416 37188
rect 24952 37247 25004 37256
rect 24952 37213 24961 37247
rect 24961 37213 24995 37247
rect 24995 37213 25004 37247
rect 24952 37204 25004 37213
rect 25504 37204 25556 37256
rect 25780 37247 25832 37256
rect 25780 37213 25789 37247
rect 25789 37213 25823 37247
rect 25823 37213 25832 37247
rect 25780 37204 25832 37213
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 27160 37204 27212 37256
rect 25228 37136 25280 37188
rect 20904 37111 20956 37120
rect 20904 37077 20913 37111
rect 20913 37077 20947 37111
rect 20947 37077 20956 37111
rect 20904 37068 20956 37077
rect 25044 37068 25096 37120
rect 26700 37111 26752 37120
rect 26700 37077 26709 37111
rect 26709 37077 26743 37111
rect 26743 37077 26752 37111
rect 26700 37068 26752 37077
rect 27436 37179 27488 37188
rect 27436 37145 27445 37179
rect 27445 37145 27479 37179
rect 27479 37145 27488 37179
rect 27436 37136 27488 37145
rect 27620 37179 27672 37188
rect 27620 37145 27629 37179
rect 27629 37145 27663 37179
rect 27663 37145 27672 37179
rect 27620 37136 27672 37145
rect 27896 37204 27948 37256
rect 29092 37247 29144 37256
rect 29092 37213 29101 37247
rect 29101 37213 29135 37247
rect 29135 37213 29144 37247
rect 29092 37204 29144 37213
rect 30196 37204 30248 37256
rect 31852 37272 31904 37324
rect 36452 37408 36504 37460
rect 37188 37408 37240 37460
rect 37464 37408 37516 37460
rect 33324 37340 33376 37392
rect 35808 37383 35860 37392
rect 35808 37349 35817 37383
rect 35817 37349 35851 37383
rect 35851 37349 35860 37383
rect 39304 37408 39356 37460
rect 39488 37451 39540 37460
rect 39488 37417 39497 37451
rect 39497 37417 39531 37451
rect 39531 37417 39540 37451
rect 39488 37408 39540 37417
rect 35808 37340 35860 37349
rect 37648 37340 37700 37392
rect 40500 37340 40552 37392
rect 41420 37340 41472 37392
rect 35440 37272 35492 37324
rect 32036 37204 32088 37256
rect 32496 37204 32548 37256
rect 32680 37247 32732 37256
rect 32680 37213 32689 37247
rect 32689 37213 32723 37247
rect 32723 37213 32732 37247
rect 32680 37204 32732 37213
rect 28724 37068 28776 37120
rect 28816 37068 28868 37120
rect 31484 37179 31536 37188
rect 31484 37145 31493 37179
rect 31493 37145 31527 37179
rect 31527 37145 31536 37179
rect 31484 37136 31536 37145
rect 31576 37136 31628 37188
rect 32772 37068 32824 37120
rect 33876 37247 33928 37256
rect 33876 37213 33885 37247
rect 33885 37213 33919 37247
rect 33919 37213 33928 37247
rect 33876 37204 33928 37213
rect 33968 37247 34020 37256
rect 33968 37213 33977 37247
rect 33977 37213 34011 37247
rect 34011 37213 34020 37247
rect 33968 37204 34020 37213
rect 34244 37204 34296 37256
rect 35716 37247 35768 37256
rect 35716 37213 35725 37247
rect 35725 37213 35759 37247
rect 35759 37213 35768 37247
rect 35716 37204 35768 37213
rect 38292 37272 38344 37324
rect 38660 37272 38712 37324
rect 35532 37136 35584 37188
rect 37188 37204 37240 37256
rect 36636 37068 36688 37120
rect 36912 37179 36964 37188
rect 36912 37145 36921 37179
rect 36921 37145 36955 37179
rect 36955 37145 36964 37179
rect 36912 37136 36964 37145
rect 37280 37136 37332 37188
rect 39120 37179 39172 37188
rect 39120 37145 39129 37179
rect 39129 37145 39163 37179
rect 39163 37145 39172 37179
rect 39120 37136 39172 37145
rect 39396 37204 39448 37256
rect 39488 37204 39540 37256
rect 39856 37136 39908 37188
rect 40500 37247 40552 37256
rect 40500 37213 40509 37247
rect 40509 37213 40543 37247
rect 40543 37213 40552 37247
rect 40500 37204 40552 37213
rect 41144 37204 41196 37256
rect 41788 37204 41840 37256
rect 40408 37179 40460 37188
rect 40408 37145 40417 37179
rect 40417 37145 40451 37179
rect 40451 37145 40460 37179
rect 40408 37136 40460 37145
rect 42616 37136 42668 37188
rect 42984 37068 43036 37120
rect 43076 37111 43128 37120
rect 43076 37077 43085 37111
rect 43085 37077 43119 37111
rect 43119 37077 43128 37111
rect 43076 37068 43128 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 8116 36864 8168 36916
rect 9956 36864 10008 36916
rect 12348 36864 12400 36916
rect 14004 36864 14056 36916
rect 7840 36771 7892 36780
rect 7840 36737 7849 36771
rect 7849 36737 7883 36771
rect 7883 36737 7892 36771
rect 7840 36728 7892 36737
rect 8024 36771 8076 36780
rect 8024 36737 8033 36771
rect 8033 36737 8067 36771
rect 8067 36737 8076 36771
rect 8024 36728 8076 36737
rect 8944 36771 8996 36780
rect 8944 36737 8953 36771
rect 8953 36737 8987 36771
rect 8987 36737 8996 36771
rect 8944 36728 8996 36737
rect 10692 36796 10744 36848
rect 15016 36864 15068 36916
rect 17132 36907 17184 36916
rect 17132 36873 17141 36907
rect 17141 36873 17175 36907
rect 17175 36873 17184 36907
rect 17132 36864 17184 36873
rect 20628 36864 20680 36916
rect 24584 36864 24636 36916
rect 9680 36728 9732 36780
rect 10232 36728 10284 36780
rect 10416 36728 10468 36780
rect 8208 36660 8260 36712
rect 10048 36703 10100 36712
rect 10048 36669 10057 36703
rect 10057 36669 10091 36703
rect 10091 36669 10100 36703
rect 10048 36660 10100 36669
rect 10508 36660 10560 36712
rect 11428 36728 11480 36780
rect 16488 36796 16540 36848
rect 16580 36796 16632 36848
rect 17868 36796 17920 36848
rect 22008 36796 22060 36848
rect 12624 36728 12676 36780
rect 13084 36728 13136 36780
rect 13636 36728 13688 36780
rect 14648 36771 14700 36780
rect 14648 36737 14662 36771
rect 14662 36737 14696 36771
rect 14696 36737 14700 36771
rect 14648 36728 14700 36737
rect 15476 36771 15528 36780
rect 15476 36737 15485 36771
rect 15485 36737 15519 36771
rect 15519 36737 15528 36771
rect 15476 36728 15528 36737
rect 15568 36771 15620 36780
rect 15568 36737 15577 36771
rect 15577 36737 15611 36771
rect 15611 36737 15620 36771
rect 15568 36728 15620 36737
rect 16856 36771 16908 36780
rect 16856 36737 16865 36771
rect 16865 36737 16899 36771
rect 16899 36737 16908 36771
rect 16856 36728 16908 36737
rect 17040 36728 17092 36780
rect 8852 36592 8904 36644
rect 9772 36592 9824 36644
rect 11428 36592 11480 36644
rect 6736 36567 6788 36576
rect 6736 36533 6745 36567
rect 6745 36533 6779 36567
rect 6779 36533 6788 36567
rect 6736 36524 6788 36533
rect 7288 36524 7340 36576
rect 7564 36524 7616 36576
rect 10876 36524 10928 36576
rect 10968 36524 11020 36576
rect 14740 36703 14792 36712
rect 14740 36669 14749 36703
rect 14749 36669 14783 36703
rect 14783 36669 14792 36703
rect 14740 36660 14792 36669
rect 12992 36524 13044 36576
rect 14556 36524 14608 36576
rect 15752 36592 15804 36644
rect 15844 36592 15896 36644
rect 19156 36771 19208 36780
rect 19156 36737 19165 36771
rect 19165 36737 19199 36771
rect 19199 36737 19208 36771
rect 19156 36728 19208 36737
rect 17776 36660 17828 36712
rect 22100 36771 22152 36780
rect 22100 36737 22109 36771
rect 22109 36737 22143 36771
rect 22143 36737 22152 36771
rect 22100 36728 22152 36737
rect 22284 36771 22336 36780
rect 22284 36737 22293 36771
rect 22293 36737 22327 36771
rect 22327 36737 22336 36771
rect 22284 36728 22336 36737
rect 25872 36796 25924 36848
rect 27528 36796 27580 36848
rect 19432 36703 19484 36712
rect 19432 36669 19441 36703
rect 19441 36669 19475 36703
rect 19475 36669 19484 36703
rect 19432 36660 19484 36669
rect 20536 36703 20588 36712
rect 20536 36669 20545 36703
rect 20545 36669 20579 36703
rect 20579 36669 20588 36703
rect 20536 36660 20588 36669
rect 20812 36660 20864 36712
rect 24860 36771 24912 36780
rect 24860 36737 24869 36771
rect 24869 36737 24903 36771
rect 24903 36737 24912 36771
rect 24860 36728 24912 36737
rect 25044 36771 25096 36780
rect 25044 36737 25053 36771
rect 25053 36737 25087 36771
rect 25087 36737 25096 36771
rect 25044 36728 25096 36737
rect 27344 36771 27396 36780
rect 27344 36737 27353 36771
rect 27353 36737 27387 36771
rect 27387 36737 27396 36771
rect 27344 36728 27396 36737
rect 33140 36864 33192 36916
rect 34428 36864 34480 36916
rect 30380 36796 30432 36848
rect 27160 36660 27212 36712
rect 27528 36660 27580 36712
rect 18880 36592 18932 36644
rect 15016 36567 15068 36576
rect 15016 36533 15025 36567
rect 15025 36533 15059 36567
rect 15059 36533 15068 36567
rect 15016 36524 15068 36533
rect 15108 36524 15160 36576
rect 15568 36524 15620 36576
rect 16396 36524 16448 36576
rect 24860 36592 24912 36644
rect 22468 36567 22520 36576
rect 22468 36533 22477 36567
rect 22477 36533 22511 36567
rect 22511 36533 22520 36567
rect 22468 36524 22520 36533
rect 23664 36524 23716 36576
rect 25596 36524 25648 36576
rect 25964 36524 26016 36576
rect 28816 36660 28868 36712
rect 31024 36771 31076 36780
rect 31024 36737 31033 36771
rect 31033 36737 31067 36771
rect 31067 36737 31076 36771
rect 31024 36728 31076 36737
rect 29920 36703 29972 36712
rect 29920 36669 29929 36703
rect 29929 36669 29963 36703
rect 29963 36669 29972 36703
rect 29920 36660 29972 36669
rect 30748 36703 30800 36712
rect 30748 36669 30757 36703
rect 30757 36669 30791 36703
rect 30791 36669 30800 36703
rect 30748 36660 30800 36669
rect 31668 36728 31720 36780
rect 32588 36771 32640 36780
rect 32588 36737 32597 36771
rect 32597 36737 32631 36771
rect 32631 36737 32640 36771
rect 32588 36728 32640 36737
rect 33048 36796 33100 36848
rect 33416 36728 33468 36780
rect 33600 36728 33652 36780
rect 34060 36728 34112 36780
rect 34796 36796 34848 36848
rect 36636 36864 36688 36916
rect 39120 36864 39172 36916
rect 39948 36864 40000 36916
rect 42616 36907 42668 36916
rect 42616 36873 42625 36907
rect 42625 36873 42659 36907
rect 42659 36873 42668 36907
rect 42616 36864 42668 36873
rect 42984 36864 43036 36916
rect 27712 36567 27764 36576
rect 27712 36533 27721 36567
rect 27721 36533 27755 36567
rect 27755 36533 27764 36567
rect 27712 36524 27764 36533
rect 27988 36524 28040 36576
rect 28080 36524 28132 36576
rect 34244 36660 34296 36712
rect 34796 36703 34848 36712
rect 34796 36669 34805 36703
rect 34805 36669 34839 36703
rect 34839 36669 34848 36703
rect 34796 36660 34848 36669
rect 41604 36728 41656 36780
rect 43076 36728 43128 36780
rect 36820 36660 36872 36712
rect 43168 36703 43220 36712
rect 43168 36669 43177 36703
rect 43177 36669 43211 36703
rect 43211 36669 43220 36703
rect 43168 36660 43220 36669
rect 31484 36524 31536 36576
rect 33416 36592 33468 36644
rect 37832 36524 37884 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 6736 36320 6788 36372
rect 9956 36320 10008 36372
rect 11520 36320 11572 36372
rect 11704 36320 11756 36372
rect 13636 36363 13688 36372
rect 13636 36329 13645 36363
rect 13645 36329 13679 36363
rect 13679 36329 13688 36363
rect 13636 36320 13688 36329
rect 14556 36363 14608 36372
rect 14556 36329 14565 36363
rect 14565 36329 14599 36363
rect 14599 36329 14608 36363
rect 14556 36320 14608 36329
rect 15844 36320 15896 36372
rect 16028 36363 16080 36372
rect 16028 36329 16037 36363
rect 16037 36329 16071 36363
rect 16071 36329 16080 36363
rect 16028 36320 16080 36329
rect 17132 36363 17184 36372
rect 17132 36329 17141 36363
rect 17141 36329 17175 36363
rect 17175 36329 17184 36363
rect 17132 36320 17184 36329
rect 17684 36320 17736 36372
rect 17776 36363 17828 36372
rect 17776 36329 17785 36363
rect 17785 36329 17819 36363
rect 17819 36329 17828 36363
rect 17776 36320 17828 36329
rect 17868 36320 17920 36372
rect 19064 36320 19116 36372
rect 19892 36320 19944 36372
rect 20352 36320 20404 36372
rect 20536 36320 20588 36372
rect 22468 36320 22520 36372
rect 23756 36320 23808 36372
rect 8024 36252 8076 36304
rect 10232 36252 10284 36304
rect 10508 36252 10560 36304
rect 11060 36252 11112 36304
rect 12808 36252 12860 36304
rect 15568 36252 15620 36304
rect 15660 36295 15712 36304
rect 15660 36261 15669 36295
rect 15669 36261 15703 36295
rect 15703 36261 15712 36295
rect 15660 36252 15712 36261
rect 15936 36252 15988 36304
rect 4620 36116 4672 36168
rect 4988 36048 5040 36100
rect 6828 36159 6880 36168
rect 6828 36125 6837 36159
rect 6837 36125 6871 36159
rect 6871 36125 6880 36159
rect 6828 36116 6880 36125
rect 6920 36159 6972 36168
rect 6920 36125 6929 36159
rect 6929 36125 6963 36159
rect 6963 36125 6972 36159
rect 6920 36116 6972 36125
rect 7196 36159 7248 36168
rect 7196 36125 7205 36159
rect 7205 36125 7239 36159
rect 7239 36125 7248 36159
rect 7196 36116 7248 36125
rect 8116 36116 8168 36168
rect 9772 36116 9824 36168
rect 7564 36048 7616 36100
rect 8852 36048 8904 36100
rect 5540 35980 5592 36032
rect 6644 36023 6696 36032
rect 6644 35989 6653 36023
rect 6653 35989 6687 36023
rect 6687 35989 6696 36023
rect 6644 35980 6696 35989
rect 8300 35980 8352 36032
rect 8576 35980 8628 36032
rect 10324 36159 10376 36168
rect 10324 36125 10333 36159
rect 10333 36125 10367 36159
rect 10367 36125 10376 36159
rect 10324 36116 10376 36125
rect 11060 36159 11112 36168
rect 11060 36125 11069 36159
rect 11069 36125 11103 36159
rect 11103 36125 11112 36159
rect 11060 36116 11112 36125
rect 11336 36159 11388 36168
rect 11336 36125 11345 36159
rect 11345 36125 11379 36159
rect 11379 36125 11388 36159
rect 11336 36116 11388 36125
rect 11520 36159 11572 36168
rect 11520 36125 11529 36159
rect 11529 36125 11563 36159
rect 11563 36125 11572 36159
rect 11520 36116 11572 36125
rect 11888 36116 11940 36168
rect 12532 36159 12584 36168
rect 12532 36125 12541 36159
rect 12541 36125 12575 36159
rect 12575 36125 12584 36159
rect 12532 36116 12584 36125
rect 12900 36116 12952 36168
rect 13084 36116 13136 36168
rect 14648 36184 14700 36236
rect 17316 36227 17368 36236
rect 17316 36193 17325 36227
rect 17325 36193 17359 36227
rect 17359 36193 17368 36227
rect 17316 36184 17368 36193
rect 14188 36116 14240 36168
rect 11980 36048 12032 36100
rect 15108 36116 15160 36168
rect 16948 36116 17000 36168
rect 17684 36116 17736 36168
rect 15016 36048 15068 36100
rect 22100 36252 22152 36304
rect 23388 36252 23440 36304
rect 17960 36159 18012 36168
rect 17960 36125 17969 36159
rect 17969 36125 18003 36159
rect 18003 36125 18012 36159
rect 17960 36116 18012 36125
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 19064 36116 19116 36168
rect 19432 36159 19484 36168
rect 19432 36125 19441 36159
rect 19441 36125 19475 36159
rect 19475 36125 19484 36159
rect 19432 36116 19484 36125
rect 10508 35980 10560 36032
rect 11244 36023 11296 36032
rect 11244 35989 11253 36023
rect 11253 35989 11287 36023
rect 11287 35989 11296 36023
rect 11244 35980 11296 35989
rect 11520 35980 11572 36032
rect 12716 35980 12768 36032
rect 17132 35980 17184 36032
rect 19892 36116 19944 36168
rect 20812 36159 20864 36168
rect 20812 36125 20821 36159
rect 20821 36125 20855 36159
rect 20855 36125 20864 36159
rect 20812 36116 20864 36125
rect 21088 36159 21140 36168
rect 21088 36125 21097 36159
rect 21097 36125 21131 36159
rect 21131 36125 21140 36159
rect 21088 36116 21140 36125
rect 21272 36159 21324 36168
rect 21272 36125 21281 36159
rect 21281 36125 21315 36159
rect 21315 36125 21324 36159
rect 21272 36116 21324 36125
rect 22100 36116 22152 36168
rect 22468 36116 22520 36168
rect 24492 36184 24544 36236
rect 23664 36159 23716 36168
rect 22284 36048 22336 36100
rect 23664 36125 23673 36159
rect 23673 36125 23707 36159
rect 23707 36125 23716 36159
rect 23664 36116 23716 36125
rect 24952 36252 25004 36304
rect 27528 36363 27580 36372
rect 27528 36329 27537 36363
rect 27537 36329 27571 36363
rect 27571 36329 27580 36363
rect 27528 36320 27580 36329
rect 28632 36363 28684 36372
rect 28632 36329 28641 36363
rect 28641 36329 28675 36363
rect 28675 36329 28684 36363
rect 28632 36320 28684 36329
rect 30012 36363 30064 36372
rect 30012 36329 30021 36363
rect 30021 36329 30055 36363
rect 30055 36329 30064 36363
rect 30012 36320 30064 36329
rect 30288 36363 30340 36372
rect 30288 36329 30316 36363
rect 30316 36329 30340 36363
rect 30288 36320 30340 36329
rect 37372 36363 37424 36372
rect 37372 36329 37381 36363
rect 37381 36329 37415 36363
rect 37415 36329 37424 36363
rect 37372 36320 37424 36329
rect 29368 36252 29420 36304
rect 29920 36252 29972 36304
rect 21916 35980 21968 36032
rect 23480 36091 23532 36100
rect 23480 36057 23489 36091
rect 23489 36057 23523 36091
rect 23523 36057 23532 36091
rect 23480 36048 23532 36057
rect 26884 36184 26936 36236
rect 27160 36184 27212 36236
rect 27896 36227 27948 36236
rect 27896 36193 27905 36227
rect 27905 36193 27939 36227
rect 27939 36193 27948 36227
rect 27896 36184 27948 36193
rect 28080 36184 28132 36236
rect 32680 36252 32732 36304
rect 33232 36295 33284 36304
rect 33232 36261 33241 36295
rect 33241 36261 33275 36295
rect 33275 36261 33284 36295
rect 33232 36252 33284 36261
rect 35716 36252 35768 36304
rect 31024 36184 31076 36236
rect 31944 36184 31996 36236
rect 25044 36159 25096 36168
rect 25044 36125 25053 36159
rect 25053 36125 25087 36159
rect 25087 36125 25096 36159
rect 25044 36116 25096 36125
rect 26516 36116 26568 36168
rect 27712 36159 27764 36168
rect 27712 36125 27721 36159
rect 27721 36125 27755 36159
rect 27755 36125 27764 36159
rect 27712 36116 27764 36125
rect 25136 35980 25188 36032
rect 25412 35980 25464 36032
rect 27436 35980 27488 36032
rect 27620 36048 27672 36100
rect 28448 36116 28500 36168
rect 27896 36048 27948 36100
rect 28816 36116 28868 36168
rect 28908 36159 28960 36168
rect 28908 36125 28917 36159
rect 28917 36125 28951 36159
rect 28951 36125 28960 36159
rect 28908 36116 28960 36125
rect 30288 36116 30340 36168
rect 30380 36116 30432 36168
rect 30564 36116 30616 36168
rect 31668 36116 31720 36168
rect 32128 36116 32180 36168
rect 32588 36116 32640 36168
rect 32956 36159 33008 36168
rect 32956 36125 32965 36159
rect 32965 36125 32999 36159
rect 32999 36125 33008 36159
rect 32956 36116 33008 36125
rect 33140 36116 33192 36168
rect 34060 36159 34112 36168
rect 34060 36125 34069 36159
rect 34069 36125 34103 36159
rect 34103 36125 34112 36159
rect 34060 36116 34112 36125
rect 34796 36184 34848 36236
rect 36176 36184 36228 36236
rect 35072 36159 35124 36168
rect 35072 36125 35081 36159
rect 35081 36125 35115 36159
rect 35115 36125 35124 36159
rect 35072 36116 35124 36125
rect 30748 36048 30800 36100
rect 29184 36023 29236 36032
rect 29184 35989 29193 36023
rect 29193 35989 29227 36023
rect 29227 35989 29236 36023
rect 29184 35980 29236 35989
rect 32772 35980 32824 36032
rect 33324 36048 33376 36100
rect 33416 36048 33468 36100
rect 33692 35980 33744 36032
rect 34520 35980 34572 36032
rect 36084 36116 36136 36168
rect 36636 36116 36688 36168
rect 36912 36159 36964 36168
rect 36912 36125 36919 36159
rect 36919 36125 36964 36159
rect 36912 36116 36964 36125
rect 36360 36048 36412 36100
rect 37004 36091 37056 36100
rect 37004 36057 37013 36091
rect 37013 36057 37047 36091
rect 37047 36057 37056 36091
rect 37004 36048 37056 36057
rect 35992 35980 36044 36032
rect 36452 35980 36504 36032
rect 38016 36116 38068 36168
rect 38752 36159 38804 36168
rect 38752 36125 38761 36159
rect 38761 36125 38795 36159
rect 38795 36125 38804 36159
rect 38752 36116 38804 36125
rect 39764 36184 39816 36236
rect 37924 36023 37976 36032
rect 37924 35989 37933 36023
rect 37933 35989 37967 36023
rect 37967 35989 37976 36023
rect 37924 35980 37976 35989
rect 38016 35980 38068 36032
rect 39396 36048 39448 36100
rect 41880 36159 41932 36168
rect 41880 36125 41889 36159
rect 41889 36125 41923 36159
rect 41923 36125 41932 36159
rect 41880 36116 41932 36125
rect 39120 35980 39172 36032
rect 39304 35980 39356 36032
rect 39948 35980 40000 36032
rect 42616 36048 42668 36100
rect 40960 35980 41012 36032
rect 43260 36023 43312 36032
rect 43260 35989 43269 36023
rect 43269 35989 43303 36023
rect 43303 35989 43312 36023
rect 43260 35980 43312 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4988 35819 5040 35828
rect 4988 35785 4997 35819
rect 4997 35785 5031 35819
rect 5031 35785 5040 35819
rect 4988 35776 5040 35785
rect 6828 35776 6880 35828
rect 7196 35708 7248 35760
rect 8208 35776 8260 35828
rect 8944 35776 8996 35828
rect 9772 35776 9824 35828
rect 10324 35776 10376 35828
rect 11980 35776 12032 35828
rect 10048 35708 10100 35760
rect 11888 35751 11940 35760
rect 11888 35717 11897 35751
rect 11897 35717 11931 35751
rect 11931 35717 11940 35751
rect 11888 35708 11940 35717
rect 5172 35615 5224 35624
rect 5172 35581 5181 35615
rect 5181 35581 5215 35615
rect 5215 35581 5224 35615
rect 5172 35572 5224 35581
rect 5356 35615 5408 35624
rect 5356 35581 5365 35615
rect 5365 35581 5399 35615
rect 5399 35581 5408 35615
rect 5356 35572 5408 35581
rect 5448 35615 5500 35624
rect 5448 35581 5457 35615
rect 5457 35581 5491 35615
rect 5491 35581 5500 35615
rect 5448 35572 5500 35581
rect 7840 35640 7892 35692
rect 8760 35640 8812 35692
rect 8852 35640 8904 35692
rect 9220 35683 9272 35692
rect 9220 35649 9229 35683
rect 9229 35649 9263 35683
rect 9263 35649 9272 35683
rect 9220 35640 9272 35649
rect 9680 35683 9732 35692
rect 9680 35649 9689 35683
rect 9689 35649 9723 35683
rect 9723 35649 9732 35683
rect 9680 35640 9732 35649
rect 9956 35640 10008 35692
rect 10140 35683 10192 35692
rect 10140 35649 10149 35683
rect 10149 35649 10183 35683
rect 10183 35649 10192 35683
rect 10140 35640 10192 35649
rect 10600 35640 10652 35692
rect 11612 35640 11664 35692
rect 12808 35819 12860 35828
rect 12808 35785 12817 35819
rect 12817 35785 12851 35819
rect 12851 35785 12860 35819
rect 12808 35776 12860 35785
rect 13360 35776 13412 35828
rect 15200 35776 15252 35828
rect 16028 35776 16080 35828
rect 12716 35708 12768 35760
rect 13544 35708 13596 35760
rect 14464 35708 14516 35760
rect 12992 35640 13044 35692
rect 14556 35683 14608 35692
rect 14556 35649 14565 35683
rect 14565 35649 14599 35683
rect 14599 35649 14608 35683
rect 14556 35640 14608 35649
rect 14832 35640 14884 35692
rect 14372 35615 14424 35624
rect 14372 35581 14381 35615
rect 14381 35581 14415 35615
rect 14415 35581 14424 35615
rect 14372 35572 14424 35581
rect 15384 35683 15436 35692
rect 15384 35649 15393 35683
rect 15393 35649 15427 35683
rect 15427 35649 15436 35683
rect 15384 35640 15436 35649
rect 15752 35640 15804 35692
rect 17040 35708 17092 35760
rect 16948 35683 17000 35692
rect 16948 35649 16957 35683
rect 16957 35649 16991 35683
rect 16991 35649 17000 35683
rect 16948 35640 17000 35649
rect 17132 35683 17184 35692
rect 17132 35649 17141 35683
rect 17141 35649 17175 35683
rect 17175 35649 17184 35683
rect 17132 35640 17184 35649
rect 19340 35776 19392 35828
rect 19892 35776 19944 35828
rect 20076 35776 20128 35828
rect 20720 35776 20772 35828
rect 21088 35776 21140 35828
rect 23480 35819 23532 35828
rect 23480 35785 23489 35819
rect 23489 35785 23523 35819
rect 23523 35785 23532 35819
rect 23480 35776 23532 35785
rect 23848 35776 23900 35828
rect 24584 35776 24636 35828
rect 18144 35708 18196 35760
rect 17868 35683 17920 35692
rect 17868 35649 17877 35683
rect 17877 35649 17911 35683
rect 17911 35649 17920 35683
rect 17868 35640 17920 35649
rect 18052 35683 18104 35692
rect 18052 35649 18061 35683
rect 18061 35649 18095 35683
rect 18095 35649 18104 35683
rect 18052 35640 18104 35649
rect 18880 35683 18932 35692
rect 18880 35649 18889 35683
rect 18889 35649 18923 35683
rect 18923 35649 18932 35683
rect 18880 35640 18932 35649
rect 21272 35640 21324 35692
rect 7012 35504 7064 35556
rect 8392 35504 8444 35556
rect 9680 35504 9732 35556
rect 10968 35504 11020 35556
rect 12716 35504 12768 35556
rect 15660 35572 15712 35624
rect 21916 35572 21968 35624
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 22560 35640 22612 35692
rect 23296 35640 23348 35692
rect 25044 35708 25096 35760
rect 25136 35708 25188 35760
rect 24032 35640 24084 35692
rect 24216 35683 24268 35692
rect 24216 35649 24225 35683
rect 24225 35649 24259 35683
rect 24259 35649 24268 35683
rect 24216 35640 24268 35649
rect 25688 35640 25740 35692
rect 27068 35640 27120 35692
rect 22192 35504 22244 35556
rect 22468 35615 22520 35624
rect 22468 35581 22477 35615
rect 22477 35581 22511 35615
rect 22511 35581 22520 35615
rect 22468 35572 22520 35581
rect 23388 35504 23440 35556
rect 25136 35615 25188 35624
rect 25136 35581 25145 35615
rect 25145 35581 25179 35615
rect 25179 35581 25188 35615
rect 25136 35572 25188 35581
rect 26332 35572 26384 35624
rect 27620 35776 27672 35828
rect 27712 35776 27764 35828
rect 31944 35776 31996 35828
rect 33048 35776 33100 35828
rect 36912 35776 36964 35828
rect 38752 35776 38804 35828
rect 42616 35819 42668 35828
rect 42616 35785 42625 35819
rect 42625 35785 42659 35819
rect 42659 35785 42668 35819
rect 42616 35776 42668 35785
rect 28356 35708 28408 35760
rect 28908 35708 28960 35760
rect 30380 35708 30432 35760
rect 27712 35640 27764 35692
rect 27896 35640 27948 35692
rect 30104 35683 30156 35692
rect 30104 35649 30113 35683
rect 30113 35649 30147 35683
rect 30147 35649 30156 35683
rect 30104 35640 30156 35649
rect 30564 35640 30616 35692
rect 28356 35572 28408 35624
rect 7104 35479 7156 35488
rect 7104 35445 7113 35479
rect 7113 35445 7147 35479
rect 7147 35445 7156 35479
rect 7104 35436 7156 35445
rect 8116 35436 8168 35488
rect 14280 35479 14332 35488
rect 14280 35445 14289 35479
rect 14289 35445 14323 35479
rect 14323 35445 14332 35479
rect 14280 35436 14332 35445
rect 18236 35479 18288 35488
rect 18236 35445 18245 35479
rect 18245 35445 18279 35479
rect 18279 35445 18288 35479
rect 18236 35436 18288 35445
rect 20444 35479 20496 35488
rect 20444 35445 20453 35479
rect 20453 35445 20487 35479
rect 20487 35445 20496 35479
rect 20444 35436 20496 35445
rect 22560 35436 22612 35488
rect 24216 35436 24268 35488
rect 24768 35436 24820 35488
rect 25412 35504 25464 35556
rect 26148 35436 26200 35488
rect 26608 35479 26660 35488
rect 26608 35445 26617 35479
rect 26617 35445 26651 35479
rect 26651 35445 26660 35479
rect 26608 35436 26660 35445
rect 27988 35504 28040 35556
rect 30380 35615 30432 35624
rect 30380 35581 30389 35615
rect 30389 35581 30423 35615
rect 30423 35581 30432 35615
rect 30380 35572 30432 35581
rect 30840 35572 30892 35624
rect 30932 35504 30984 35556
rect 31484 35640 31536 35692
rect 32680 35708 32732 35760
rect 36176 35708 36228 35760
rect 37924 35751 37976 35760
rect 37924 35717 37933 35751
rect 37933 35717 37967 35751
rect 37967 35717 37976 35751
rect 37924 35708 37976 35717
rect 38016 35708 38068 35760
rect 33324 35640 33376 35692
rect 33416 35683 33468 35692
rect 33416 35649 33425 35683
rect 33425 35649 33459 35683
rect 33459 35649 33468 35683
rect 33416 35640 33468 35649
rect 34244 35640 34296 35692
rect 34336 35683 34388 35692
rect 34336 35649 34345 35683
rect 34345 35649 34379 35683
rect 34379 35649 34388 35683
rect 34336 35640 34388 35649
rect 38384 35640 38436 35692
rect 31208 35615 31260 35624
rect 31208 35581 31217 35615
rect 31217 35581 31251 35615
rect 31251 35581 31260 35615
rect 31208 35572 31260 35581
rect 31760 35572 31812 35624
rect 32036 35572 32088 35624
rect 33140 35615 33192 35624
rect 33140 35581 33149 35615
rect 33149 35581 33183 35615
rect 33183 35581 33192 35615
rect 33140 35572 33192 35581
rect 35624 35572 35676 35624
rect 41788 35708 41840 35760
rect 43260 35708 43312 35760
rect 39120 35640 39172 35692
rect 40960 35683 41012 35692
rect 40960 35649 40969 35683
rect 40969 35649 41003 35683
rect 41003 35649 41012 35683
rect 40960 35640 41012 35649
rect 29000 35436 29052 35488
rect 29644 35436 29696 35488
rect 36912 35504 36964 35556
rect 41236 35683 41288 35692
rect 41236 35649 41245 35683
rect 41245 35649 41279 35683
rect 41279 35649 41288 35683
rect 41236 35640 41288 35649
rect 41328 35683 41380 35692
rect 41328 35649 41337 35683
rect 41337 35649 41371 35683
rect 41371 35649 41380 35683
rect 41328 35640 41380 35649
rect 32128 35436 32180 35488
rect 33600 35436 33652 35488
rect 38108 35479 38160 35488
rect 38108 35445 38117 35479
rect 38117 35445 38151 35479
rect 38151 35445 38160 35479
rect 38108 35436 38160 35445
rect 40316 35436 40368 35488
rect 41144 35504 41196 35556
rect 41972 35572 42024 35624
rect 43260 35615 43312 35624
rect 43260 35581 43269 35615
rect 43269 35581 43303 35615
rect 43303 35581 43312 35615
rect 43260 35572 43312 35581
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5448 35232 5500 35284
rect 9588 35232 9640 35284
rect 5172 35164 5224 35216
rect 7564 35139 7616 35148
rect 7564 35105 7573 35139
rect 7573 35105 7607 35139
rect 7607 35105 7616 35139
rect 7564 35096 7616 35105
rect 5540 35071 5592 35080
rect 5540 35037 5549 35071
rect 5549 35037 5583 35071
rect 5583 35037 5592 35071
rect 5540 35028 5592 35037
rect 5632 35071 5684 35080
rect 5632 35037 5641 35071
rect 5641 35037 5675 35071
rect 5675 35037 5684 35071
rect 5632 35028 5684 35037
rect 7288 35071 7340 35080
rect 7288 35037 7297 35071
rect 7297 35037 7331 35071
rect 7331 35037 7340 35071
rect 7288 35028 7340 35037
rect 7656 35071 7708 35080
rect 7656 35037 7665 35071
rect 7665 35037 7699 35071
rect 7699 35037 7708 35071
rect 7656 35028 7708 35037
rect 7932 35096 7984 35148
rect 7932 34960 7984 35012
rect 7564 34892 7616 34944
rect 8760 35164 8812 35216
rect 11704 35164 11756 35216
rect 12256 35232 12308 35284
rect 12624 35232 12676 35284
rect 15660 35275 15712 35284
rect 15660 35241 15669 35275
rect 15669 35241 15703 35275
rect 15703 35241 15712 35275
rect 15660 35232 15712 35241
rect 17868 35232 17920 35284
rect 20444 35232 20496 35284
rect 22284 35275 22336 35284
rect 22284 35241 22293 35275
rect 22293 35241 22327 35275
rect 22327 35241 22336 35275
rect 22284 35232 22336 35241
rect 25136 35275 25188 35284
rect 25136 35241 25145 35275
rect 25145 35241 25179 35275
rect 25179 35241 25188 35275
rect 25136 35232 25188 35241
rect 27068 35275 27120 35284
rect 27068 35241 27077 35275
rect 27077 35241 27111 35275
rect 27111 35241 27120 35275
rect 27068 35232 27120 35241
rect 27804 35232 27856 35284
rect 27896 35275 27948 35284
rect 27896 35241 27905 35275
rect 27905 35241 27939 35275
rect 27939 35241 27948 35275
rect 27896 35232 27948 35241
rect 29552 35232 29604 35284
rect 9496 35071 9548 35080
rect 9496 35037 9505 35071
rect 9505 35037 9539 35071
rect 9539 35037 9548 35071
rect 9496 35028 9548 35037
rect 10232 35028 10284 35080
rect 10784 35071 10836 35080
rect 10784 35037 10793 35071
rect 10793 35037 10827 35071
rect 10827 35037 10836 35071
rect 10784 35028 10836 35037
rect 11704 35028 11756 35080
rect 11796 35028 11848 35080
rect 12532 35071 12584 35080
rect 12532 35037 12541 35071
rect 12541 35037 12575 35071
rect 12575 35037 12584 35071
rect 12532 35028 12584 35037
rect 14372 35139 14424 35148
rect 14372 35105 14381 35139
rect 14381 35105 14415 35139
rect 14415 35105 14424 35139
rect 14372 35096 14424 35105
rect 14464 35028 14516 35080
rect 14556 35071 14608 35080
rect 14556 35037 14565 35071
rect 14565 35037 14599 35071
rect 14599 35037 14608 35071
rect 14556 35028 14608 35037
rect 19892 35164 19944 35216
rect 22100 35164 22152 35216
rect 22560 35164 22612 35216
rect 23296 35096 23348 35148
rect 23388 35096 23440 35148
rect 27988 35164 28040 35216
rect 31208 35232 31260 35284
rect 27068 35096 27120 35148
rect 8484 34960 8536 35012
rect 9772 34960 9824 35012
rect 15476 35003 15528 35012
rect 15476 34969 15485 35003
rect 15485 34969 15519 35003
rect 15519 34969 15528 35003
rect 15476 34960 15528 34969
rect 17224 35003 17276 35012
rect 17224 34969 17233 35003
rect 17233 34969 17267 35003
rect 17267 34969 17276 35003
rect 17224 34960 17276 34969
rect 17500 34960 17552 35012
rect 11060 34935 11112 34944
rect 11060 34901 11069 34935
rect 11069 34901 11103 34935
rect 11103 34901 11112 34935
rect 11060 34892 11112 34901
rect 11336 34892 11388 34944
rect 15384 34892 15436 34944
rect 22468 35071 22520 35080
rect 22468 35037 22477 35071
rect 22477 35037 22511 35071
rect 22511 35037 22520 35071
rect 22468 35028 22520 35037
rect 23020 35028 23072 35080
rect 23112 35003 23164 35012
rect 23112 34969 23121 35003
rect 23121 34969 23155 35003
rect 23155 34969 23164 35003
rect 23112 34960 23164 34969
rect 23204 34960 23256 35012
rect 23940 35028 23992 35080
rect 25780 35028 25832 35080
rect 26148 35071 26200 35080
rect 26148 35037 26157 35071
rect 26157 35037 26191 35071
rect 26191 35037 26200 35071
rect 26148 35028 26200 35037
rect 26240 35071 26292 35080
rect 26240 35037 26249 35071
rect 26249 35037 26283 35071
rect 26283 35037 26292 35071
rect 26240 35028 26292 35037
rect 27528 35028 27580 35080
rect 27620 35028 27672 35080
rect 28540 35096 28592 35148
rect 30840 35207 30892 35216
rect 30840 35173 30849 35207
rect 30849 35173 30883 35207
rect 30883 35173 30892 35207
rect 30840 35164 30892 35173
rect 30932 35207 30984 35216
rect 30932 35173 30941 35207
rect 30941 35173 30975 35207
rect 30975 35173 30984 35207
rect 32588 35232 32640 35284
rect 34888 35232 34940 35284
rect 35808 35232 35860 35284
rect 38016 35232 38068 35284
rect 30932 35164 30984 35173
rect 31392 35164 31444 35216
rect 32128 35096 32180 35148
rect 32772 35139 32824 35148
rect 32772 35105 32781 35139
rect 32781 35105 32815 35139
rect 32815 35105 32824 35139
rect 32772 35096 32824 35105
rect 32956 35096 33008 35148
rect 36084 35164 36136 35216
rect 28448 35028 28500 35080
rect 28816 35071 28868 35080
rect 28816 35037 28825 35071
rect 28825 35037 28859 35071
rect 28859 35037 28868 35071
rect 28816 35028 28868 35037
rect 24860 34960 24912 35012
rect 25044 34960 25096 35012
rect 25872 34960 25924 35012
rect 27068 34960 27120 35012
rect 29460 35028 29512 35080
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 31392 35028 31444 35080
rect 32036 35028 32088 35080
rect 25412 34892 25464 34944
rect 27620 34892 27672 34944
rect 28908 34892 28960 34944
rect 29552 34960 29604 35012
rect 30380 34892 30432 34944
rect 30472 34935 30524 34944
rect 30472 34901 30481 34935
rect 30481 34901 30515 34935
rect 30515 34901 30524 34935
rect 30472 34892 30524 34901
rect 30656 34892 30708 34944
rect 33416 35028 33468 35080
rect 33968 35028 34020 35080
rect 36728 35096 36780 35148
rect 38108 35164 38160 35216
rect 35808 35071 35860 35080
rect 35808 35037 35817 35071
rect 35817 35037 35851 35071
rect 35851 35037 35860 35071
rect 35808 35028 35860 35037
rect 35900 35071 35952 35080
rect 35900 35037 35910 35071
rect 35910 35037 35944 35071
rect 35944 35037 35952 35071
rect 35900 35028 35952 35037
rect 35716 34960 35768 35012
rect 36084 35003 36136 35012
rect 36084 34969 36093 35003
rect 36093 34969 36127 35003
rect 36127 34969 36136 35003
rect 36084 34960 36136 34969
rect 36176 35003 36228 35012
rect 36176 34969 36185 35003
rect 36185 34969 36219 35003
rect 36219 34969 36228 35003
rect 36176 34960 36228 34969
rect 33048 34892 33100 34944
rect 34244 34935 34296 34944
rect 34244 34901 34253 34935
rect 34253 34901 34287 34935
rect 34287 34901 34296 34935
rect 34244 34892 34296 34901
rect 35348 34892 35400 34944
rect 36452 35028 36504 35080
rect 36912 35071 36964 35080
rect 36912 35037 36921 35071
rect 36921 35037 36955 35071
rect 36955 35037 36964 35071
rect 36912 35028 36964 35037
rect 37740 35096 37792 35148
rect 37372 35028 37424 35080
rect 37832 35028 37884 35080
rect 38384 35028 38436 35080
rect 37280 35003 37332 35012
rect 37280 34969 37289 35003
rect 37289 34969 37323 35003
rect 37323 34969 37332 35003
rect 37280 34960 37332 34969
rect 40040 35139 40092 35148
rect 40040 35105 40049 35139
rect 40049 35105 40083 35139
rect 40083 35105 40092 35139
rect 40040 35096 40092 35105
rect 43996 35096 44048 35148
rect 41420 35028 41472 35080
rect 41880 35028 41932 35080
rect 41972 35071 42024 35080
rect 41972 35037 41981 35071
rect 41981 35037 42015 35071
rect 42015 35037 42024 35071
rect 41972 35028 42024 35037
rect 42892 35071 42944 35080
rect 42892 35037 42901 35071
rect 42901 35037 42935 35071
rect 42935 35037 42944 35071
rect 42892 35028 42944 35037
rect 40592 34960 40644 35012
rect 41236 34960 41288 35012
rect 43996 34960 44048 35012
rect 40776 34892 40828 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 8944 34688 8996 34740
rect 9404 34688 9456 34740
rect 9864 34688 9916 34740
rect 4620 34620 4672 34672
rect 7564 34663 7616 34672
rect 7564 34629 7573 34663
rect 7573 34629 7607 34663
rect 7607 34629 7616 34663
rect 7564 34620 7616 34629
rect 5816 34552 5868 34604
rect 7104 34595 7156 34604
rect 7104 34561 7113 34595
rect 7113 34561 7147 34595
rect 7147 34561 7156 34595
rect 7104 34552 7156 34561
rect 7288 34595 7340 34604
rect 7288 34561 7297 34595
rect 7297 34561 7331 34595
rect 7331 34561 7340 34595
rect 7288 34552 7340 34561
rect 8484 34595 8536 34604
rect 8484 34561 8493 34595
rect 8493 34561 8527 34595
rect 8527 34561 8536 34595
rect 8484 34552 8536 34561
rect 9680 34620 9732 34672
rect 10600 34620 10652 34672
rect 9404 34595 9456 34604
rect 9404 34561 9413 34595
rect 9413 34561 9447 34595
rect 9447 34561 9456 34595
rect 9404 34552 9456 34561
rect 10048 34595 10100 34604
rect 10048 34561 10057 34595
rect 10057 34561 10091 34595
rect 10091 34561 10100 34595
rect 10048 34552 10100 34561
rect 8392 34527 8444 34536
rect 8392 34493 8401 34527
rect 8401 34493 8435 34527
rect 8435 34493 8444 34527
rect 8392 34484 8444 34493
rect 7564 34416 7616 34468
rect 8852 34484 8904 34536
rect 9220 34484 9272 34536
rect 11704 34595 11756 34604
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 12440 34620 12492 34672
rect 13084 34663 13136 34672
rect 13084 34629 13093 34663
rect 13093 34629 13127 34663
rect 13127 34629 13136 34663
rect 13084 34620 13136 34629
rect 13728 34620 13780 34672
rect 12716 34595 12768 34604
rect 10324 34484 10376 34536
rect 12716 34561 12725 34595
rect 12725 34561 12759 34595
rect 12759 34561 12768 34595
rect 12716 34552 12768 34561
rect 13544 34595 13596 34604
rect 13544 34561 13553 34595
rect 13553 34561 13587 34595
rect 13587 34561 13596 34595
rect 13544 34552 13596 34561
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 17960 34688 18012 34740
rect 22744 34688 22796 34740
rect 24584 34688 24636 34740
rect 28172 34688 28224 34740
rect 28448 34688 28500 34740
rect 31300 34688 31352 34740
rect 31484 34688 31536 34740
rect 32588 34688 32640 34740
rect 33048 34731 33100 34740
rect 33048 34697 33057 34731
rect 33057 34697 33091 34731
rect 33091 34697 33100 34731
rect 33048 34688 33100 34697
rect 33140 34688 33192 34740
rect 34428 34688 34480 34740
rect 35808 34688 35860 34740
rect 36728 34688 36780 34740
rect 38476 34688 38528 34740
rect 14464 34484 14516 34536
rect 10232 34416 10284 34468
rect 6368 34348 6420 34400
rect 6920 34391 6972 34400
rect 6920 34357 6929 34391
rect 6929 34357 6963 34391
rect 6963 34357 6972 34391
rect 6920 34348 6972 34357
rect 7472 34391 7524 34400
rect 7472 34357 7481 34391
rect 7481 34357 7515 34391
rect 7515 34357 7524 34391
rect 7472 34348 7524 34357
rect 9680 34348 9732 34400
rect 12900 34416 12952 34468
rect 13544 34416 13596 34468
rect 17040 34620 17092 34672
rect 18236 34620 18288 34672
rect 24860 34663 24912 34672
rect 17224 34552 17276 34604
rect 15476 34484 15528 34536
rect 19524 34552 19576 34604
rect 19156 34484 19208 34536
rect 24860 34629 24869 34663
rect 24869 34629 24903 34663
rect 24903 34629 24912 34663
rect 24860 34620 24912 34629
rect 25780 34663 25832 34672
rect 25780 34629 25789 34663
rect 25789 34629 25823 34663
rect 25823 34629 25832 34663
rect 25780 34620 25832 34629
rect 22468 34552 22520 34604
rect 23388 34552 23440 34604
rect 23940 34552 23992 34604
rect 24308 34552 24360 34604
rect 25320 34552 25372 34604
rect 27160 34620 27212 34672
rect 26332 34552 26384 34604
rect 28080 34620 28132 34672
rect 28632 34620 28684 34672
rect 25044 34484 25096 34536
rect 25872 34484 25924 34536
rect 28356 34595 28408 34604
rect 28356 34561 28365 34595
rect 28365 34561 28399 34595
rect 28399 34561 28408 34595
rect 28908 34620 28960 34672
rect 29184 34620 29236 34672
rect 35900 34620 35952 34672
rect 40316 34620 40368 34672
rect 28356 34552 28408 34561
rect 23112 34416 23164 34468
rect 24768 34416 24820 34468
rect 27712 34484 27764 34536
rect 27804 34484 27856 34536
rect 29460 34484 29512 34536
rect 31300 34595 31352 34604
rect 31300 34561 31309 34595
rect 31309 34561 31343 34595
rect 31343 34561 31352 34595
rect 31300 34552 31352 34561
rect 33232 34595 33284 34604
rect 33232 34561 33241 34595
rect 33241 34561 33275 34595
rect 33275 34561 33284 34595
rect 33232 34552 33284 34561
rect 33692 34595 33744 34604
rect 33692 34561 33701 34595
rect 33701 34561 33735 34595
rect 33735 34561 33744 34595
rect 33692 34552 33744 34561
rect 34428 34552 34480 34604
rect 35992 34552 36044 34604
rect 31392 34484 31444 34536
rect 32496 34484 32548 34536
rect 34888 34527 34940 34536
rect 34888 34493 34897 34527
rect 34897 34493 34931 34527
rect 34931 34493 34940 34527
rect 34888 34484 34940 34493
rect 36360 34595 36412 34604
rect 36360 34561 36369 34595
rect 36369 34561 36403 34595
rect 36403 34561 36412 34595
rect 36360 34552 36412 34561
rect 36452 34595 36504 34604
rect 36452 34561 36497 34595
rect 36497 34561 36504 34595
rect 36452 34552 36504 34561
rect 36636 34595 36688 34604
rect 36636 34561 36645 34595
rect 36645 34561 36679 34595
rect 36679 34561 36688 34595
rect 36636 34552 36688 34561
rect 14280 34348 14332 34400
rect 25412 34348 25464 34400
rect 26976 34416 27028 34468
rect 29092 34416 29144 34468
rect 29644 34416 29696 34468
rect 34152 34416 34204 34468
rect 34244 34416 34296 34468
rect 28448 34348 28500 34400
rect 29000 34348 29052 34400
rect 30012 34391 30064 34400
rect 30012 34357 30021 34391
rect 30021 34357 30055 34391
rect 30055 34357 30064 34391
rect 30012 34348 30064 34357
rect 32864 34348 32916 34400
rect 33048 34348 33100 34400
rect 33600 34391 33652 34400
rect 33600 34357 33609 34391
rect 33609 34357 33643 34391
rect 33643 34357 33652 34391
rect 33600 34348 33652 34357
rect 35808 34348 35860 34400
rect 36176 34416 36228 34468
rect 38200 34484 38252 34536
rect 43260 34348 43312 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5816 34187 5868 34196
rect 5816 34153 5825 34187
rect 5825 34153 5859 34187
rect 5859 34153 5868 34187
rect 5816 34144 5868 34153
rect 7472 34144 7524 34196
rect 8116 34144 8168 34196
rect 7104 34076 7156 34128
rect 10784 34076 10836 34128
rect 6644 34008 6696 34060
rect 6368 33940 6420 33992
rect 6460 33983 6512 33992
rect 6460 33949 6469 33983
rect 6469 33949 6503 33983
rect 6503 33949 6512 33983
rect 6460 33940 6512 33949
rect 7012 33940 7064 33992
rect 8484 34008 8536 34060
rect 8576 34008 8628 34060
rect 10232 34051 10284 34060
rect 10232 34017 10241 34051
rect 10241 34017 10275 34051
rect 10275 34017 10284 34051
rect 10232 34008 10284 34017
rect 10324 34051 10376 34060
rect 10324 34017 10333 34051
rect 10333 34017 10367 34051
rect 10367 34017 10376 34051
rect 10324 34008 10376 34017
rect 10968 34008 11020 34060
rect 11152 34076 11204 34128
rect 11428 34076 11480 34128
rect 12164 34076 12216 34128
rect 6736 33872 6788 33924
rect 7840 33872 7892 33924
rect 7932 33872 7984 33924
rect 9404 33940 9456 33992
rect 9680 33872 9732 33924
rect 7012 33847 7064 33856
rect 7012 33813 7021 33847
rect 7021 33813 7055 33847
rect 7055 33813 7064 33847
rect 7012 33804 7064 33813
rect 9864 33847 9916 33856
rect 9864 33813 9873 33847
rect 9873 33813 9907 33847
rect 9907 33813 9916 33847
rect 9864 33804 9916 33813
rect 11060 33915 11112 33924
rect 11060 33881 11077 33915
rect 11077 33881 11112 33915
rect 11060 33872 11112 33881
rect 11152 33915 11204 33924
rect 11152 33881 11161 33915
rect 11161 33881 11195 33915
rect 11195 33881 11204 33915
rect 11152 33872 11204 33881
rect 12164 33915 12216 33924
rect 12164 33881 12173 33915
rect 12173 33881 12207 33915
rect 12207 33881 12216 33915
rect 12164 33872 12216 33881
rect 12900 33915 12952 33924
rect 12900 33881 12909 33915
rect 12909 33881 12943 33915
rect 12943 33881 12952 33915
rect 12900 33872 12952 33881
rect 13820 33940 13872 33992
rect 16948 33940 17000 33992
rect 26792 34144 26844 34196
rect 28264 34144 28316 34196
rect 28448 34144 28500 34196
rect 23020 34076 23072 34128
rect 25872 34076 25924 34128
rect 27988 34076 28040 34128
rect 30196 34076 30248 34128
rect 31668 34144 31720 34196
rect 32772 34144 32824 34196
rect 33784 34187 33836 34196
rect 33784 34153 33793 34187
rect 33793 34153 33827 34187
rect 33827 34153 33836 34187
rect 33784 34144 33836 34153
rect 31024 34076 31076 34128
rect 20352 34008 20404 34060
rect 14280 33872 14332 33924
rect 17408 33872 17460 33924
rect 17500 33915 17552 33924
rect 17500 33881 17509 33915
rect 17509 33881 17543 33915
rect 17543 33881 17552 33915
rect 17500 33872 17552 33881
rect 19524 33983 19576 33992
rect 19524 33949 19533 33983
rect 19533 33949 19567 33983
rect 19567 33949 19576 33983
rect 19524 33940 19576 33949
rect 20260 33940 20312 33992
rect 23112 34008 23164 34060
rect 19248 33872 19300 33924
rect 23020 33983 23072 33992
rect 23020 33949 23029 33983
rect 23029 33949 23063 33983
rect 23063 33949 23072 33983
rect 23020 33940 23072 33949
rect 25504 34008 25556 34060
rect 11336 33804 11388 33856
rect 15108 33804 15160 33856
rect 17868 33804 17920 33856
rect 22928 33872 22980 33924
rect 24860 33940 24912 33992
rect 26240 33940 26292 33992
rect 26884 33940 26936 33992
rect 27160 33940 27212 33992
rect 27528 33983 27580 33992
rect 27528 33949 27537 33983
rect 27537 33949 27571 33983
rect 27571 33949 27580 33983
rect 27528 33940 27580 33949
rect 29000 34008 29052 34060
rect 29276 34008 29328 34060
rect 23848 33872 23900 33924
rect 25964 33872 26016 33924
rect 26056 33872 26108 33924
rect 28080 33940 28132 33992
rect 29920 33983 29972 33992
rect 29920 33949 29929 33983
rect 29929 33949 29963 33983
rect 29963 33949 29972 33983
rect 29920 33940 29972 33949
rect 30564 33983 30616 33992
rect 30564 33949 30573 33983
rect 30573 33949 30607 33983
rect 30607 33949 30616 33983
rect 30564 33940 30616 33949
rect 30840 33983 30892 33992
rect 30840 33949 30849 33983
rect 30849 33949 30883 33983
rect 30883 33949 30892 33983
rect 30840 33940 30892 33949
rect 31760 33940 31812 33992
rect 33692 34008 33744 34060
rect 34520 34076 34572 34128
rect 35992 34144 36044 34196
rect 36636 34144 36688 34196
rect 19984 33804 20036 33856
rect 22284 33804 22336 33856
rect 22468 33847 22520 33856
rect 22468 33813 22477 33847
rect 22477 33813 22511 33847
rect 22511 33813 22520 33847
rect 22468 33804 22520 33813
rect 26884 33847 26936 33856
rect 26884 33813 26893 33847
rect 26893 33813 26927 33847
rect 26927 33813 26936 33847
rect 26884 33804 26936 33813
rect 27528 33804 27580 33856
rect 27896 33804 27948 33856
rect 30104 33804 30156 33856
rect 30564 33804 30616 33856
rect 31484 33872 31536 33924
rect 32404 33872 32456 33924
rect 33968 33983 34020 33992
rect 33968 33949 33977 33983
rect 33977 33949 34011 33983
rect 34011 33949 34020 33983
rect 33968 33940 34020 33949
rect 35440 34008 35492 34060
rect 41788 34008 41840 34060
rect 34152 33940 34204 33992
rect 34428 33872 34480 33924
rect 31392 33804 31444 33856
rect 31944 33847 31996 33856
rect 31944 33813 31971 33847
rect 31971 33813 31996 33847
rect 31944 33804 31996 33813
rect 33600 33804 33652 33856
rect 34520 33804 34572 33856
rect 35256 33915 35308 33924
rect 35256 33881 35265 33915
rect 35265 33881 35299 33915
rect 35299 33881 35308 33915
rect 35256 33872 35308 33881
rect 35716 33983 35768 33992
rect 35716 33949 35725 33983
rect 35725 33949 35759 33983
rect 35759 33949 35768 33983
rect 35716 33940 35768 33949
rect 37556 33872 37608 33924
rect 42616 33872 42668 33924
rect 35716 33804 35768 33856
rect 35808 33804 35860 33856
rect 42984 33804 43036 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 8116 33600 8168 33652
rect 10232 33600 10284 33652
rect 20168 33600 20220 33652
rect 25964 33600 26016 33652
rect 26424 33600 26476 33652
rect 6368 33532 6420 33584
rect 6276 33464 6328 33516
rect 6828 33507 6880 33516
rect 6828 33473 6837 33507
rect 6837 33473 6871 33507
rect 6871 33473 6880 33507
rect 6828 33464 6880 33473
rect 7012 33464 7064 33516
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 6644 33439 6696 33448
rect 6644 33405 6653 33439
rect 6653 33405 6687 33439
rect 6687 33405 6696 33439
rect 6644 33396 6696 33405
rect 9496 33532 9548 33584
rect 10692 33532 10744 33584
rect 9312 33507 9364 33516
rect 9312 33473 9321 33507
rect 9321 33473 9355 33507
rect 9355 33473 9364 33507
rect 9772 33507 9824 33516
rect 9312 33464 9364 33473
rect 9772 33473 9781 33507
rect 9781 33473 9815 33507
rect 9815 33473 9824 33507
rect 9772 33464 9824 33473
rect 10416 33464 10468 33516
rect 10784 33464 10836 33516
rect 10968 33464 11020 33516
rect 12072 33575 12124 33584
rect 12072 33541 12081 33575
rect 12081 33541 12115 33575
rect 12115 33541 12124 33575
rect 12072 33532 12124 33541
rect 12900 33575 12952 33584
rect 12900 33541 12909 33575
rect 12909 33541 12943 33575
rect 12943 33541 12952 33575
rect 12900 33532 12952 33541
rect 17500 33532 17552 33584
rect 19984 33532 20036 33584
rect 13544 33507 13596 33516
rect 13544 33473 13553 33507
rect 13553 33473 13587 33507
rect 13587 33473 13596 33507
rect 13544 33464 13596 33473
rect 14188 33464 14240 33516
rect 7564 33328 7616 33380
rect 7932 33328 7984 33380
rect 4896 33303 4948 33312
rect 4896 33269 4905 33303
rect 4905 33269 4939 33303
rect 4939 33269 4948 33303
rect 4896 33260 4948 33269
rect 5264 33303 5316 33312
rect 5264 33269 5273 33303
rect 5273 33269 5307 33303
rect 5307 33269 5316 33303
rect 5264 33260 5316 33269
rect 8760 33303 8812 33312
rect 8760 33269 8769 33303
rect 8769 33269 8803 33303
rect 8803 33269 8812 33303
rect 8760 33260 8812 33269
rect 8852 33260 8904 33312
rect 13360 33396 13412 33448
rect 13728 33396 13780 33448
rect 14556 33464 14608 33516
rect 16948 33464 17000 33516
rect 17132 33507 17184 33516
rect 17132 33473 17166 33507
rect 17166 33473 17184 33507
rect 17132 33464 17184 33473
rect 23848 33532 23900 33584
rect 25504 33532 25556 33584
rect 26792 33532 26844 33584
rect 26884 33532 26936 33584
rect 28448 33600 28500 33652
rect 30656 33600 30708 33652
rect 31116 33600 31168 33652
rect 31760 33643 31812 33652
rect 31760 33609 31769 33643
rect 31769 33609 31803 33643
rect 31803 33609 31812 33643
rect 31760 33600 31812 33609
rect 32956 33600 33008 33652
rect 36452 33600 36504 33652
rect 37096 33600 37148 33652
rect 32496 33532 32548 33584
rect 33048 33532 33100 33584
rect 34796 33532 34848 33584
rect 35532 33532 35584 33584
rect 36176 33532 36228 33584
rect 19248 33396 19300 33448
rect 16488 33328 16540 33380
rect 20628 33328 20680 33380
rect 22284 33464 22336 33516
rect 24308 33507 24360 33516
rect 24308 33473 24317 33507
rect 24317 33473 24351 33507
rect 24351 33473 24360 33507
rect 24308 33464 24360 33473
rect 24860 33464 24912 33516
rect 25412 33507 25464 33516
rect 25412 33473 25421 33507
rect 25421 33473 25455 33507
rect 25455 33473 25464 33507
rect 25412 33464 25464 33473
rect 22468 33439 22520 33448
rect 22468 33405 22477 33439
rect 22477 33405 22511 33439
rect 22511 33405 22520 33439
rect 22468 33396 22520 33405
rect 23664 33396 23716 33448
rect 26608 33464 26660 33516
rect 27252 33464 27304 33516
rect 28540 33464 28592 33516
rect 28908 33507 28960 33516
rect 28908 33473 28917 33507
rect 28917 33473 28951 33507
rect 28951 33473 28960 33507
rect 28908 33464 28960 33473
rect 27528 33396 27580 33448
rect 27620 33439 27672 33448
rect 27620 33405 27629 33439
rect 27629 33405 27663 33439
rect 27663 33405 27672 33439
rect 27620 33396 27672 33405
rect 22376 33328 22428 33380
rect 28816 33396 28868 33448
rect 30564 33464 30616 33516
rect 30748 33464 30800 33516
rect 31208 33464 31260 33516
rect 31300 33507 31352 33516
rect 31300 33473 31309 33507
rect 31309 33473 31343 33507
rect 31343 33473 31352 33507
rect 31300 33464 31352 33473
rect 31392 33507 31444 33516
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 31576 33464 31628 33516
rect 30196 33439 30248 33448
rect 30196 33405 30205 33439
rect 30205 33405 30239 33439
rect 30239 33405 30248 33439
rect 30196 33396 30248 33405
rect 37740 33464 37792 33516
rect 39304 33575 39356 33584
rect 39304 33541 39313 33575
rect 39313 33541 39347 33575
rect 39347 33541 39356 33575
rect 39304 33532 39356 33541
rect 42616 33643 42668 33652
rect 42616 33609 42625 33643
rect 42625 33609 42659 33643
rect 42659 33609 42668 33643
rect 42616 33600 42668 33609
rect 40316 33532 40368 33584
rect 42984 33575 43036 33584
rect 33416 33396 33468 33448
rect 36728 33439 36780 33448
rect 36728 33405 36737 33439
rect 36737 33405 36771 33439
rect 36771 33405 36780 33439
rect 36728 33396 36780 33405
rect 38660 33396 38712 33448
rect 39396 33396 39448 33448
rect 28448 33371 28500 33380
rect 28448 33337 28457 33371
rect 28457 33337 28491 33371
rect 28491 33337 28500 33371
rect 28448 33328 28500 33337
rect 9772 33303 9824 33312
rect 9772 33269 9781 33303
rect 9781 33269 9815 33303
rect 9815 33269 9824 33303
rect 9772 33260 9824 33269
rect 12992 33260 13044 33312
rect 13544 33303 13596 33312
rect 13544 33269 13553 33303
rect 13553 33269 13587 33303
rect 13587 33269 13596 33303
rect 13544 33260 13596 33269
rect 13912 33260 13964 33312
rect 20076 33260 20128 33312
rect 22284 33260 22336 33312
rect 24860 33260 24912 33312
rect 27160 33260 27212 33312
rect 27804 33303 27856 33312
rect 27804 33269 27813 33303
rect 27813 33269 27847 33303
rect 27847 33269 27856 33303
rect 27804 33260 27856 33269
rect 28080 33260 28132 33312
rect 31668 33328 31720 33380
rect 40592 33464 40644 33516
rect 41144 33464 41196 33516
rect 42984 33541 42993 33575
rect 42993 33541 43027 33575
rect 43027 33541 43036 33575
rect 42984 33532 43036 33541
rect 28632 33303 28684 33312
rect 28632 33269 28641 33303
rect 28641 33269 28675 33303
rect 28675 33269 28684 33303
rect 28632 33260 28684 33269
rect 30748 33260 30800 33312
rect 34428 33303 34480 33312
rect 34428 33269 34437 33303
rect 34437 33269 34471 33303
rect 34471 33269 34480 33303
rect 34428 33260 34480 33269
rect 35348 33303 35400 33312
rect 35348 33269 35357 33303
rect 35357 33269 35391 33303
rect 35391 33269 35400 33303
rect 35348 33260 35400 33269
rect 36452 33260 36504 33312
rect 42892 33328 42944 33380
rect 43260 33439 43312 33448
rect 43260 33405 43269 33439
rect 43269 33405 43303 33439
rect 43303 33405 43312 33439
rect 43260 33396 43312 33405
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 6276 33099 6328 33108
rect 6276 33065 6285 33099
rect 6285 33065 6319 33099
rect 6319 33065 6328 33099
rect 6276 33056 6328 33065
rect 7564 33056 7616 33108
rect 7840 33099 7892 33108
rect 7840 33065 7849 33099
rect 7849 33065 7883 33099
rect 7883 33065 7892 33099
rect 7840 33056 7892 33065
rect 9312 33056 9364 33108
rect 10416 33056 10468 33108
rect 10600 33056 10652 33108
rect 10968 33099 11020 33108
rect 10968 33065 10977 33099
rect 10977 33065 11011 33099
rect 11011 33065 11020 33099
rect 10968 33056 11020 33065
rect 12256 33099 12308 33108
rect 12256 33065 12265 33099
rect 12265 33065 12299 33099
rect 12299 33065 12308 33099
rect 12256 33056 12308 33065
rect 5356 32988 5408 33040
rect 17408 33056 17460 33108
rect 18052 33056 18104 33108
rect 18696 33056 18748 33108
rect 19156 33056 19208 33108
rect 19340 33056 19392 33108
rect 19984 33056 20036 33108
rect 21364 33056 21416 33108
rect 23204 33056 23256 33108
rect 7012 32920 7064 32972
rect 4160 32852 4212 32904
rect 4896 32852 4948 32904
rect 6736 32895 6788 32904
rect 6736 32861 6745 32895
rect 6745 32861 6779 32895
rect 6779 32861 6788 32895
rect 9772 32920 9824 32972
rect 15108 32920 15160 32972
rect 18052 32963 18104 32972
rect 18052 32929 18061 32963
rect 18061 32929 18095 32963
rect 18095 32929 18104 32963
rect 18052 32920 18104 32929
rect 8024 32895 8076 32904
rect 6736 32852 6788 32861
rect 7012 32784 7064 32836
rect 8024 32861 8033 32895
rect 8033 32861 8067 32895
rect 8067 32861 8076 32895
rect 8024 32852 8076 32861
rect 8116 32852 8168 32904
rect 9404 32895 9456 32904
rect 9404 32861 9413 32895
rect 9413 32861 9447 32895
rect 9447 32861 9456 32895
rect 9404 32852 9456 32861
rect 7656 32784 7708 32836
rect 10968 32852 11020 32904
rect 11704 32852 11756 32904
rect 9956 32784 10008 32836
rect 10692 32784 10744 32836
rect 11980 32784 12032 32836
rect 12256 32852 12308 32904
rect 16396 32852 16448 32904
rect 16488 32852 16540 32904
rect 18328 32852 18380 32904
rect 19892 32852 19944 32904
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 21364 32852 21416 32861
rect 23664 32988 23716 33040
rect 22652 32963 22704 32972
rect 22652 32929 22661 32963
rect 22661 32929 22695 32963
rect 22695 32929 22704 32963
rect 22652 32920 22704 32929
rect 24124 32920 24176 32972
rect 24768 32920 24820 32972
rect 25228 33056 25280 33108
rect 26976 32988 27028 33040
rect 27620 33056 27672 33108
rect 28264 33099 28316 33108
rect 28264 33065 28273 33099
rect 28273 33065 28307 33099
rect 28307 33065 28316 33099
rect 28264 33056 28316 33065
rect 28908 33056 28960 33108
rect 35532 32988 35584 33040
rect 37372 32988 37424 33040
rect 22836 32895 22888 32904
rect 22836 32861 22845 32895
rect 22845 32861 22879 32895
rect 22879 32861 22888 32895
rect 22836 32852 22888 32861
rect 15476 32784 15528 32836
rect 17868 32827 17920 32836
rect 17868 32793 17877 32827
rect 17877 32793 17911 32827
rect 17911 32793 17920 32827
rect 17868 32784 17920 32793
rect 7748 32716 7800 32768
rect 8668 32716 8720 32768
rect 10048 32716 10100 32768
rect 10324 32716 10376 32768
rect 11336 32716 11388 32768
rect 12808 32716 12860 32768
rect 14188 32716 14240 32768
rect 19340 32784 19392 32836
rect 18420 32716 18472 32768
rect 20444 32784 20496 32836
rect 22468 32784 22520 32836
rect 23664 32895 23716 32904
rect 23664 32861 23673 32895
rect 23673 32861 23707 32895
rect 23707 32861 23716 32895
rect 23664 32852 23716 32861
rect 24308 32852 24360 32904
rect 26700 32920 26752 32972
rect 26148 32784 26200 32836
rect 26884 32852 26936 32904
rect 29736 32920 29788 32972
rect 30196 32920 30248 32972
rect 29828 32852 29880 32904
rect 30288 32895 30340 32904
rect 30288 32861 30297 32895
rect 30297 32861 30331 32895
rect 30331 32861 30340 32895
rect 30288 32852 30340 32861
rect 30472 32852 30524 32904
rect 30840 32852 30892 32904
rect 33508 32920 33560 32972
rect 33968 32920 34020 32972
rect 35256 32920 35308 32972
rect 35348 32920 35400 32972
rect 38016 32920 38068 32972
rect 33324 32895 33376 32904
rect 33324 32861 33333 32895
rect 33333 32861 33367 32895
rect 33367 32861 33376 32895
rect 33324 32852 33376 32861
rect 33416 32852 33468 32904
rect 34428 32852 34480 32904
rect 35716 32852 35768 32904
rect 35900 32852 35952 32904
rect 36176 32895 36228 32904
rect 36176 32861 36186 32895
rect 36186 32861 36220 32895
rect 36220 32861 36228 32895
rect 36176 32852 36228 32861
rect 37372 32852 37424 32904
rect 37464 32852 37516 32904
rect 28724 32784 28776 32836
rect 28816 32784 28868 32836
rect 32404 32784 32456 32836
rect 34980 32784 35032 32836
rect 19984 32716 20036 32768
rect 21180 32759 21232 32768
rect 21180 32725 21189 32759
rect 21189 32725 21223 32759
rect 21223 32725 21232 32759
rect 21180 32716 21232 32725
rect 23388 32716 23440 32768
rect 24768 32759 24820 32768
rect 24768 32725 24777 32759
rect 24777 32725 24811 32759
rect 24811 32725 24820 32759
rect 24768 32716 24820 32725
rect 26976 32716 27028 32768
rect 29644 32716 29696 32768
rect 34336 32716 34388 32768
rect 36084 32716 36136 32768
rect 36452 32827 36504 32836
rect 36452 32793 36461 32827
rect 36461 32793 36495 32827
rect 36495 32793 36504 32827
rect 36452 32784 36504 32793
rect 38016 32827 38068 32836
rect 38016 32793 38025 32827
rect 38025 32793 38059 32827
rect 38059 32793 38068 32827
rect 38016 32784 38068 32793
rect 38384 32852 38436 32904
rect 37832 32716 37884 32768
rect 38844 32784 38896 32836
rect 38936 32759 38988 32768
rect 38936 32725 38945 32759
rect 38945 32725 38979 32759
rect 38979 32725 38988 32759
rect 38936 32716 38988 32725
rect 41420 32895 41472 32904
rect 41420 32861 41429 32895
rect 41429 32861 41463 32895
rect 41463 32861 41472 32895
rect 41420 32852 41472 32861
rect 41880 32852 41932 32904
rect 42892 32895 42944 32904
rect 42892 32861 42901 32895
rect 42901 32861 42935 32895
rect 42935 32861 42944 32895
rect 42892 32852 42944 32861
rect 39580 32784 39632 32836
rect 43168 32827 43220 32836
rect 43168 32793 43177 32827
rect 43177 32793 43211 32827
rect 43211 32793 43220 32827
rect 43168 32784 43220 32793
rect 39488 32716 39540 32768
rect 40040 32759 40092 32768
rect 40040 32725 40049 32759
rect 40049 32725 40083 32759
rect 40083 32725 40092 32759
rect 40040 32716 40092 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 6644 32512 6696 32564
rect 7748 32555 7800 32564
rect 7748 32521 7757 32555
rect 7757 32521 7791 32555
rect 7791 32521 7800 32555
rect 7748 32512 7800 32521
rect 9404 32512 9456 32564
rect 11336 32512 11388 32564
rect 12716 32512 12768 32564
rect 13360 32512 13412 32564
rect 13636 32512 13688 32564
rect 9312 32444 9364 32496
rect 9588 32487 9640 32496
rect 9588 32453 9597 32487
rect 9597 32453 9631 32487
rect 9631 32453 9640 32487
rect 9588 32444 9640 32453
rect 10784 32444 10836 32496
rect 12440 32444 12492 32496
rect 4712 32376 4764 32428
rect 7288 32419 7340 32428
rect 7288 32385 7297 32419
rect 7297 32385 7331 32419
rect 7331 32385 7340 32419
rect 7288 32376 7340 32385
rect 7656 32376 7708 32428
rect 8576 32419 8628 32428
rect 8576 32385 8585 32419
rect 8585 32385 8619 32419
rect 8619 32385 8628 32419
rect 8576 32376 8628 32385
rect 7012 32308 7064 32360
rect 7564 32308 7616 32360
rect 9496 32376 9548 32428
rect 9680 32376 9732 32428
rect 10784 32308 10836 32360
rect 11704 32308 11756 32360
rect 12072 32308 12124 32360
rect 12808 32419 12860 32428
rect 12808 32385 12817 32419
rect 12817 32385 12851 32419
rect 12851 32385 12860 32419
rect 12808 32376 12860 32385
rect 13084 32419 13136 32428
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 13636 32376 13688 32428
rect 13912 32376 13964 32428
rect 16396 32512 16448 32564
rect 5356 32283 5408 32292
rect 5356 32249 5365 32283
rect 5365 32249 5399 32283
rect 5399 32249 5408 32283
rect 5356 32240 5408 32249
rect 12256 32240 12308 32292
rect 14740 32376 14792 32428
rect 14280 32308 14332 32360
rect 18144 32419 18196 32428
rect 18144 32385 18153 32419
rect 18153 32385 18187 32419
rect 18187 32385 18196 32419
rect 18144 32376 18196 32385
rect 19248 32376 19300 32428
rect 18328 32308 18380 32360
rect 18420 32351 18472 32360
rect 18420 32317 18429 32351
rect 18429 32317 18463 32351
rect 18463 32317 18472 32351
rect 18420 32308 18472 32317
rect 20260 32555 20312 32564
rect 20260 32521 20269 32555
rect 20269 32521 20303 32555
rect 20303 32521 20312 32555
rect 20260 32512 20312 32521
rect 20628 32555 20680 32564
rect 20628 32521 20637 32555
rect 20637 32521 20671 32555
rect 20671 32521 20680 32555
rect 20628 32512 20680 32521
rect 21180 32512 21232 32564
rect 22836 32512 22888 32564
rect 25320 32512 25372 32564
rect 25964 32512 26016 32564
rect 27344 32512 27396 32564
rect 27528 32512 27580 32564
rect 27712 32512 27764 32564
rect 19432 32444 19484 32496
rect 24768 32444 24820 32496
rect 20444 32419 20496 32428
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 22192 32376 22244 32428
rect 22928 32376 22980 32428
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 23020 32308 23072 32360
rect 23664 32376 23716 32428
rect 23848 32419 23900 32428
rect 23848 32385 23857 32419
rect 23857 32385 23891 32419
rect 23891 32385 23900 32419
rect 23848 32376 23900 32385
rect 25228 32376 25280 32428
rect 25780 32444 25832 32496
rect 26056 32376 26108 32428
rect 28264 32444 28316 32496
rect 26516 32419 26568 32428
rect 26516 32385 26525 32419
rect 26525 32385 26559 32419
rect 26559 32385 26568 32419
rect 26516 32376 26568 32385
rect 27528 32376 27580 32428
rect 4160 32172 4212 32224
rect 4620 32172 4672 32224
rect 8024 32172 8076 32224
rect 10324 32172 10376 32224
rect 11612 32172 11664 32224
rect 14556 32172 14608 32224
rect 16212 32215 16264 32224
rect 16212 32181 16221 32215
rect 16221 32181 16255 32215
rect 16255 32181 16264 32215
rect 16212 32172 16264 32181
rect 16304 32172 16356 32224
rect 19984 32172 20036 32224
rect 23112 32172 23164 32224
rect 23480 32172 23532 32224
rect 28448 32376 28500 32428
rect 28264 32308 28316 32360
rect 28816 32444 28868 32496
rect 29092 32376 29144 32428
rect 29828 32512 29880 32564
rect 31576 32444 31628 32496
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 30380 32308 30432 32360
rect 32496 32487 32548 32496
rect 32496 32453 32505 32487
rect 32505 32453 32539 32487
rect 32539 32453 32548 32487
rect 32496 32444 32548 32453
rect 34336 32512 34388 32564
rect 34520 32444 34572 32496
rect 36360 32512 36412 32564
rect 36912 32555 36964 32564
rect 36912 32521 36921 32555
rect 36921 32521 36955 32555
rect 36955 32521 36964 32555
rect 36912 32512 36964 32521
rect 39580 32555 39632 32564
rect 39580 32521 39589 32555
rect 39589 32521 39623 32555
rect 39623 32521 39632 32555
rect 39580 32512 39632 32521
rect 33508 32419 33560 32428
rect 33508 32385 33517 32419
rect 33517 32385 33551 32419
rect 33551 32385 33560 32419
rect 33508 32376 33560 32385
rect 34428 32376 34480 32428
rect 34980 32419 35032 32428
rect 34980 32385 34989 32419
rect 34989 32385 35023 32419
rect 35023 32385 35032 32419
rect 34980 32376 35032 32385
rect 35256 32419 35308 32428
rect 35256 32385 35265 32419
rect 35265 32385 35299 32419
rect 35299 32385 35308 32419
rect 35256 32376 35308 32385
rect 35992 32376 36044 32428
rect 37924 32444 37976 32496
rect 38936 32444 38988 32496
rect 26792 32240 26844 32292
rect 23756 32172 23808 32224
rect 27712 32240 27764 32292
rect 31300 32240 31352 32292
rect 31852 32240 31904 32292
rect 36636 32308 36688 32360
rect 37740 32351 37792 32360
rect 37740 32317 37749 32351
rect 37749 32317 37783 32351
rect 37783 32317 37792 32351
rect 37740 32308 37792 32317
rect 37832 32308 37884 32360
rect 38844 32419 38896 32428
rect 38844 32385 38853 32419
rect 38853 32385 38887 32419
rect 38887 32385 38896 32419
rect 39948 32444 40000 32496
rect 38844 32376 38896 32385
rect 39488 32419 39540 32428
rect 39488 32385 39497 32419
rect 39497 32385 39531 32419
rect 39531 32385 39540 32419
rect 39488 32376 39540 32385
rect 42984 32419 43036 32428
rect 42984 32385 42993 32419
rect 42993 32385 43027 32419
rect 43027 32385 43036 32419
rect 42984 32376 43036 32385
rect 40960 32308 41012 32360
rect 42892 32308 42944 32360
rect 43260 32351 43312 32360
rect 43260 32317 43269 32351
rect 43269 32317 43303 32351
rect 43303 32317 43312 32351
rect 43260 32308 43312 32317
rect 28080 32172 28132 32224
rect 34612 32172 34664 32224
rect 34796 32172 34848 32224
rect 35716 32172 35768 32224
rect 37740 32172 37792 32224
rect 40408 32172 40460 32224
rect 42616 32215 42668 32224
rect 42616 32181 42625 32215
rect 42625 32181 42659 32215
rect 42659 32181 42668 32215
rect 42616 32172 42668 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4712 31968 4764 32020
rect 5264 31875 5316 31884
rect 5264 31841 5273 31875
rect 5273 31841 5307 31875
rect 5307 31841 5316 31875
rect 9680 31968 9732 32020
rect 10324 32011 10376 32020
rect 10324 31977 10333 32011
rect 10333 31977 10367 32011
rect 10367 31977 10376 32011
rect 10324 31968 10376 31977
rect 8024 31900 8076 31952
rect 5264 31832 5316 31841
rect 7380 31832 7432 31884
rect 7472 31832 7524 31884
rect 8208 31832 8260 31884
rect 11152 31968 11204 32020
rect 13084 31968 13136 32020
rect 10876 31900 10928 31952
rect 11244 31900 11296 31952
rect 13360 31943 13412 31952
rect 13360 31909 13369 31943
rect 13369 31909 13403 31943
rect 13403 31909 13412 31943
rect 13360 31900 13412 31909
rect 13912 31900 13964 31952
rect 16212 31968 16264 32020
rect 16304 31900 16356 31952
rect 22744 31968 22796 32020
rect 23388 31968 23440 32020
rect 27712 31968 27764 32020
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 7012 31764 7064 31816
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 8760 31764 8812 31816
rect 5356 31696 5408 31748
rect 6276 31696 6328 31748
rect 9864 31764 9916 31816
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 11980 31832 12032 31884
rect 14188 31832 14240 31884
rect 14280 31875 14332 31884
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14556 31807 14608 31816
rect 14556 31773 14590 31807
rect 14590 31773 14608 31807
rect 14556 31764 14608 31773
rect 18144 31764 18196 31816
rect 25136 31900 25188 31952
rect 26240 31900 26292 31952
rect 23388 31875 23440 31884
rect 23388 31841 23397 31875
rect 23397 31841 23431 31875
rect 23431 31841 23440 31875
rect 23388 31832 23440 31841
rect 27160 31832 27212 31884
rect 30840 31968 30892 32020
rect 31208 31968 31260 32020
rect 35256 31968 35308 32020
rect 35900 32011 35952 32020
rect 35900 31977 35909 32011
rect 35909 31977 35943 32011
rect 35943 31977 35952 32011
rect 35900 31968 35952 31977
rect 36084 31968 36136 32020
rect 36544 31968 36596 32020
rect 37464 32011 37516 32020
rect 37464 31977 37473 32011
rect 37473 31977 37507 32011
rect 37507 31977 37516 32011
rect 37464 31968 37516 31977
rect 40960 32011 41012 32020
rect 40960 31977 40969 32011
rect 40969 31977 41003 32011
rect 41003 31977 41012 32011
rect 40960 31968 41012 31977
rect 33140 31900 33192 31952
rect 20904 31764 20956 31816
rect 12440 31739 12492 31748
rect 12440 31705 12449 31739
rect 12449 31705 12483 31739
rect 12483 31705 12492 31739
rect 12440 31696 12492 31705
rect 13636 31696 13688 31748
rect 20996 31696 21048 31748
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22008 31807 22060 31816
rect 22008 31773 22017 31807
rect 22017 31773 22051 31807
rect 22051 31773 22060 31807
rect 22008 31764 22060 31773
rect 23112 31807 23164 31816
rect 23112 31773 23121 31807
rect 23121 31773 23155 31807
rect 23155 31773 23164 31807
rect 23112 31764 23164 31773
rect 23296 31807 23348 31816
rect 23296 31773 23305 31807
rect 23305 31773 23339 31807
rect 23339 31773 23348 31807
rect 23296 31764 23348 31773
rect 23480 31764 23532 31816
rect 24676 31764 24728 31816
rect 24860 31764 24912 31816
rect 25228 31764 25280 31816
rect 25872 31764 25924 31816
rect 26056 31764 26108 31816
rect 26240 31764 26292 31816
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 27896 31764 27948 31816
rect 25688 31696 25740 31748
rect 27068 31696 27120 31748
rect 28172 31764 28224 31816
rect 28448 31807 28500 31816
rect 28448 31773 28457 31807
rect 28457 31773 28491 31807
rect 28491 31773 28500 31807
rect 28448 31764 28500 31773
rect 28540 31807 28592 31816
rect 28540 31773 28549 31807
rect 28549 31773 28583 31807
rect 28583 31773 28592 31807
rect 28540 31764 28592 31773
rect 29736 31807 29788 31816
rect 29736 31773 29745 31807
rect 29745 31773 29779 31807
rect 29779 31773 29788 31807
rect 29736 31764 29788 31773
rect 29828 31764 29880 31816
rect 31024 31764 31076 31816
rect 32496 31832 32548 31884
rect 33508 31943 33560 31952
rect 33508 31909 33517 31943
rect 33517 31909 33551 31943
rect 33551 31909 33560 31943
rect 33508 31900 33560 31909
rect 34796 31900 34848 31952
rect 35440 31900 35492 31952
rect 35716 31900 35768 31952
rect 33232 31807 33284 31816
rect 33232 31773 33241 31807
rect 33241 31773 33275 31807
rect 33275 31773 33284 31807
rect 33232 31764 33284 31773
rect 33692 31764 33744 31816
rect 35164 31764 35216 31816
rect 36636 31900 36688 31952
rect 33324 31696 33376 31748
rect 8300 31628 8352 31680
rect 9220 31628 9272 31680
rect 10324 31628 10376 31680
rect 10692 31628 10744 31680
rect 11428 31628 11480 31680
rect 13820 31628 13872 31680
rect 22928 31671 22980 31680
rect 22928 31637 22937 31671
rect 22937 31637 22971 31671
rect 22971 31637 22980 31671
rect 22928 31628 22980 31637
rect 24952 31628 25004 31680
rect 25320 31628 25372 31680
rect 26240 31628 26292 31680
rect 29000 31671 29052 31680
rect 29000 31637 29009 31671
rect 29009 31637 29043 31671
rect 29043 31637 29052 31671
rect 29000 31628 29052 31637
rect 29092 31628 29144 31680
rect 36360 31832 36412 31884
rect 37096 31832 37148 31884
rect 38108 31832 38160 31884
rect 40040 31832 40092 31884
rect 41788 31968 41840 32020
rect 35992 31764 36044 31816
rect 36912 31807 36964 31816
rect 36912 31773 36922 31807
rect 36922 31773 36956 31807
rect 36956 31773 36964 31807
rect 36912 31764 36964 31773
rect 36636 31696 36688 31748
rect 37556 31764 37608 31816
rect 38476 31807 38528 31816
rect 38476 31773 38485 31807
rect 38485 31773 38519 31807
rect 38519 31773 38528 31807
rect 38476 31764 38528 31773
rect 38660 31764 38712 31816
rect 40408 31807 40460 31816
rect 40408 31773 40418 31807
rect 40418 31773 40452 31807
rect 40452 31773 40460 31807
rect 40408 31764 40460 31773
rect 37096 31739 37148 31748
rect 37096 31705 37105 31739
rect 37105 31705 37139 31739
rect 37139 31705 37148 31739
rect 37096 31696 37148 31705
rect 35900 31628 35952 31680
rect 35992 31628 36044 31680
rect 37464 31696 37516 31748
rect 38016 31696 38068 31748
rect 38568 31696 38620 31748
rect 38752 31696 38804 31748
rect 39580 31696 39632 31748
rect 40592 31739 40644 31748
rect 40592 31705 40601 31739
rect 40601 31705 40635 31739
rect 40635 31705 40644 31739
rect 40592 31696 40644 31705
rect 41052 31696 41104 31748
rect 42616 31764 42668 31816
rect 42984 31900 43036 31952
rect 39304 31628 39356 31680
rect 40776 31628 40828 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 7564 31424 7616 31476
rect 9312 31424 9364 31476
rect 9496 31467 9548 31476
rect 9496 31433 9505 31467
rect 9505 31433 9539 31467
rect 9539 31433 9548 31467
rect 9496 31424 9548 31433
rect 8024 31356 8076 31408
rect 9220 31356 9272 31408
rect 7288 31288 7340 31340
rect 7196 31220 7248 31272
rect 8300 31331 8352 31340
rect 8300 31297 8309 31331
rect 8309 31297 8343 31331
rect 8343 31297 8352 31331
rect 8300 31288 8352 31297
rect 9312 31331 9364 31340
rect 9312 31297 9321 31331
rect 9321 31297 9355 31331
rect 9355 31297 9364 31331
rect 10232 31424 10284 31476
rect 10600 31424 10652 31476
rect 9312 31288 9364 31297
rect 6184 31152 6236 31204
rect 7196 31084 7248 31136
rect 8116 31084 8168 31136
rect 8300 31152 8352 31204
rect 8668 31152 8720 31204
rect 9864 31152 9916 31204
rect 10416 31331 10468 31340
rect 10416 31297 10425 31331
rect 10425 31297 10459 31331
rect 10459 31297 10468 31331
rect 10416 31288 10468 31297
rect 10508 31331 10560 31340
rect 10508 31297 10517 31331
rect 10517 31297 10551 31331
rect 10551 31297 10560 31331
rect 10508 31288 10560 31297
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 13360 31424 13412 31476
rect 19984 31424 20036 31476
rect 32312 31424 32364 31476
rect 34152 31467 34204 31476
rect 34152 31433 34161 31467
rect 34161 31433 34195 31467
rect 34195 31433 34204 31467
rect 34152 31424 34204 31433
rect 34336 31424 34388 31476
rect 13912 31399 13964 31408
rect 13912 31365 13937 31399
rect 13937 31365 13964 31399
rect 13912 31356 13964 31365
rect 23112 31356 23164 31408
rect 11428 31220 11480 31272
rect 18236 31288 18288 31340
rect 22928 31288 22980 31340
rect 23848 31288 23900 31340
rect 24860 31220 24912 31272
rect 10692 31084 10744 31136
rect 12808 31084 12860 31136
rect 13820 31084 13872 31136
rect 15016 31084 15068 31136
rect 19340 31084 19392 31136
rect 24492 31152 24544 31204
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 26976 31288 27028 31340
rect 28080 31331 28132 31340
rect 28080 31297 28089 31331
rect 28089 31297 28123 31331
rect 28123 31297 28132 31331
rect 28080 31288 28132 31297
rect 28264 31288 28316 31340
rect 30012 31356 30064 31408
rect 30656 31356 30708 31408
rect 30104 31288 30156 31340
rect 30840 31331 30892 31340
rect 30840 31297 30849 31331
rect 30849 31297 30883 31331
rect 30883 31297 30892 31331
rect 30840 31288 30892 31297
rect 33416 31356 33468 31408
rect 34428 31356 34480 31408
rect 36084 31356 36136 31408
rect 32404 31331 32456 31340
rect 32404 31297 32413 31331
rect 32413 31297 32447 31331
rect 32447 31297 32456 31331
rect 32404 31288 32456 31297
rect 33324 31331 33376 31340
rect 33324 31297 33333 31331
rect 33333 31297 33367 31331
rect 33367 31297 33376 31331
rect 33324 31288 33376 31297
rect 34244 31331 34296 31340
rect 34244 31297 34253 31331
rect 34253 31297 34287 31331
rect 34287 31297 34296 31331
rect 34244 31288 34296 31297
rect 34704 31288 34756 31340
rect 26424 31263 26476 31272
rect 26424 31229 26433 31263
rect 26433 31229 26467 31263
rect 26467 31229 26476 31263
rect 26424 31220 26476 31229
rect 26516 31220 26568 31272
rect 32956 31220 33008 31272
rect 35440 31220 35492 31272
rect 35992 31288 36044 31340
rect 38016 31424 38068 31476
rect 38660 31424 38712 31476
rect 41052 31467 41104 31476
rect 41052 31433 41061 31467
rect 41061 31433 41095 31467
rect 41095 31433 41104 31467
rect 41052 31424 41104 31433
rect 36452 31331 36504 31340
rect 36452 31297 36461 31331
rect 36461 31297 36495 31331
rect 36495 31297 36504 31331
rect 36452 31288 36504 31297
rect 36544 31288 36596 31340
rect 29368 31152 29420 31204
rect 30012 31152 30064 31204
rect 23572 31084 23624 31136
rect 23664 31084 23716 31136
rect 24124 31084 24176 31136
rect 25228 31127 25280 31136
rect 25228 31093 25237 31127
rect 25237 31093 25271 31127
rect 25271 31093 25280 31127
rect 25228 31084 25280 31093
rect 26424 31084 26476 31136
rect 27068 31084 27120 31136
rect 31116 31127 31168 31136
rect 31116 31093 31125 31127
rect 31125 31093 31159 31127
rect 31159 31093 31168 31127
rect 31116 31084 31168 31093
rect 35348 31152 35400 31204
rect 35808 31152 35860 31204
rect 35900 31152 35952 31204
rect 36636 31152 36688 31204
rect 37280 31288 37332 31340
rect 37924 31331 37976 31340
rect 37924 31297 37933 31331
rect 37933 31297 37967 31331
rect 37967 31297 37976 31331
rect 37924 31288 37976 31297
rect 38016 31288 38068 31340
rect 38752 31356 38804 31408
rect 39120 31288 39172 31340
rect 39396 31288 39448 31340
rect 39488 31288 39540 31340
rect 43076 31288 43128 31340
rect 38844 31220 38896 31272
rect 39212 31220 39264 31272
rect 43168 31263 43220 31272
rect 43168 31229 43177 31263
rect 43177 31229 43211 31263
rect 43211 31229 43220 31263
rect 43168 31220 43220 31229
rect 34336 31084 34388 31136
rect 34520 31084 34572 31136
rect 36084 31084 36136 31136
rect 36912 31084 36964 31136
rect 38752 31084 38804 31136
rect 39212 31084 39264 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7012 30923 7064 30932
rect 7012 30889 7021 30923
rect 7021 30889 7055 30923
rect 7055 30889 7064 30923
rect 7012 30880 7064 30889
rect 7288 30880 7340 30932
rect 7472 30880 7524 30932
rect 20260 30880 20312 30932
rect 23572 30880 23624 30932
rect 24952 30880 25004 30932
rect 25136 30880 25188 30932
rect 25412 30880 25464 30932
rect 4620 30812 4672 30864
rect 6460 30744 6512 30796
rect 7380 30744 7432 30796
rect 8300 30744 8352 30796
rect 9496 30744 9548 30796
rect 6276 30676 6328 30728
rect 7104 30676 7156 30728
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8116 30676 8168 30685
rect 8208 30719 8260 30728
rect 8208 30685 8217 30719
rect 8217 30685 8251 30719
rect 8251 30685 8260 30719
rect 8208 30676 8260 30685
rect 8760 30676 8812 30728
rect 7564 30608 7616 30660
rect 9772 30787 9824 30796
rect 9772 30753 9781 30787
rect 9781 30753 9815 30787
rect 9815 30753 9824 30787
rect 9772 30744 9824 30753
rect 10416 30744 10468 30796
rect 10784 30744 10836 30796
rect 19984 30812 20036 30864
rect 9864 30719 9916 30728
rect 9864 30685 9873 30719
rect 9873 30685 9907 30719
rect 9907 30685 9916 30719
rect 9864 30676 9916 30685
rect 10508 30676 10560 30728
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11011 30719
rect 11011 30685 11020 30719
rect 10968 30676 11020 30685
rect 10692 30608 10744 30660
rect 11520 30676 11572 30728
rect 17592 30744 17644 30796
rect 18328 30744 18380 30796
rect 24124 30812 24176 30864
rect 25228 30812 25280 30864
rect 26700 30812 26752 30864
rect 12164 30676 12216 30728
rect 14280 30676 14332 30728
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 22376 30744 22428 30796
rect 23664 30787 23716 30796
rect 23664 30753 23673 30787
rect 23673 30753 23707 30787
rect 23707 30753 23716 30787
rect 23664 30744 23716 30753
rect 23848 30787 23900 30796
rect 23848 30753 23857 30787
rect 23857 30753 23891 30787
rect 23891 30753 23900 30787
rect 23848 30744 23900 30753
rect 25044 30744 25096 30796
rect 26424 30744 26476 30796
rect 27436 30744 27488 30796
rect 31576 30880 31628 30932
rect 32956 30812 33008 30864
rect 33508 30812 33560 30864
rect 33784 30812 33836 30864
rect 29276 30744 29328 30796
rect 20260 30676 20312 30728
rect 4804 30583 4856 30592
rect 4804 30549 4813 30583
rect 4813 30549 4847 30583
rect 4847 30549 4856 30583
rect 4804 30540 4856 30549
rect 5540 30540 5592 30592
rect 8576 30583 8628 30592
rect 8576 30549 8585 30583
rect 8585 30549 8619 30583
rect 8619 30549 8628 30583
rect 8576 30540 8628 30549
rect 9496 30583 9548 30592
rect 9496 30549 9505 30583
rect 9505 30549 9539 30583
rect 9539 30549 9548 30583
rect 9496 30540 9548 30549
rect 14648 30608 14700 30660
rect 18236 30651 18288 30660
rect 18236 30617 18245 30651
rect 18245 30617 18279 30651
rect 18279 30617 18288 30651
rect 18236 30608 18288 30617
rect 20168 30608 20220 30660
rect 20812 30651 20864 30660
rect 20812 30617 20821 30651
rect 20821 30617 20855 30651
rect 20855 30617 20864 30651
rect 20812 30608 20864 30617
rect 20996 30719 21048 30728
rect 20996 30685 21005 30719
rect 21005 30685 21039 30719
rect 21039 30685 21048 30719
rect 20996 30676 21048 30685
rect 25412 30676 25464 30728
rect 25872 30719 25924 30728
rect 25872 30685 25881 30719
rect 25881 30685 25915 30719
rect 25915 30685 25924 30719
rect 25872 30676 25924 30685
rect 26240 30676 26292 30728
rect 26976 30676 27028 30728
rect 29000 30676 29052 30728
rect 30656 30719 30708 30728
rect 30656 30685 30665 30719
rect 30665 30685 30699 30719
rect 30699 30685 30708 30719
rect 30656 30676 30708 30685
rect 30840 30676 30892 30728
rect 33140 30719 33192 30728
rect 33140 30685 33149 30719
rect 33149 30685 33183 30719
rect 33183 30685 33192 30719
rect 33140 30676 33192 30685
rect 33692 30676 33744 30728
rect 34244 30719 34296 30728
rect 34244 30685 34253 30719
rect 34253 30685 34287 30719
rect 34287 30685 34296 30719
rect 34244 30676 34296 30685
rect 36268 30880 36320 30932
rect 37004 30880 37056 30932
rect 37556 30880 37608 30932
rect 38936 30880 38988 30932
rect 39212 30880 39264 30932
rect 42984 30880 43036 30932
rect 36544 30812 36596 30864
rect 37464 30744 37516 30796
rect 34980 30719 35032 30728
rect 34980 30685 34989 30719
rect 34989 30685 35023 30719
rect 35023 30685 35032 30719
rect 34980 30676 35032 30685
rect 35164 30719 35216 30728
rect 35164 30685 35173 30719
rect 35173 30685 35207 30719
rect 35207 30685 35216 30719
rect 35164 30676 35216 30685
rect 36084 30719 36136 30728
rect 36084 30685 36093 30719
rect 36093 30685 36127 30719
rect 36127 30685 36136 30719
rect 36084 30676 36136 30685
rect 36176 30719 36228 30728
rect 36176 30685 36185 30719
rect 36185 30685 36219 30719
rect 36219 30685 36228 30719
rect 36176 30676 36228 30685
rect 36360 30719 36412 30728
rect 36360 30685 36369 30719
rect 36369 30685 36403 30719
rect 36403 30685 36412 30719
rect 36360 30676 36412 30685
rect 37556 30676 37608 30728
rect 38384 30676 38436 30728
rect 11704 30540 11756 30592
rect 14464 30540 14516 30592
rect 15936 30583 15988 30592
rect 15936 30549 15945 30583
rect 15945 30549 15979 30583
rect 15979 30549 15988 30583
rect 15936 30540 15988 30549
rect 17592 30540 17644 30592
rect 18880 30540 18932 30592
rect 20260 30583 20312 30592
rect 20260 30549 20269 30583
rect 20269 30549 20303 30583
rect 20303 30549 20312 30583
rect 20260 30540 20312 30549
rect 23204 30583 23256 30592
rect 23204 30549 23213 30583
rect 23213 30549 23247 30583
rect 23247 30549 23256 30583
rect 23204 30540 23256 30549
rect 23572 30583 23624 30592
rect 23572 30549 23581 30583
rect 23581 30549 23615 30583
rect 23615 30549 23624 30583
rect 23572 30540 23624 30549
rect 24860 30540 24912 30592
rect 27988 30583 28040 30592
rect 27988 30549 27997 30583
rect 27997 30549 28031 30583
rect 28031 30549 28040 30583
rect 27988 30540 28040 30549
rect 28448 30608 28500 30660
rect 29092 30608 29144 30660
rect 30932 30608 30984 30660
rect 32312 30608 32364 30660
rect 28632 30583 28684 30592
rect 28632 30549 28641 30583
rect 28641 30549 28675 30583
rect 28675 30549 28684 30583
rect 28632 30540 28684 30549
rect 31484 30583 31536 30592
rect 31484 30549 31493 30583
rect 31493 30549 31527 30583
rect 31527 30549 31536 30583
rect 31484 30540 31536 30549
rect 33416 30583 33468 30592
rect 33416 30549 33425 30583
rect 33425 30549 33459 30583
rect 33459 30549 33468 30583
rect 33416 30540 33468 30549
rect 33968 30651 34020 30660
rect 33968 30617 33977 30651
rect 33977 30617 34011 30651
rect 34011 30617 34020 30651
rect 33968 30608 34020 30617
rect 38108 30608 38160 30660
rect 38752 30719 38804 30728
rect 38752 30685 38761 30719
rect 38761 30685 38795 30719
rect 38795 30685 38804 30719
rect 38752 30676 38804 30685
rect 39580 30744 39632 30796
rect 40040 30787 40092 30796
rect 40040 30753 40049 30787
rect 40049 30753 40083 30787
rect 40083 30753 40092 30787
rect 40040 30744 40092 30753
rect 40408 30744 40460 30796
rect 41696 30744 41748 30796
rect 39120 30719 39172 30728
rect 39120 30685 39129 30719
rect 39129 30685 39163 30719
rect 39163 30685 39172 30719
rect 39120 30676 39172 30685
rect 40224 30676 40276 30728
rect 42616 30608 42668 30660
rect 37924 30540 37976 30592
rect 39212 30540 39264 30592
rect 43076 30540 43128 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5540 30379 5592 30388
rect 5540 30345 5549 30379
rect 5549 30345 5583 30379
rect 5583 30345 5592 30379
rect 5540 30336 5592 30345
rect 7472 30336 7524 30388
rect 14648 30336 14700 30388
rect 19432 30336 19484 30388
rect 20812 30336 20864 30388
rect 4620 30268 4672 30320
rect 9404 30268 9456 30320
rect 13820 30268 13872 30320
rect 14464 30268 14516 30320
rect 4804 30200 4856 30252
rect 9772 30200 9824 30252
rect 10692 30200 10744 30252
rect 11152 30243 11204 30252
rect 11152 30209 11161 30243
rect 11161 30209 11195 30243
rect 11195 30209 11204 30243
rect 11152 30200 11204 30209
rect 12348 30200 12400 30252
rect 13268 30243 13320 30252
rect 13268 30209 13277 30243
rect 13277 30209 13311 30243
rect 13311 30209 13320 30243
rect 13268 30200 13320 30209
rect 13912 30200 13964 30252
rect 11612 30132 11664 30184
rect 14372 30243 14424 30252
rect 14372 30209 14381 30243
rect 14381 30209 14415 30243
rect 14415 30209 14424 30243
rect 14372 30200 14424 30209
rect 17960 30243 18012 30252
rect 17960 30209 17969 30243
rect 17969 30209 18003 30243
rect 18003 30209 18012 30243
rect 17960 30200 18012 30209
rect 18880 30311 18932 30320
rect 18880 30277 18889 30311
rect 18889 30277 18923 30311
rect 18923 30277 18932 30311
rect 18880 30268 18932 30277
rect 19248 30268 19300 30320
rect 23572 30336 23624 30388
rect 25780 30336 25832 30388
rect 29276 30336 29328 30388
rect 29552 30336 29604 30388
rect 30288 30336 30340 30388
rect 31116 30336 31168 30388
rect 18972 30200 19024 30252
rect 15936 30132 15988 30184
rect 18420 30132 18472 30184
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 19800 30243 19852 30252
rect 19800 30209 19809 30243
rect 19809 30209 19843 30243
rect 19843 30209 19852 30243
rect 19800 30200 19852 30209
rect 20812 30200 20864 30252
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 21456 30243 21508 30252
rect 21456 30209 21465 30243
rect 21465 30209 21499 30243
rect 21499 30209 21508 30243
rect 21456 30200 21508 30209
rect 13176 30064 13228 30116
rect 10692 30039 10744 30048
rect 10692 30005 10701 30039
rect 10701 30005 10735 30039
rect 10735 30005 10744 30039
rect 10692 29996 10744 30005
rect 11612 29996 11664 30048
rect 18236 29996 18288 30048
rect 19248 30064 19300 30116
rect 24308 30243 24360 30252
rect 24308 30209 24317 30243
rect 24317 30209 24351 30243
rect 24351 30209 24360 30243
rect 24308 30200 24360 30209
rect 25044 30200 25096 30252
rect 23572 30132 23624 30184
rect 24492 30175 24544 30184
rect 24492 30141 24501 30175
rect 24501 30141 24535 30175
rect 24535 30141 24544 30175
rect 24492 30132 24544 30141
rect 19800 29996 19852 30048
rect 19892 29996 19944 30048
rect 20996 29996 21048 30048
rect 21456 29996 21508 30048
rect 24032 30064 24084 30116
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25596 30200 25648 30252
rect 25872 30268 25924 30320
rect 26332 30243 26384 30252
rect 26332 30209 26341 30243
rect 26341 30209 26375 30243
rect 26375 30209 26384 30243
rect 26332 30200 26384 30209
rect 28080 30243 28132 30252
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 28356 30243 28408 30252
rect 28356 30209 28365 30243
rect 28365 30209 28399 30243
rect 28399 30209 28408 30243
rect 28356 30200 28408 30209
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 29368 30200 29420 30252
rect 29552 30200 29604 30252
rect 24308 29996 24360 30048
rect 26056 30064 26108 30116
rect 28264 30064 28316 30116
rect 28724 30064 28776 30116
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 32404 30200 32456 30252
rect 31668 30132 31720 30184
rect 32312 30175 32364 30184
rect 32312 30141 32321 30175
rect 32321 30141 32355 30175
rect 32355 30141 32364 30175
rect 32312 30132 32364 30141
rect 30288 30064 30340 30116
rect 35164 30268 35216 30320
rect 34060 30200 34112 30252
rect 34520 30132 34572 30184
rect 34888 30200 34940 30252
rect 35440 30243 35492 30252
rect 35440 30209 35449 30243
rect 35449 30209 35483 30243
rect 35483 30209 35492 30243
rect 35440 30200 35492 30209
rect 35716 30336 35768 30388
rect 36176 30336 36228 30388
rect 37832 30336 37884 30388
rect 35716 30243 35768 30252
rect 35716 30209 35725 30243
rect 35725 30209 35759 30243
rect 35759 30209 35768 30243
rect 35716 30200 35768 30209
rect 35808 30243 35860 30252
rect 35808 30209 35817 30243
rect 35817 30209 35851 30243
rect 35851 30209 35860 30243
rect 35808 30200 35860 30209
rect 35900 30132 35952 30184
rect 30380 29996 30432 30048
rect 34796 30064 34848 30116
rect 34980 30064 35032 30116
rect 35532 30064 35584 30116
rect 36636 30200 36688 30252
rect 39212 30268 39264 30320
rect 42616 30379 42668 30388
rect 42616 30345 42625 30379
rect 42625 30345 42659 30379
rect 42659 30345 42668 30379
rect 42616 30336 42668 30345
rect 42984 30379 43036 30388
rect 42984 30345 42993 30379
rect 42993 30345 43027 30379
rect 43027 30345 43036 30379
rect 42984 30336 43036 30345
rect 43076 30379 43128 30388
rect 43076 30345 43085 30379
rect 43085 30345 43119 30379
rect 43119 30345 43128 30379
rect 43076 30336 43128 30345
rect 37280 30132 37332 30184
rect 37924 30175 37976 30184
rect 37924 30141 37933 30175
rect 37933 30141 37967 30175
rect 37967 30141 37976 30175
rect 37924 30132 37976 30141
rect 38108 30175 38160 30184
rect 38108 30141 38117 30175
rect 38117 30141 38151 30175
rect 38151 30141 38160 30175
rect 38108 30132 38160 30141
rect 38936 30132 38988 30184
rect 39304 30243 39356 30252
rect 39304 30209 39313 30243
rect 39313 30209 39347 30243
rect 39347 30209 39356 30243
rect 39304 30200 39356 30209
rect 40224 30268 40276 30320
rect 39948 30200 40000 30252
rect 40132 30175 40184 30184
rect 40132 30141 40141 30175
rect 40141 30141 40175 30175
rect 40175 30141 40184 30175
rect 40132 30132 40184 30141
rect 40316 30243 40368 30252
rect 40316 30209 40325 30243
rect 40325 30209 40359 30243
rect 40359 30209 40368 30243
rect 40316 30200 40368 30209
rect 43260 30064 43312 30116
rect 34336 29996 34388 30048
rect 36728 29996 36780 30048
rect 37096 29996 37148 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 37556 29996 37608 30048
rect 41052 29996 41104 30048
rect 41144 30039 41196 30048
rect 41144 30005 41153 30039
rect 41153 30005 41187 30039
rect 41187 30005 41196 30039
rect 41144 29996 41196 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 9220 29792 9272 29844
rect 11520 29792 11572 29844
rect 11612 29835 11664 29844
rect 11612 29801 11621 29835
rect 11621 29801 11655 29835
rect 11655 29801 11664 29835
rect 11612 29792 11664 29801
rect 17224 29792 17276 29844
rect 8116 29724 8168 29776
rect 18788 29835 18840 29844
rect 18788 29801 18797 29835
rect 18797 29801 18831 29835
rect 18831 29801 18840 29835
rect 18788 29792 18840 29801
rect 19248 29792 19300 29844
rect 22836 29792 22888 29844
rect 23572 29835 23624 29844
rect 23572 29801 23581 29835
rect 23581 29801 23615 29835
rect 23615 29801 23624 29835
rect 23572 29792 23624 29801
rect 24308 29792 24360 29844
rect 32128 29792 32180 29844
rect 33232 29792 33284 29844
rect 33324 29792 33376 29844
rect 33968 29792 34020 29844
rect 34520 29792 34572 29844
rect 35532 29792 35584 29844
rect 36176 29792 36228 29844
rect 36636 29792 36688 29844
rect 7104 29656 7156 29708
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 18052 29656 18104 29708
rect 18236 29656 18288 29708
rect 6644 29495 6696 29504
rect 6644 29461 6653 29495
rect 6653 29461 6687 29495
rect 6687 29461 6696 29495
rect 6644 29452 6696 29461
rect 7104 29520 7156 29572
rect 7380 29520 7432 29572
rect 7840 29520 7892 29572
rect 9312 29588 9364 29640
rect 11704 29588 11756 29640
rect 12348 29588 12400 29640
rect 12808 29631 12860 29640
rect 12808 29597 12817 29631
rect 12817 29597 12851 29631
rect 12851 29597 12860 29631
rect 12808 29588 12860 29597
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 17776 29588 17828 29640
rect 18972 29656 19024 29708
rect 20260 29656 20312 29708
rect 10692 29520 10744 29572
rect 8392 29452 8444 29504
rect 13360 29452 13412 29504
rect 16212 29495 16264 29504
rect 16212 29461 16221 29495
rect 16221 29461 16255 29495
rect 16255 29461 16264 29495
rect 16212 29452 16264 29461
rect 16580 29495 16632 29504
rect 16580 29461 16589 29495
rect 16589 29461 16623 29495
rect 16623 29461 16632 29495
rect 16580 29452 16632 29461
rect 16856 29452 16908 29504
rect 18236 29452 18288 29504
rect 19800 29631 19852 29640
rect 19800 29597 19809 29631
rect 19809 29597 19843 29631
rect 19843 29597 19852 29631
rect 19800 29588 19852 29597
rect 19892 29631 19944 29640
rect 19892 29597 19901 29631
rect 19901 29597 19935 29631
rect 19935 29597 19944 29631
rect 19892 29588 19944 29597
rect 20812 29588 20864 29640
rect 25688 29724 25740 29776
rect 22928 29699 22980 29708
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 23204 29656 23256 29708
rect 30012 29724 30064 29776
rect 27252 29656 27304 29708
rect 30104 29699 30156 29708
rect 30104 29665 30113 29699
rect 30113 29665 30147 29699
rect 30147 29665 30156 29699
rect 30104 29656 30156 29665
rect 30380 29699 30432 29708
rect 30380 29665 30389 29699
rect 30389 29665 30423 29699
rect 30423 29665 30432 29699
rect 30380 29656 30432 29665
rect 31300 29656 31352 29708
rect 31576 29656 31628 29708
rect 25320 29588 25372 29640
rect 26976 29631 27028 29640
rect 26976 29597 26985 29631
rect 26985 29597 27019 29631
rect 27019 29597 27028 29631
rect 26976 29588 27028 29597
rect 27988 29631 28040 29640
rect 27988 29597 27997 29631
rect 27997 29597 28031 29631
rect 28031 29597 28040 29631
rect 27988 29588 28040 29597
rect 28080 29588 28132 29640
rect 31392 29588 31444 29640
rect 19340 29520 19392 29572
rect 22376 29520 22428 29572
rect 26516 29520 26568 29572
rect 27528 29520 27580 29572
rect 19432 29452 19484 29504
rect 23204 29495 23256 29504
rect 23204 29461 23213 29495
rect 23213 29461 23247 29495
rect 23247 29461 23256 29495
rect 31116 29520 31168 29572
rect 31208 29520 31260 29572
rect 31852 29631 31904 29640
rect 31852 29597 31861 29631
rect 31861 29597 31895 29631
rect 31895 29597 31904 29631
rect 31852 29588 31904 29597
rect 32128 29588 32180 29640
rect 32956 29631 33008 29640
rect 32956 29597 32965 29631
rect 32965 29597 32999 29631
rect 32999 29597 33008 29631
rect 32956 29588 33008 29597
rect 33140 29631 33192 29640
rect 33140 29597 33147 29631
rect 33147 29597 33192 29631
rect 33140 29588 33192 29597
rect 33416 29631 33468 29640
rect 33416 29597 33449 29631
rect 33449 29597 33468 29631
rect 33416 29588 33468 29597
rect 31760 29520 31812 29572
rect 34520 29588 34572 29640
rect 35808 29656 35860 29708
rect 34980 29631 35032 29640
rect 34980 29597 34989 29631
rect 34989 29597 35023 29631
rect 35023 29597 35032 29631
rect 34980 29588 35032 29597
rect 34152 29520 34204 29572
rect 35992 29588 36044 29640
rect 36728 29520 36780 29572
rect 23204 29452 23256 29461
rect 28724 29495 28776 29504
rect 28724 29461 28733 29495
rect 28733 29461 28767 29495
rect 28767 29461 28776 29495
rect 28724 29452 28776 29461
rect 30472 29452 30524 29504
rect 37096 29588 37148 29640
rect 41696 29792 41748 29844
rect 41144 29588 41196 29640
rect 37464 29520 37516 29572
rect 37924 29520 37976 29572
rect 43168 29563 43220 29572
rect 43168 29529 43177 29563
rect 43177 29529 43211 29563
rect 43211 29529 43220 29563
rect 43168 29520 43220 29529
rect 39396 29452 39448 29504
rect 40040 29452 40092 29504
rect 41052 29452 41104 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 8300 29248 8352 29300
rect 9220 29248 9272 29300
rect 16856 29291 16908 29300
rect 16856 29257 16865 29291
rect 16865 29257 16899 29291
rect 16899 29257 16908 29291
rect 16856 29248 16908 29257
rect 18052 29291 18104 29300
rect 18052 29257 18061 29291
rect 18061 29257 18095 29291
rect 18095 29257 18104 29291
rect 18052 29248 18104 29257
rect 6920 29112 6972 29164
rect 9128 29180 9180 29232
rect 17224 29223 17276 29232
rect 17224 29189 17233 29223
rect 17233 29189 17267 29223
rect 17267 29189 17276 29223
rect 17224 29180 17276 29189
rect 19340 29248 19392 29300
rect 26148 29248 26200 29300
rect 28080 29248 28132 29300
rect 28632 29248 28684 29300
rect 7932 29155 7984 29164
rect 7932 29121 7966 29155
rect 7966 29121 7984 29155
rect 7932 29112 7984 29121
rect 8208 29112 8260 29164
rect 11704 29112 11756 29164
rect 13636 29155 13688 29164
rect 13636 29121 13670 29155
rect 13670 29121 13688 29155
rect 13636 29112 13688 29121
rect 15936 29112 15988 29164
rect 17868 29112 17920 29164
rect 18420 29112 18472 29164
rect 18512 29155 18564 29164
rect 18512 29121 18521 29155
rect 18521 29121 18555 29155
rect 18555 29121 18564 29155
rect 18512 29112 18564 29121
rect 13176 29044 13228 29096
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 17592 29044 17644 29096
rect 14464 28976 14516 29028
rect 17868 28976 17920 29028
rect 22928 29180 22980 29232
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 19984 29112 20036 29164
rect 26424 29112 26476 29164
rect 27896 29180 27948 29232
rect 28356 29223 28408 29232
rect 28356 29189 28365 29223
rect 28365 29189 28399 29223
rect 28399 29189 28408 29223
rect 28356 29180 28408 29189
rect 28724 29180 28776 29232
rect 19156 29044 19208 29096
rect 25412 29087 25464 29096
rect 19064 28976 19116 29028
rect 25412 29053 25421 29087
rect 25421 29053 25455 29087
rect 25455 29053 25464 29087
rect 25412 29044 25464 29053
rect 26700 29044 26752 29096
rect 28540 29112 28592 29164
rect 29828 29112 29880 29164
rect 28448 29044 28500 29096
rect 31116 29248 31168 29300
rect 32312 29248 32364 29300
rect 34520 29248 34572 29300
rect 32404 29180 32456 29232
rect 30748 29112 30800 29164
rect 31116 29112 31168 29164
rect 31484 29112 31536 29164
rect 33232 29180 33284 29232
rect 36728 29248 36780 29300
rect 37372 29248 37424 29300
rect 38476 29248 38528 29300
rect 39212 29248 39264 29300
rect 35624 29223 35676 29232
rect 35624 29189 35633 29223
rect 35633 29189 35667 29223
rect 35667 29189 35676 29223
rect 35624 29180 35676 29189
rect 33140 29155 33192 29164
rect 33140 29121 33149 29155
rect 33149 29121 33183 29155
rect 33183 29121 33192 29155
rect 33140 29112 33192 29121
rect 34428 29155 34480 29164
rect 34428 29121 34437 29155
rect 34437 29121 34471 29155
rect 34471 29121 34480 29155
rect 34428 29112 34480 29121
rect 31300 29044 31352 29096
rect 33968 29044 34020 29096
rect 34796 29155 34848 29164
rect 34796 29121 34805 29155
rect 34805 29121 34839 29155
rect 34839 29121 34848 29155
rect 34796 29112 34848 29121
rect 35992 29112 36044 29164
rect 37280 29112 37332 29164
rect 37556 29112 37608 29164
rect 37648 29112 37700 29164
rect 38292 29112 38344 29164
rect 38660 29112 38712 29164
rect 39120 29155 39172 29164
rect 39120 29121 39127 29155
rect 39127 29121 39172 29155
rect 39120 29112 39172 29121
rect 39212 29155 39264 29164
rect 39212 29121 39221 29155
rect 39221 29121 39255 29155
rect 39255 29121 39264 29155
rect 39212 29112 39264 29121
rect 14004 28908 14056 28960
rect 14648 28908 14700 28960
rect 26056 28976 26108 29028
rect 22560 28908 22612 28960
rect 27436 28976 27488 29028
rect 34796 28976 34848 29028
rect 38108 29044 38160 29096
rect 38200 29044 38252 29096
rect 38752 29044 38804 29096
rect 39396 29155 39448 29164
rect 39396 29121 39410 29155
rect 39410 29121 39444 29155
rect 39444 29121 39448 29155
rect 39396 29112 39448 29121
rect 39948 29180 40000 29232
rect 41052 29291 41104 29300
rect 41052 29257 41061 29291
rect 41061 29257 41095 29291
rect 41095 29257 41104 29291
rect 41052 29248 41104 29257
rect 40132 29155 40184 29164
rect 40132 29121 40141 29155
rect 40141 29121 40175 29155
rect 40175 29121 40184 29155
rect 40132 29112 40184 29121
rect 40316 29155 40368 29164
rect 40316 29121 40325 29155
rect 40325 29121 40359 29155
rect 40359 29121 40368 29155
rect 40316 29112 40368 29121
rect 41144 29155 41196 29164
rect 41144 29121 41153 29155
rect 41153 29121 41187 29155
rect 41187 29121 41196 29155
rect 41144 29112 41196 29121
rect 40224 29044 40276 29096
rect 40040 28976 40092 29028
rect 32036 28908 32088 28960
rect 36912 28908 36964 28960
rect 37372 28908 37424 28960
rect 39304 28908 39356 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 7932 28704 7984 28756
rect 8116 28704 8168 28756
rect 11152 28704 11204 28756
rect 12348 28704 12400 28756
rect 13636 28704 13688 28756
rect 7104 28636 7156 28688
rect 8208 28636 8260 28688
rect 5632 28500 5684 28552
rect 6828 28500 6880 28552
rect 8116 28500 8168 28552
rect 8300 28543 8352 28552
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 8576 28543 8628 28552
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 9404 28543 9456 28552
rect 9404 28509 9438 28543
rect 9438 28509 9456 28543
rect 9404 28500 9456 28509
rect 12716 28500 12768 28552
rect 14464 28568 14516 28620
rect 14004 28500 14056 28552
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 18512 28704 18564 28756
rect 20904 28747 20956 28756
rect 20904 28713 20913 28747
rect 20913 28713 20947 28747
rect 20947 28713 20956 28747
rect 20904 28704 20956 28713
rect 22836 28747 22888 28756
rect 22836 28713 22845 28747
rect 22845 28713 22879 28747
rect 22879 28713 22888 28747
rect 22836 28704 22888 28713
rect 27160 28704 27212 28756
rect 32496 28704 32548 28756
rect 32956 28704 33008 28756
rect 36912 28704 36964 28756
rect 38108 28704 38160 28756
rect 39120 28704 39172 28756
rect 16580 28636 16632 28688
rect 19524 28636 19576 28688
rect 27620 28636 27672 28688
rect 28264 28636 28316 28688
rect 18420 28611 18472 28620
rect 18420 28577 18429 28611
rect 18429 28577 18463 28611
rect 18463 28577 18472 28611
rect 18420 28568 18472 28577
rect 6644 28432 6696 28484
rect 8392 28475 8444 28484
rect 8392 28441 8401 28475
rect 8401 28441 8435 28475
rect 8435 28441 8444 28475
rect 8392 28432 8444 28441
rect 12440 28432 12492 28484
rect 13360 28475 13412 28484
rect 13360 28441 13369 28475
rect 13369 28441 13403 28475
rect 13403 28441 13412 28475
rect 13360 28432 13412 28441
rect 13820 28432 13872 28484
rect 14740 28500 14792 28552
rect 15200 28500 15252 28552
rect 18144 28500 18196 28552
rect 14464 28475 14516 28484
rect 14464 28441 14473 28475
rect 14473 28441 14507 28475
rect 14507 28441 14516 28475
rect 14464 28432 14516 28441
rect 14832 28407 14884 28416
rect 14832 28373 14841 28407
rect 14841 28373 14875 28407
rect 14875 28373 14884 28407
rect 14832 28364 14884 28373
rect 16212 28432 16264 28484
rect 21548 28500 21600 28552
rect 24584 28568 24636 28620
rect 20076 28432 20128 28484
rect 20444 28432 20496 28484
rect 17684 28364 17736 28416
rect 17960 28364 18012 28416
rect 18512 28364 18564 28416
rect 19524 28364 19576 28416
rect 20812 28432 20864 28484
rect 20904 28432 20956 28484
rect 23020 28500 23072 28552
rect 23204 28500 23256 28552
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 23112 28475 23164 28484
rect 23112 28441 23121 28475
rect 23121 28441 23155 28475
rect 23155 28441 23164 28475
rect 23112 28432 23164 28441
rect 24124 28432 24176 28484
rect 27160 28475 27212 28484
rect 27160 28441 27169 28475
rect 27169 28441 27203 28475
rect 27203 28441 27212 28475
rect 27160 28432 27212 28441
rect 21088 28364 21140 28416
rect 23020 28364 23072 28416
rect 26424 28364 26476 28416
rect 27988 28543 28040 28552
rect 27988 28509 27997 28543
rect 27997 28509 28031 28543
rect 28031 28509 28040 28543
rect 27988 28500 28040 28509
rect 30380 28636 30432 28688
rect 28908 28568 28960 28620
rect 39028 28636 39080 28688
rect 32496 28568 32548 28620
rect 34152 28568 34204 28620
rect 29460 28500 29512 28552
rect 29828 28500 29880 28552
rect 30288 28500 30340 28552
rect 30472 28543 30524 28552
rect 30472 28509 30481 28543
rect 30481 28509 30515 28543
rect 30515 28509 30524 28543
rect 30472 28500 30524 28509
rect 30840 28500 30892 28552
rect 31208 28500 31260 28552
rect 31576 28500 31628 28552
rect 32036 28500 32088 28552
rect 32220 28500 32272 28552
rect 32588 28500 32640 28552
rect 33232 28543 33284 28552
rect 33232 28509 33241 28543
rect 33241 28509 33275 28543
rect 33275 28509 33284 28543
rect 33232 28500 33284 28509
rect 34336 28500 34388 28552
rect 35072 28500 35124 28552
rect 29552 28364 29604 28416
rect 31208 28364 31260 28416
rect 31852 28432 31904 28484
rect 32864 28432 32916 28484
rect 33140 28432 33192 28484
rect 34244 28432 34296 28484
rect 34428 28432 34480 28484
rect 35440 28500 35492 28552
rect 36912 28543 36964 28552
rect 36912 28509 36921 28543
rect 36921 28509 36955 28543
rect 36955 28509 36964 28543
rect 36912 28500 36964 28509
rect 37648 28568 37700 28620
rect 37372 28543 37424 28552
rect 37372 28509 37381 28543
rect 37381 28509 37415 28543
rect 37415 28509 37424 28543
rect 37372 28500 37424 28509
rect 37556 28543 37608 28552
rect 37556 28509 37565 28543
rect 37565 28509 37599 28543
rect 37599 28509 37608 28543
rect 37556 28500 37608 28509
rect 38844 28543 38896 28552
rect 38844 28509 38853 28543
rect 38853 28509 38887 28543
rect 38887 28509 38896 28543
rect 38844 28500 38896 28509
rect 35256 28432 35308 28484
rect 42984 28704 43036 28756
rect 40224 28568 40276 28620
rect 39304 28543 39356 28552
rect 39304 28509 39318 28543
rect 39318 28509 39352 28543
rect 39352 28509 39356 28543
rect 39304 28500 39356 28509
rect 40040 28543 40092 28552
rect 40040 28509 40049 28543
rect 40049 28509 40083 28543
rect 40083 28509 40092 28543
rect 40040 28500 40092 28509
rect 40316 28543 40368 28552
rect 40316 28509 40325 28543
rect 40325 28509 40359 28543
rect 40359 28509 40368 28543
rect 40316 28500 40368 28509
rect 41880 28543 41932 28552
rect 41880 28509 41889 28543
rect 41889 28509 41923 28543
rect 41923 28509 41932 28543
rect 41880 28500 41932 28509
rect 39028 28432 39080 28484
rect 42616 28432 42668 28484
rect 34612 28364 34664 28416
rect 36912 28364 36964 28416
rect 37372 28364 37424 28416
rect 39488 28364 39540 28416
rect 43076 28364 43128 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 7012 28203 7064 28212
rect 7012 28169 7021 28203
rect 7021 28169 7055 28203
rect 7055 28169 7064 28203
rect 7012 28160 7064 28169
rect 12072 28160 12124 28212
rect 14280 28160 14332 28212
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 17684 28203 17736 28212
rect 17684 28169 17693 28203
rect 17693 28169 17727 28203
rect 17727 28169 17736 28203
rect 17684 28160 17736 28169
rect 18420 28160 18472 28212
rect 20904 28160 20956 28212
rect 24124 28160 24176 28212
rect 27988 28160 28040 28212
rect 6920 28067 6972 28076
rect 6920 28033 6929 28067
rect 6929 28033 6963 28067
rect 6963 28033 6972 28067
rect 6920 28024 6972 28033
rect 7840 28024 7892 28076
rect 8944 28024 8996 28076
rect 13452 28092 13504 28144
rect 14832 28092 14884 28144
rect 22928 28092 22980 28144
rect 12348 28067 12400 28076
rect 12348 28033 12357 28067
rect 12357 28033 12391 28067
rect 12391 28033 12400 28067
rect 12348 28024 12400 28033
rect 13360 28024 13412 28076
rect 14464 28024 14516 28076
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 12440 27956 12492 28008
rect 16672 27956 16724 28008
rect 19064 28024 19116 28076
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 18236 27956 18288 28008
rect 21364 27999 21416 28008
rect 21364 27965 21373 27999
rect 21373 27965 21407 27999
rect 21407 27965 21416 27999
rect 21364 27956 21416 27965
rect 23296 27999 23348 28008
rect 23296 27965 23305 27999
rect 23305 27965 23339 27999
rect 23339 27965 23348 27999
rect 23296 27956 23348 27965
rect 23572 28024 23624 28076
rect 24032 27999 24084 28008
rect 24032 27965 24041 27999
rect 24041 27965 24075 27999
rect 24075 27965 24084 27999
rect 24032 27956 24084 27965
rect 24676 28092 24728 28144
rect 26884 28092 26936 28144
rect 27712 28092 27764 28144
rect 28632 28092 28684 28144
rect 29644 28092 29696 28144
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 24952 28024 25004 28076
rect 25412 28024 25464 28076
rect 25044 27956 25096 28008
rect 27160 28024 27212 28076
rect 29368 28024 29420 28076
rect 29736 28024 29788 28076
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 35256 28160 35308 28212
rect 40316 28160 40368 28212
rect 42616 28203 42668 28212
rect 42616 28169 42625 28203
rect 42625 28169 42659 28203
rect 42659 28169 42668 28203
rect 42616 28160 42668 28169
rect 42984 28203 43036 28212
rect 42984 28169 42993 28203
rect 42993 28169 43027 28203
rect 43027 28169 43036 28203
rect 42984 28160 43036 28169
rect 43076 28203 43128 28212
rect 43076 28169 43085 28203
rect 43085 28169 43119 28203
rect 43119 28169 43128 28203
rect 43076 28160 43128 28169
rect 31760 28092 31812 28144
rect 33508 28135 33560 28144
rect 33508 28101 33517 28135
rect 33517 28101 33551 28135
rect 33551 28101 33560 28135
rect 33508 28092 33560 28101
rect 31668 28024 31720 28076
rect 28356 27999 28408 28008
rect 28356 27965 28365 27999
rect 28365 27965 28399 27999
rect 28399 27965 28408 27999
rect 28356 27956 28408 27965
rect 28448 27999 28500 28008
rect 28448 27965 28457 27999
rect 28457 27965 28491 27999
rect 28491 27965 28500 27999
rect 28448 27956 28500 27965
rect 28540 27999 28592 28008
rect 28540 27965 28549 27999
rect 28549 27965 28583 27999
rect 28583 27965 28592 27999
rect 28540 27956 28592 27965
rect 28632 27999 28684 28008
rect 28632 27965 28641 27999
rect 28641 27965 28675 27999
rect 28675 27965 28684 27999
rect 28632 27956 28684 27965
rect 32588 28067 32640 28076
rect 32588 28033 32597 28067
rect 32597 28033 32631 28067
rect 32631 28033 32640 28067
rect 32588 28024 32640 28033
rect 32772 28024 32824 28076
rect 32036 27956 32088 28008
rect 32956 27956 33008 28008
rect 33232 27956 33284 28008
rect 13820 27931 13872 27940
rect 13820 27897 13829 27931
rect 13829 27897 13863 27931
rect 13863 27897 13872 27931
rect 13820 27888 13872 27897
rect 20812 27888 20864 27940
rect 36084 28092 36136 28144
rect 37096 28092 37148 28144
rect 37648 28092 37700 28144
rect 38844 28092 38896 28144
rect 34336 28024 34388 28076
rect 35072 28024 35124 28076
rect 35624 28024 35676 28076
rect 35992 28067 36044 28076
rect 35992 28033 36001 28067
rect 36001 28033 36035 28067
rect 36035 28033 36044 28067
rect 35992 28024 36044 28033
rect 37832 28067 37884 28076
rect 34428 27956 34480 28008
rect 37832 28033 37841 28067
rect 37841 28033 37875 28067
rect 37875 28033 37884 28067
rect 37832 28024 37884 28033
rect 39488 28067 39540 28076
rect 39488 28033 39497 28067
rect 39497 28033 39531 28067
rect 39531 28033 39540 28067
rect 39488 28024 39540 28033
rect 36912 27888 36964 27940
rect 37924 27999 37976 28008
rect 37924 27965 37933 27999
rect 37933 27965 37967 27999
rect 37967 27965 37976 27999
rect 37924 27956 37976 27965
rect 43260 27999 43312 28008
rect 43260 27965 43269 27999
rect 43269 27965 43303 27999
rect 43303 27965 43312 27999
rect 43260 27956 43312 27965
rect 38752 27888 38804 27940
rect 5540 27820 5592 27872
rect 8208 27863 8260 27872
rect 8208 27829 8217 27863
rect 8217 27829 8251 27863
rect 8251 27829 8260 27863
rect 8208 27820 8260 27829
rect 12532 27863 12584 27872
rect 12532 27829 12541 27863
rect 12541 27829 12575 27863
rect 12575 27829 12584 27863
rect 12532 27820 12584 27829
rect 20720 27863 20772 27872
rect 20720 27829 20729 27863
rect 20729 27829 20763 27863
rect 20763 27829 20772 27863
rect 20720 27820 20772 27829
rect 24124 27820 24176 27872
rect 27712 27820 27764 27872
rect 27804 27820 27856 27872
rect 30840 27820 30892 27872
rect 32312 27863 32364 27872
rect 32312 27829 32321 27863
rect 32321 27829 32355 27863
rect 32355 27829 32364 27863
rect 32312 27820 32364 27829
rect 32404 27820 32456 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 17960 27548 18012 27600
rect 8208 27480 8260 27532
rect 11704 27523 11756 27532
rect 11704 27489 11713 27523
rect 11713 27489 11747 27523
rect 11747 27489 11756 27523
rect 11704 27480 11756 27489
rect 22560 27616 22612 27668
rect 23204 27616 23256 27668
rect 25780 27616 25832 27668
rect 23572 27548 23624 27600
rect 24676 27548 24728 27600
rect 25964 27659 26016 27668
rect 25964 27625 25973 27659
rect 25973 27625 26007 27659
rect 26007 27625 26016 27659
rect 25964 27616 26016 27625
rect 21640 27480 21692 27532
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 8116 27412 8168 27464
rect 9128 27412 9180 27464
rect 10968 27412 11020 27464
rect 5540 27387 5592 27396
rect 5540 27353 5574 27387
rect 5574 27353 5592 27387
rect 5540 27344 5592 27353
rect 5632 27344 5684 27396
rect 6920 27344 6972 27396
rect 7748 27319 7800 27328
rect 7748 27285 7757 27319
rect 7757 27285 7791 27319
rect 7791 27285 7800 27319
rect 7748 27276 7800 27285
rect 8392 27387 8444 27396
rect 8392 27353 8401 27387
rect 8401 27353 8435 27387
rect 8435 27353 8444 27387
rect 8392 27344 8444 27353
rect 10324 27344 10376 27396
rect 16488 27412 16540 27464
rect 16580 27455 16632 27464
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 18788 27412 18840 27464
rect 20352 27412 20404 27464
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 20720 27412 20772 27464
rect 23020 27412 23072 27464
rect 12164 27344 12216 27396
rect 10692 27276 10744 27328
rect 21180 27344 21232 27396
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 24860 27480 24912 27532
rect 26608 27548 26660 27600
rect 32772 27616 32824 27668
rect 34520 27616 34572 27668
rect 35992 27616 36044 27668
rect 37096 27616 37148 27668
rect 29552 27548 29604 27600
rect 30564 27548 30616 27600
rect 31024 27548 31076 27600
rect 31576 27548 31628 27600
rect 32956 27548 33008 27600
rect 33968 27548 34020 27600
rect 26976 27480 27028 27532
rect 25044 27455 25096 27464
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 17132 27276 17184 27328
rect 18696 27276 18748 27328
rect 20812 27276 20864 27328
rect 21088 27276 21140 27328
rect 22744 27276 22796 27328
rect 23020 27319 23072 27328
rect 23020 27285 23029 27319
rect 23029 27285 23063 27319
rect 23063 27285 23072 27319
rect 23020 27276 23072 27285
rect 23204 27276 23256 27328
rect 25044 27421 25053 27455
rect 25053 27421 25087 27455
rect 25087 27421 25096 27455
rect 25044 27412 25096 27421
rect 25688 27387 25740 27396
rect 25688 27353 25697 27387
rect 25697 27353 25731 27387
rect 25731 27353 25740 27387
rect 25688 27344 25740 27353
rect 26516 27412 26568 27464
rect 27068 27412 27120 27464
rect 27436 27455 27488 27464
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 27528 27455 27580 27464
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 29736 27412 29788 27464
rect 30012 27455 30064 27464
rect 30012 27421 30021 27455
rect 30021 27421 30055 27455
rect 30055 27421 30064 27455
rect 30012 27412 30064 27421
rect 31944 27480 31996 27532
rect 32036 27480 32088 27532
rect 30932 27455 30984 27464
rect 30932 27421 30941 27455
rect 30941 27421 30975 27455
rect 30975 27421 30984 27455
rect 30932 27412 30984 27421
rect 31668 27412 31720 27464
rect 32588 27480 32640 27532
rect 33876 27480 33928 27532
rect 34796 27480 34848 27532
rect 33140 27412 33192 27464
rect 34980 27455 35032 27464
rect 34980 27421 34989 27455
rect 34989 27421 35023 27455
rect 35023 27421 35032 27455
rect 34980 27412 35032 27421
rect 35624 27548 35676 27600
rect 29276 27344 29328 27396
rect 25228 27319 25280 27328
rect 25228 27285 25237 27319
rect 25237 27285 25271 27319
rect 25271 27285 25280 27319
rect 25228 27276 25280 27285
rect 26516 27276 26568 27328
rect 27344 27276 27396 27328
rect 31760 27344 31812 27396
rect 32956 27344 33008 27396
rect 36084 27455 36136 27464
rect 36084 27421 36093 27455
rect 36093 27421 36127 27455
rect 36127 27421 36136 27455
rect 36084 27412 36136 27421
rect 36360 27455 36412 27464
rect 36360 27421 36369 27455
rect 36369 27421 36403 27455
rect 36403 27421 36412 27455
rect 36360 27412 36412 27421
rect 37096 27455 37148 27464
rect 37096 27421 37105 27455
rect 37105 27421 37139 27455
rect 37139 27421 37148 27455
rect 37096 27412 37148 27421
rect 38384 27548 38436 27600
rect 39028 27548 39080 27600
rect 40132 27548 40184 27600
rect 35440 27344 35492 27396
rect 36728 27344 36780 27396
rect 39028 27455 39080 27464
rect 39028 27421 39037 27455
rect 39037 27421 39071 27455
rect 39071 27421 39080 27455
rect 39028 27412 39080 27421
rect 40684 27412 40736 27464
rect 43996 27480 44048 27532
rect 41880 27412 41932 27464
rect 43076 27412 43128 27464
rect 29736 27319 29788 27328
rect 29736 27285 29745 27319
rect 29745 27285 29779 27319
rect 29779 27285 29788 27319
rect 29736 27276 29788 27285
rect 30932 27276 30984 27328
rect 32772 27276 32824 27328
rect 34704 27276 34756 27328
rect 36084 27276 36136 27328
rect 38476 27319 38528 27328
rect 38476 27285 38485 27319
rect 38485 27285 38519 27319
rect 38519 27285 38528 27319
rect 38476 27276 38528 27285
rect 40316 27344 40368 27396
rect 40776 27276 40828 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8116 27072 8168 27124
rect 9128 27004 9180 27056
rect 7748 26936 7800 26988
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 10324 27115 10376 27124
rect 10324 27081 10333 27115
rect 10333 27081 10367 27115
rect 10367 27081 10376 27115
rect 10324 27072 10376 27081
rect 10692 27115 10744 27124
rect 10692 27081 10701 27115
rect 10701 27081 10735 27115
rect 10735 27081 10744 27115
rect 10692 27072 10744 27081
rect 10876 27072 10928 27124
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 14924 27072 14976 27124
rect 17224 27115 17276 27124
rect 17224 27081 17233 27115
rect 17233 27081 17267 27115
rect 17267 27081 17276 27115
rect 17224 27072 17276 27081
rect 18052 27072 18104 27124
rect 18328 27072 18380 27124
rect 21272 27072 21324 27124
rect 21364 27072 21416 27124
rect 23112 27072 23164 27124
rect 26240 27115 26292 27124
rect 26240 27081 26249 27115
rect 26249 27081 26283 27115
rect 26283 27081 26292 27115
rect 26240 27072 26292 27081
rect 27988 27072 28040 27124
rect 28264 27072 28316 27124
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 12532 27004 12584 27056
rect 16488 27004 16540 27056
rect 10968 26936 11020 26988
rect 11704 26936 11756 26988
rect 14740 26936 14792 26988
rect 10232 26868 10284 26920
rect 10876 26911 10928 26920
rect 10876 26877 10885 26911
rect 10885 26877 10919 26911
rect 10919 26877 10928 26911
rect 10876 26868 10928 26877
rect 13452 26868 13504 26920
rect 16948 26936 17000 26988
rect 17040 26868 17092 26920
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 17408 26911 17460 26920
rect 17408 26877 17417 26911
rect 17417 26877 17451 26911
rect 17451 26877 17460 26911
rect 17408 26868 17460 26877
rect 8392 26800 8444 26852
rect 9680 26732 9732 26784
rect 17684 26800 17736 26852
rect 18420 26936 18472 26988
rect 20812 26936 20864 26988
rect 21088 26979 21140 26988
rect 21088 26945 21097 26979
rect 21097 26945 21131 26979
rect 21131 26945 21140 26979
rect 21088 26936 21140 26945
rect 21180 26979 21232 26988
rect 21180 26945 21189 26979
rect 21189 26945 21223 26979
rect 21223 26945 21232 26979
rect 21180 26936 21232 26945
rect 21272 26936 21324 26988
rect 21640 26936 21692 26988
rect 22928 26936 22980 26988
rect 24032 27004 24084 27056
rect 27252 27004 27304 27056
rect 30564 27072 30616 27124
rect 31024 27072 31076 27124
rect 23572 26979 23624 26988
rect 23572 26945 23581 26979
rect 23581 26945 23615 26979
rect 23615 26945 23624 26979
rect 23572 26936 23624 26945
rect 23756 26936 23808 26988
rect 24860 26936 24912 26988
rect 12256 26732 12308 26784
rect 13084 26732 13136 26784
rect 16580 26732 16632 26784
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 17408 26732 17460 26784
rect 21180 26800 21232 26852
rect 21456 26800 21508 26852
rect 18052 26775 18104 26784
rect 18052 26741 18061 26775
rect 18061 26741 18095 26775
rect 18095 26741 18104 26775
rect 18052 26732 18104 26741
rect 18972 26732 19024 26784
rect 19340 26732 19392 26784
rect 19616 26775 19668 26784
rect 19616 26741 19625 26775
rect 19625 26741 19659 26775
rect 19659 26741 19668 26775
rect 19616 26732 19668 26741
rect 20076 26732 20128 26784
rect 20168 26732 20220 26784
rect 23204 26868 23256 26920
rect 24216 26868 24268 26920
rect 25228 26911 25280 26920
rect 25228 26877 25237 26911
rect 25237 26877 25271 26911
rect 25271 26877 25280 26911
rect 25228 26868 25280 26877
rect 25964 26936 26016 26988
rect 30472 27004 30524 27056
rect 30656 27004 30708 27056
rect 31668 27072 31720 27124
rect 28540 26979 28592 26988
rect 28540 26945 28549 26979
rect 28549 26945 28583 26979
rect 28583 26945 28592 26979
rect 28540 26936 28592 26945
rect 28816 26979 28868 26988
rect 28816 26945 28825 26979
rect 28825 26945 28859 26979
rect 28859 26945 28868 26979
rect 28816 26936 28868 26945
rect 29368 26979 29420 26988
rect 29368 26945 29377 26979
rect 29377 26945 29411 26979
rect 29411 26945 29420 26979
rect 29368 26936 29420 26945
rect 29460 26979 29512 26988
rect 29460 26945 29469 26979
rect 29469 26945 29503 26979
rect 29503 26945 29512 26979
rect 29460 26936 29512 26945
rect 29828 26936 29880 26988
rect 26792 26868 26844 26920
rect 28908 26868 28960 26920
rect 30840 26979 30892 26988
rect 30840 26945 30849 26979
rect 30849 26945 30883 26979
rect 30883 26945 30892 26979
rect 30840 26936 30892 26945
rect 30932 26979 30984 26988
rect 30932 26945 30941 26979
rect 30941 26945 30975 26979
rect 30975 26945 30984 26979
rect 30932 26936 30984 26945
rect 31852 26936 31904 26988
rect 32496 26936 32548 26988
rect 33140 26936 33192 26988
rect 31484 26868 31536 26920
rect 31944 26868 31996 26920
rect 34152 26979 34204 26988
rect 34152 26945 34161 26979
rect 34161 26945 34195 26979
rect 34195 26945 34204 26979
rect 34152 26936 34204 26945
rect 34244 26936 34296 26988
rect 34796 26936 34848 26988
rect 34980 27072 35032 27124
rect 35900 27004 35952 27056
rect 36728 27047 36780 27056
rect 36728 27013 36737 27047
rect 36737 27013 36771 27047
rect 36771 27013 36780 27047
rect 36728 27004 36780 27013
rect 37096 27004 37148 27056
rect 37740 27004 37792 27056
rect 37924 26936 37976 26988
rect 38660 26936 38712 26988
rect 39028 26979 39080 26988
rect 39028 26945 39035 26979
rect 39035 26945 39080 26979
rect 39028 26936 39080 26945
rect 39120 26979 39172 26988
rect 39120 26945 39129 26979
rect 39129 26945 39163 26979
rect 39163 26945 39172 26979
rect 39120 26936 39172 26945
rect 36176 26868 36228 26920
rect 22744 26800 22796 26852
rect 23388 26732 23440 26784
rect 24676 26732 24728 26784
rect 26240 26732 26292 26784
rect 26884 26800 26936 26852
rect 33784 26800 33836 26852
rect 36912 26868 36964 26920
rect 38200 26911 38252 26920
rect 38200 26877 38209 26911
rect 38209 26877 38243 26911
rect 38243 26877 38252 26911
rect 38200 26868 38252 26877
rect 32956 26732 33008 26784
rect 33416 26732 33468 26784
rect 36820 26800 36872 26852
rect 37004 26800 37056 26852
rect 37740 26800 37792 26852
rect 40776 26936 40828 26988
rect 41972 26936 42024 26988
rect 42984 26979 43036 26988
rect 42984 26945 42993 26979
rect 42993 26945 43027 26979
rect 43027 26945 43036 26979
rect 42984 26936 43036 26945
rect 43076 26911 43128 26920
rect 43076 26877 43085 26911
rect 43085 26877 43119 26911
rect 43119 26877 43128 26911
rect 43076 26868 43128 26877
rect 43260 26911 43312 26920
rect 43260 26877 43269 26911
rect 43269 26877 43303 26911
rect 43303 26877 43312 26911
rect 43260 26868 43312 26877
rect 39488 26775 39540 26784
rect 39488 26741 39497 26775
rect 39497 26741 39531 26775
rect 39531 26741 39540 26775
rect 39488 26732 39540 26741
rect 40040 26732 40092 26784
rect 42616 26775 42668 26784
rect 42616 26741 42625 26775
rect 42625 26741 42659 26775
rect 42659 26741 42668 26775
rect 42616 26732 42668 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 12164 26571 12216 26580
rect 12164 26537 12173 26571
rect 12173 26537 12207 26571
rect 12207 26537 12216 26571
rect 12164 26528 12216 26537
rect 12256 26528 12308 26580
rect 17408 26528 17460 26580
rect 17500 26528 17552 26580
rect 9036 26460 9088 26512
rect 10968 26435 11020 26444
rect 10968 26401 10977 26435
rect 10977 26401 11011 26435
rect 11011 26401 11020 26435
rect 10968 26392 11020 26401
rect 8116 26324 8168 26376
rect 9496 26367 9548 26376
rect 9496 26333 9505 26367
rect 9505 26333 9539 26367
rect 9539 26333 9548 26367
rect 9496 26324 9548 26333
rect 9680 26367 9732 26376
rect 9680 26333 9689 26367
rect 9689 26333 9723 26367
rect 9723 26333 9732 26367
rect 9680 26324 9732 26333
rect 13268 26460 13320 26512
rect 12440 26392 12492 26444
rect 12716 26367 12768 26376
rect 12716 26333 12725 26367
rect 12725 26333 12759 26367
rect 12759 26333 12768 26367
rect 12716 26324 12768 26333
rect 18328 26503 18380 26512
rect 18328 26469 18337 26503
rect 18337 26469 18371 26503
rect 18371 26469 18380 26503
rect 18328 26460 18380 26469
rect 16948 26435 17000 26444
rect 16948 26401 16957 26435
rect 16957 26401 16991 26435
rect 16991 26401 17000 26435
rect 16948 26392 17000 26401
rect 17040 26392 17092 26444
rect 19340 26392 19392 26444
rect 15200 26324 15252 26376
rect 15752 26367 15804 26376
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 13084 26256 13136 26308
rect 15844 26256 15896 26308
rect 17316 26256 17368 26308
rect 17684 26324 17736 26376
rect 18788 26324 18840 26376
rect 12624 26188 12676 26240
rect 17868 26256 17920 26308
rect 18328 26256 18380 26308
rect 18696 26256 18748 26308
rect 18144 26188 18196 26240
rect 20628 26324 20680 26376
rect 19524 26256 19576 26308
rect 20076 26188 20128 26240
rect 20444 26188 20496 26240
rect 23020 26392 23072 26444
rect 25596 26460 25648 26512
rect 28080 26528 28132 26580
rect 34612 26528 34664 26580
rect 35532 26528 35584 26580
rect 37188 26528 37240 26580
rect 40776 26571 40828 26580
rect 40776 26537 40785 26571
rect 40785 26537 40819 26571
rect 40819 26537 40828 26571
rect 40776 26528 40828 26537
rect 42984 26528 43036 26580
rect 26884 26392 26936 26444
rect 28080 26392 28132 26444
rect 30012 26460 30064 26512
rect 31300 26460 31352 26512
rect 34244 26460 34296 26512
rect 35808 26460 35860 26512
rect 38200 26460 38252 26512
rect 30196 26392 30248 26444
rect 35992 26392 36044 26444
rect 21548 26324 21600 26376
rect 23204 26324 23256 26376
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 26792 26324 26844 26376
rect 26976 26324 27028 26376
rect 22928 26231 22980 26240
rect 22928 26197 22937 26231
rect 22937 26197 22971 26231
rect 22971 26197 22980 26231
rect 22928 26188 22980 26197
rect 27436 26324 27488 26376
rect 27896 26188 27948 26240
rect 28908 26324 28960 26376
rect 29736 26367 29788 26376
rect 29736 26333 29745 26367
rect 29745 26333 29779 26367
rect 29779 26333 29788 26367
rect 29736 26324 29788 26333
rect 29828 26324 29880 26376
rect 31208 26367 31260 26376
rect 31208 26333 31217 26367
rect 31217 26333 31251 26367
rect 31251 26333 31260 26367
rect 31208 26324 31260 26333
rect 31484 26367 31536 26376
rect 31484 26333 31493 26367
rect 31493 26333 31527 26367
rect 31527 26333 31536 26367
rect 32772 26367 32824 26376
rect 31484 26324 31536 26333
rect 28540 26256 28592 26308
rect 28632 26231 28684 26240
rect 28632 26197 28641 26231
rect 28641 26197 28675 26231
rect 28675 26197 28684 26231
rect 28632 26188 28684 26197
rect 30288 26256 30340 26308
rect 31116 26256 31168 26308
rect 31576 26256 31628 26308
rect 32772 26333 32776 26367
rect 32776 26333 32810 26367
rect 32810 26333 32824 26367
rect 32772 26324 32824 26333
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 32864 26324 32916 26333
rect 33232 26367 33284 26376
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33232 26324 33284 26333
rect 33784 26367 33836 26376
rect 33784 26333 33793 26367
rect 33793 26333 33827 26367
rect 33827 26333 33836 26367
rect 33784 26324 33836 26333
rect 33968 26367 34020 26376
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 34244 26324 34296 26376
rect 34428 26324 34480 26376
rect 35164 26367 35216 26376
rect 35164 26333 35173 26367
rect 35173 26333 35207 26367
rect 35207 26333 35216 26367
rect 35164 26324 35216 26333
rect 36452 26324 36504 26376
rect 36636 26367 36688 26376
rect 36636 26333 36645 26367
rect 36645 26333 36679 26367
rect 36679 26333 36688 26367
rect 36636 26324 36688 26333
rect 36728 26367 36780 26376
rect 36728 26333 36737 26367
rect 36737 26333 36771 26367
rect 36771 26333 36780 26367
rect 36728 26324 36780 26333
rect 30932 26188 30984 26240
rect 33508 26256 33560 26308
rect 34060 26299 34112 26308
rect 34060 26265 34069 26299
rect 34069 26265 34103 26299
rect 34103 26265 34112 26299
rect 34060 26256 34112 26265
rect 36176 26256 36228 26308
rect 37004 26367 37056 26376
rect 37004 26333 37013 26367
rect 37013 26333 37047 26367
rect 37047 26333 37056 26367
rect 37004 26324 37056 26333
rect 37556 26367 37608 26376
rect 37556 26333 37565 26367
rect 37565 26333 37599 26367
rect 37599 26333 37608 26367
rect 37556 26324 37608 26333
rect 37740 26324 37792 26376
rect 37832 26324 37884 26376
rect 33140 26188 33192 26240
rect 38660 26367 38712 26376
rect 38660 26333 38669 26367
rect 38669 26333 38703 26367
rect 38703 26333 38712 26367
rect 38660 26324 38712 26333
rect 39672 26392 39724 26444
rect 40316 26435 40368 26444
rect 40316 26401 40325 26435
rect 40325 26401 40359 26435
rect 40359 26401 40368 26435
rect 40316 26392 40368 26401
rect 41972 26435 42024 26444
rect 41972 26401 41981 26435
rect 41981 26401 42015 26435
rect 42015 26401 42024 26435
rect 41972 26392 42024 26401
rect 39304 26324 39356 26376
rect 40684 26324 40736 26376
rect 42616 26324 42668 26376
rect 35164 26188 35216 26240
rect 35532 26188 35584 26240
rect 36268 26188 36320 26240
rect 36452 26188 36504 26240
rect 36544 26188 36596 26240
rect 38936 26299 38988 26308
rect 38936 26265 38945 26299
rect 38945 26265 38979 26299
rect 38979 26265 38988 26299
rect 38936 26256 38988 26265
rect 39028 26299 39080 26308
rect 39028 26265 39037 26299
rect 39037 26265 39071 26299
rect 39071 26265 39080 26299
rect 39028 26256 39080 26265
rect 38844 26188 38896 26240
rect 39120 26188 39172 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 15844 26027 15896 26036
rect 15844 25993 15853 26027
rect 15853 25993 15887 26027
rect 15887 25993 15896 26027
rect 15844 25984 15896 25993
rect 19432 25984 19484 26036
rect 21272 25984 21324 26036
rect 12624 25959 12676 25968
rect 12624 25925 12633 25959
rect 12633 25925 12667 25959
rect 12667 25925 12676 25959
rect 12624 25916 12676 25925
rect 17500 25916 17552 25968
rect 18144 25959 18196 25968
rect 18144 25925 18153 25959
rect 18153 25925 18187 25959
rect 18187 25925 18196 25959
rect 18144 25916 18196 25925
rect 20076 25916 20128 25968
rect 22928 25916 22980 25968
rect 23204 25916 23256 25968
rect 23940 25916 23992 25968
rect 15200 25848 15252 25900
rect 19984 25891 20036 25900
rect 19984 25857 19993 25891
rect 19993 25857 20027 25891
rect 20027 25857 20036 25891
rect 19984 25848 20036 25857
rect 20168 25891 20220 25900
rect 20168 25857 20177 25891
rect 20177 25857 20211 25891
rect 20211 25857 20220 25891
rect 20168 25848 20220 25857
rect 22560 25891 22612 25900
rect 22560 25857 22569 25891
rect 22569 25857 22603 25891
rect 22603 25857 22612 25891
rect 22560 25848 22612 25857
rect 11888 25823 11940 25832
rect 11888 25789 11897 25823
rect 11897 25789 11931 25823
rect 11931 25789 11940 25823
rect 11888 25780 11940 25789
rect 16856 25780 16908 25832
rect 18972 25823 19024 25832
rect 18972 25789 18981 25823
rect 18981 25789 19015 25823
rect 19015 25789 19024 25823
rect 18972 25780 19024 25789
rect 19064 25823 19116 25832
rect 19064 25789 19073 25823
rect 19073 25789 19107 25823
rect 19107 25789 19116 25823
rect 19064 25780 19116 25789
rect 20076 25780 20128 25832
rect 24952 25848 25004 25900
rect 27252 26027 27304 26036
rect 27252 25993 27261 26027
rect 27261 25993 27295 26027
rect 27295 25993 27304 26027
rect 27252 25984 27304 25993
rect 28816 25984 28868 26036
rect 28908 25984 28960 26036
rect 32956 25984 33008 26036
rect 30748 25959 30800 25968
rect 30748 25925 30757 25959
rect 30757 25925 30791 25959
rect 30791 25925 30800 25959
rect 30748 25916 30800 25925
rect 26424 25891 26476 25900
rect 26424 25857 26433 25891
rect 26433 25857 26467 25891
rect 26467 25857 26476 25891
rect 26424 25848 26476 25857
rect 26516 25848 26568 25900
rect 27712 25848 27764 25900
rect 27252 25780 27304 25832
rect 17868 25712 17920 25764
rect 18236 25712 18288 25764
rect 20352 25687 20404 25696
rect 20352 25653 20361 25687
rect 20361 25653 20395 25687
rect 20395 25653 20404 25687
rect 20352 25644 20404 25653
rect 23940 25687 23992 25696
rect 23940 25653 23949 25687
rect 23949 25653 23983 25687
rect 23983 25653 23992 25687
rect 23940 25644 23992 25653
rect 24768 25644 24820 25696
rect 26884 25712 26936 25764
rect 30656 25848 30708 25900
rect 28080 25823 28132 25832
rect 28080 25789 28089 25823
rect 28089 25789 28123 25823
rect 28123 25789 28132 25823
rect 28080 25780 28132 25789
rect 31300 25916 31352 25968
rect 32680 25916 32732 25968
rect 33048 25959 33100 25968
rect 33048 25925 33057 25959
rect 33057 25925 33091 25959
rect 33091 25925 33100 25959
rect 33048 25916 33100 25925
rect 33140 25959 33192 25968
rect 33140 25925 33149 25959
rect 33149 25925 33183 25959
rect 33183 25925 33192 25959
rect 33140 25916 33192 25925
rect 31208 25848 31260 25900
rect 31392 25848 31444 25900
rect 32772 25848 32824 25900
rect 36452 25984 36504 26036
rect 36544 25984 36596 26036
rect 40040 26027 40092 26036
rect 35992 25916 36044 25968
rect 33416 25891 33468 25900
rect 33416 25857 33425 25891
rect 33425 25857 33459 25891
rect 33459 25857 33468 25891
rect 33416 25848 33468 25857
rect 34428 25848 34480 25900
rect 34796 25848 34848 25900
rect 35808 25848 35860 25900
rect 37004 25848 37056 25900
rect 38660 25848 38712 25900
rect 40040 25993 40049 26027
rect 40049 25993 40083 26027
rect 40083 25993 40092 26027
rect 40040 25984 40092 25993
rect 39488 25916 39540 25968
rect 43168 25959 43220 25968
rect 43168 25925 43177 25959
rect 43177 25925 43211 25959
rect 43211 25925 43220 25959
rect 43168 25916 43220 25925
rect 38844 25848 38896 25900
rect 39120 25891 39172 25900
rect 39120 25857 39129 25891
rect 39129 25857 39163 25891
rect 39163 25857 39172 25891
rect 39120 25848 39172 25857
rect 40132 25891 40184 25900
rect 40132 25857 40141 25891
rect 40141 25857 40175 25891
rect 40175 25857 40184 25891
rect 40132 25848 40184 25857
rect 41144 25848 41196 25900
rect 35624 25780 35676 25832
rect 37464 25780 37516 25832
rect 43076 25848 43128 25900
rect 36268 25755 36320 25764
rect 36268 25721 36277 25755
rect 36277 25721 36311 25755
rect 36311 25721 36320 25755
rect 36268 25712 36320 25721
rect 27896 25644 27948 25696
rect 31024 25644 31076 25696
rect 31944 25644 31996 25696
rect 34060 25644 34112 25696
rect 38568 25712 38620 25764
rect 40316 25712 40368 25764
rect 36820 25687 36872 25696
rect 36820 25653 36829 25687
rect 36829 25653 36863 25687
rect 36863 25653 36872 25687
rect 36820 25644 36872 25653
rect 39028 25644 39080 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10600 25440 10652 25492
rect 10876 25372 10928 25424
rect 18604 25440 18656 25492
rect 19064 25440 19116 25492
rect 19984 25440 20036 25492
rect 21548 25440 21600 25492
rect 24492 25440 24544 25492
rect 27712 25440 27764 25492
rect 31392 25440 31444 25492
rect 32220 25440 32272 25492
rect 33232 25440 33284 25492
rect 36176 25440 36228 25492
rect 40684 25483 40736 25492
rect 40684 25449 40693 25483
rect 40693 25449 40727 25483
rect 40727 25449 40736 25483
rect 40684 25440 40736 25449
rect 20076 25372 20128 25424
rect 22192 25372 22244 25424
rect 30840 25372 30892 25424
rect 31300 25372 31352 25424
rect 31760 25372 31812 25424
rect 31852 25415 31904 25424
rect 31852 25381 31861 25415
rect 31861 25381 31895 25415
rect 31895 25381 31904 25415
rect 31852 25372 31904 25381
rect 10968 25236 11020 25288
rect 10232 25168 10284 25220
rect 10692 25168 10744 25220
rect 12716 25236 12768 25288
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 13912 25236 13964 25288
rect 14372 25236 14424 25288
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 15200 25279 15252 25288
rect 15200 25245 15209 25279
rect 15209 25245 15243 25279
rect 15243 25245 15252 25279
rect 15200 25236 15252 25245
rect 17040 25236 17092 25288
rect 11704 25143 11756 25152
rect 11704 25109 11713 25143
rect 11713 25109 11747 25143
rect 11747 25109 11756 25143
rect 11704 25100 11756 25109
rect 13360 25168 13412 25220
rect 12808 25143 12860 25152
rect 12808 25109 12817 25143
rect 12817 25109 12851 25143
rect 12851 25109 12860 25143
rect 12808 25100 12860 25109
rect 14740 25100 14792 25152
rect 15108 25168 15160 25220
rect 17316 25236 17368 25288
rect 15844 25100 15896 25152
rect 17776 25168 17828 25220
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 20628 25347 20680 25356
rect 20628 25313 20637 25347
rect 20637 25313 20671 25347
rect 20671 25313 20680 25347
rect 20628 25304 20680 25313
rect 28172 25304 28224 25356
rect 31944 25304 31996 25356
rect 20352 25236 20404 25288
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 25872 25236 25924 25288
rect 27068 25279 27120 25288
rect 27068 25245 27117 25279
rect 27117 25245 27120 25279
rect 27068 25236 27120 25245
rect 27344 25279 27396 25288
rect 27344 25245 27353 25279
rect 27353 25245 27387 25279
rect 27387 25245 27396 25279
rect 27344 25236 27396 25245
rect 27896 25236 27948 25288
rect 18788 25168 18840 25220
rect 23296 25168 23348 25220
rect 26884 25168 26936 25220
rect 28172 25168 28224 25220
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 30564 25236 30616 25288
rect 30932 25279 30984 25288
rect 30932 25245 30941 25279
rect 30941 25245 30975 25279
rect 30975 25245 30984 25279
rect 30932 25236 30984 25245
rect 31300 25236 31352 25288
rect 31484 25236 31536 25288
rect 32312 25236 32364 25288
rect 32496 25236 32548 25288
rect 34244 25304 34296 25356
rect 35440 25279 35492 25288
rect 35440 25245 35449 25279
rect 35449 25245 35483 25279
rect 35483 25245 35492 25279
rect 35440 25236 35492 25245
rect 35624 25279 35676 25288
rect 35624 25245 35631 25279
rect 35631 25245 35676 25279
rect 35624 25236 35676 25245
rect 39028 25347 39080 25356
rect 39028 25313 39037 25347
rect 39037 25313 39071 25347
rect 39071 25313 39080 25347
rect 39028 25304 39080 25313
rect 40224 25304 40276 25356
rect 30104 25168 30156 25220
rect 30472 25168 30524 25220
rect 32772 25168 32824 25220
rect 35716 25211 35768 25220
rect 35716 25177 35725 25211
rect 35725 25177 35759 25211
rect 35759 25177 35768 25211
rect 35716 25168 35768 25177
rect 35808 25211 35860 25220
rect 35808 25177 35817 25211
rect 35817 25177 35851 25211
rect 35851 25177 35860 25211
rect 35808 25168 35860 25177
rect 18052 25100 18104 25152
rect 26976 25100 27028 25152
rect 29276 25100 29328 25152
rect 30288 25100 30340 25152
rect 31392 25100 31444 25152
rect 36728 25236 36780 25288
rect 36912 25236 36964 25288
rect 37648 25279 37700 25288
rect 37648 25245 37657 25279
rect 37657 25245 37691 25279
rect 37691 25245 37700 25279
rect 37648 25236 37700 25245
rect 38936 25279 38988 25288
rect 38936 25245 38945 25279
rect 38945 25245 38979 25279
rect 38979 25245 38988 25279
rect 38936 25236 38988 25245
rect 39212 25279 39264 25288
rect 39212 25245 39221 25279
rect 39221 25245 39255 25279
rect 39255 25245 39264 25279
rect 39212 25236 39264 25245
rect 39304 25279 39356 25288
rect 39304 25245 39313 25279
rect 39313 25245 39347 25279
rect 39347 25245 39356 25279
rect 39304 25236 39356 25245
rect 43076 25236 43128 25288
rect 40316 25211 40368 25220
rect 40316 25177 40325 25211
rect 40325 25177 40359 25211
rect 40359 25177 40368 25211
rect 40316 25168 40368 25177
rect 40408 25168 40460 25220
rect 43996 25168 44048 25220
rect 36912 25143 36964 25152
rect 36912 25109 36921 25143
rect 36921 25109 36955 25143
rect 36955 25109 36964 25143
rect 36912 25100 36964 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 10232 24939 10284 24948
rect 10232 24905 10241 24939
rect 10241 24905 10275 24939
rect 10275 24905 10284 24939
rect 10232 24896 10284 24905
rect 10600 24939 10652 24948
rect 10600 24905 10609 24939
rect 10609 24905 10643 24939
rect 10643 24905 10652 24939
rect 10600 24896 10652 24905
rect 17316 24896 17368 24948
rect 25688 24896 25740 24948
rect 25872 24896 25924 24948
rect 12808 24871 12860 24880
rect 12808 24837 12842 24871
rect 12842 24837 12860 24871
rect 12808 24828 12860 24837
rect 17500 24828 17552 24880
rect 9036 24803 9088 24812
rect 9036 24769 9054 24803
rect 9054 24769 9088 24803
rect 9036 24760 9088 24769
rect 10692 24803 10744 24812
rect 10692 24769 10701 24803
rect 10701 24769 10735 24803
rect 10735 24769 10744 24803
rect 10692 24760 10744 24769
rect 14740 24803 14792 24812
rect 14740 24769 14774 24803
rect 14774 24769 14792 24803
rect 14740 24760 14792 24769
rect 21088 24760 21140 24812
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 10876 24735 10928 24744
rect 10876 24701 10885 24735
rect 10885 24701 10919 24735
rect 10919 24701 10928 24735
rect 10876 24692 10928 24701
rect 11888 24692 11940 24744
rect 11060 24624 11112 24676
rect 8300 24556 8352 24608
rect 13912 24599 13964 24608
rect 13912 24565 13921 24599
rect 13921 24565 13955 24599
rect 13955 24565 13964 24599
rect 13912 24556 13964 24565
rect 16856 24692 16908 24744
rect 24952 24828 25004 24880
rect 28540 24896 28592 24948
rect 33508 24896 33560 24948
rect 35808 24896 35860 24948
rect 38936 24896 38988 24948
rect 39304 24896 39356 24948
rect 43076 24939 43128 24948
rect 43076 24905 43085 24939
rect 43085 24905 43119 24939
rect 43119 24905 43128 24939
rect 43076 24896 43128 24905
rect 15752 24624 15804 24676
rect 22744 24692 22796 24744
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 23480 24692 23532 24744
rect 15844 24599 15896 24608
rect 15844 24565 15853 24599
rect 15853 24565 15887 24599
rect 15887 24565 15896 24599
rect 22836 24624 22888 24676
rect 24860 24692 24912 24744
rect 25412 24760 25464 24812
rect 31392 24828 31444 24880
rect 32680 24871 32732 24880
rect 32680 24837 32689 24871
rect 32689 24837 32723 24871
rect 32723 24837 32732 24871
rect 32680 24828 32732 24837
rect 35716 24828 35768 24880
rect 28356 24760 28408 24812
rect 29460 24760 29512 24812
rect 15844 24556 15896 24565
rect 19340 24556 19392 24608
rect 22376 24556 22428 24608
rect 27712 24624 27764 24676
rect 23848 24556 23900 24608
rect 29276 24735 29328 24744
rect 29276 24701 29285 24735
rect 29285 24701 29319 24735
rect 29319 24701 29328 24735
rect 29276 24692 29328 24701
rect 30104 24760 30156 24812
rect 30564 24760 30616 24812
rect 30748 24803 30800 24812
rect 30748 24769 30757 24803
rect 30757 24769 30791 24803
rect 30791 24769 30800 24803
rect 30748 24760 30800 24769
rect 30840 24803 30892 24812
rect 30840 24769 30869 24803
rect 30869 24769 30892 24803
rect 30840 24760 30892 24769
rect 31760 24760 31812 24812
rect 29736 24735 29788 24744
rect 29736 24701 29745 24735
rect 29745 24701 29779 24735
rect 29779 24701 29788 24735
rect 29736 24692 29788 24701
rect 30472 24735 30524 24744
rect 30472 24701 30481 24735
rect 30481 24701 30515 24735
rect 30515 24701 30524 24735
rect 30472 24692 30524 24701
rect 32220 24692 32272 24744
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 35992 24760 36044 24812
rect 30656 24624 30708 24676
rect 31576 24624 31628 24676
rect 36268 24624 36320 24676
rect 30840 24556 30892 24608
rect 31024 24599 31076 24608
rect 31024 24565 31033 24599
rect 31033 24565 31067 24599
rect 31067 24565 31076 24599
rect 31024 24556 31076 24565
rect 32588 24556 32640 24608
rect 35900 24556 35952 24608
rect 38568 24803 38620 24812
rect 38568 24769 38577 24803
rect 38577 24769 38611 24803
rect 38611 24769 38620 24803
rect 38568 24760 38620 24769
rect 38016 24692 38068 24744
rect 36728 24556 36780 24608
rect 38660 24556 38712 24608
rect 38844 24803 38896 24812
rect 38844 24769 38853 24803
rect 38853 24769 38887 24803
rect 38887 24769 38896 24803
rect 38844 24760 38896 24769
rect 38936 24803 38988 24812
rect 38936 24769 38945 24803
rect 38945 24769 38979 24803
rect 38979 24769 38988 24803
rect 38936 24760 38988 24769
rect 39396 24760 39448 24812
rect 39488 24760 39540 24812
rect 39948 24803 40000 24812
rect 39948 24769 39957 24803
rect 39957 24769 39991 24803
rect 39991 24769 40000 24803
rect 39948 24760 40000 24769
rect 40132 24760 40184 24812
rect 40776 24760 40828 24812
rect 41972 24760 42024 24812
rect 42984 24803 43036 24812
rect 42984 24769 42993 24803
rect 42993 24769 43027 24803
rect 43027 24769 43036 24803
rect 42984 24760 43036 24769
rect 39120 24624 39172 24676
rect 40316 24624 40368 24676
rect 39764 24556 39816 24608
rect 43260 24735 43312 24744
rect 43260 24701 43269 24735
rect 43269 24701 43303 24735
rect 43303 24701 43312 24735
rect 43260 24692 43312 24701
rect 42616 24599 42668 24608
rect 42616 24565 42625 24599
rect 42625 24565 42659 24599
rect 42659 24565 42668 24599
rect 42616 24556 42668 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8300 24352 8352 24404
rect 9404 24352 9456 24404
rect 10140 24216 10192 24268
rect 10876 24216 10928 24268
rect 14556 24352 14608 24404
rect 13912 24284 13964 24336
rect 22468 24352 22520 24404
rect 22836 24352 22888 24404
rect 27252 24352 27304 24404
rect 28080 24352 28132 24404
rect 30104 24352 30156 24404
rect 30748 24352 30800 24404
rect 39212 24352 39264 24404
rect 39488 24395 39540 24404
rect 39488 24361 39497 24395
rect 39497 24361 39531 24395
rect 39531 24361 39540 24395
rect 39488 24352 39540 24361
rect 40776 24395 40828 24404
rect 40776 24361 40785 24395
rect 40785 24361 40819 24395
rect 40819 24361 40828 24395
rect 40776 24352 40828 24361
rect 15384 24216 15436 24268
rect 11060 24148 11112 24200
rect 11888 24148 11940 24200
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 16856 24148 16908 24200
rect 11704 24080 11756 24132
rect 9864 24055 9916 24064
rect 9864 24021 9873 24055
rect 9873 24021 9907 24055
rect 9907 24021 9916 24055
rect 9864 24012 9916 24021
rect 10232 24055 10284 24064
rect 10232 24021 10241 24055
rect 10241 24021 10275 24055
rect 10275 24021 10284 24055
rect 10232 24012 10284 24021
rect 12716 24055 12768 24064
rect 12716 24021 12725 24055
rect 12725 24021 12759 24055
rect 12759 24021 12768 24055
rect 19984 24216 20036 24268
rect 21088 24284 21140 24336
rect 22008 24284 22060 24336
rect 25320 24284 25372 24336
rect 20168 24216 20220 24268
rect 20536 24148 20588 24200
rect 22376 24148 22428 24200
rect 22744 24148 22796 24200
rect 23756 24216 23808 24268
rect 23480 24191 23532 24200
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 27068 24191 27120 24200
rect 27068 24157 27072 24191
rect 27072 24157 27106 24191
rect 27106 24157 27120 24191
rect 24492 24080 24544 24132
rect 27068 24148 27120 24157
rect 35808 24284 35860 24336
rect 38936 24284 38988 24336
rect 42984 24352 43036 24404
rect 27712 24216 27764 24268
rect 29184 24216 29236 24268
rect 29736 24216 29788 24268
rect 31208 24216 31260 24268
rect 27344 24148 27396 24200
rect 27528 24148 27580 24200
rect 28264 24148 28316 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 28540 24148 28592 24200
rect 28908 24148 28960 24200
rect 12716 24012 12768 24021
rect 19432 24012 19484 24064
rect 21088 24012 21140 24064
rect 22468 24012 22520 24064
rect 24676 24055 24728 24064
rect 24676 24021 24685 24055
rect 24685 24021 24719 24055
rect 24719 24021 24728 24055
rect 24676 24012 24728 24021
rect 27712 24080 27764 24132
rect 28632 24012 28684 24064
rect 30104 24191 30156 24200
rect 30104 24157 30113 24191
rect 30113 24157 30147 24191
rect 30147 24157 30156 24191
rect 30104 24148 30156 24157
rect 34428 24216 34480 24268
rect 37556 24259 37608 24268
rect 37556 24225 37565 24259
rect 37565 24225 37599 24259
rect 37599 24225 37608 24259
rect 37556 24216 37608 24225
rect 37648 24216 37700 24268
rect 38016 24259 38068 24268
rect 38016 24225 38025 24259
rect 38025 24225 38059 24259
rect 38059 24225 38068 24259
rect 38016 24216 38068 24225
rect 33048 24148 33100 24200
rect 30288 24080 30340 24132
rect 30932 24123 30984 24132
rect 30932 24089 30941 24123
rect 30941 24089 30975 24123
rect 30975 24089 30984 24123
rect 30932 24080 30984 24089
rect 30472 24012 30524 24064
rect 30840 24012 30892 24064
rect 32956 24080 33008 24132
rect 35348 24148 35400 24200
rect 37832 24148 37884 24200
rect 38844 24191 38896 24200
rect 38844 24157 38853 24191
rect 38853 24157 38887 24191
rect 38887 24157 38896 24191
rect 38844 24148 38896 24157
rect 40316 24259 40368 24268
rect 40316 24225 40325 24259
rect 40325 24225 40359 24259
rect 40359 24225 40368 24259
rect 40316 24216 40368 24225
rect 41972 24259 42024 24268
rect 41972 24225 41981 24259
rect 41981 24225 42015 24259
rect 42015 24225 42024 24259
rect 41972 24216 42024 24225
rect 39028 24148 39080 24200
rect 39580 24148 39632 24200
rect 40408 24191 40460 24200
rect 40408 24157 40417 24191
rect 40417 24157 40451 24191
rect 40451 24157 40460 24191
rect 40408 24148 40460 24157
rect 42616 24148 42668 24200
rect 34612 24080 34664 24132
rect 35532 24080 35584 24132
rect 39212 24123 39264 24132
rect 39212 24089 39218 24123
rect 39218 24089 39252 24123
rect 39252 24089 39264 24123
rect 39212 24080 39264 24089
rect 35256 24012 35308 24064
rect 38660 24012 38712 24064
rect 38936 24012 38988 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 14740 23808 14792 23860
rect 11060 23740 11112 23792
rect 9864 23672 9916 23724
rect 20260 23808 20312 23860
rect 10232 23604 10284 23656
rect 16212 23604 16264 23656
rect 16948 23604 17000 23656
rect 19432 23672 19484 23724
rect 18052 23468 18104 23520
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20536 23672 20588 23724
rect 22008 23740 22060 23792
rect 22468 23783 22520 23792
rect 22468 23749 22477 23783
rect 22477 23749 22511 23783
rect 22511 23749 22520 23783
rect 22468 23740 22520 23749
rect 24400 23851 24452 23860
rect 24400 23817 24409 23851
rect 24409 23817 24443 23851
rect 24443 23817 24452 23851
rect 24400 23808 24452 23817
rect 24584 23808 24636 23860
rect 26976 23808 27028 23860
rect 28080 23851 28132 23860
rect 28080 23817 28089 23851
rect 28089 23817 28123 23851
rect 28123 23817 28132 23851
rect 28080 23808 28132 23817
rect 28264 23808 28316 23860
rect 31208 23808 31260 23860
rect 33140 23808 33192 23860
rect 24676 23783 24728 23792
rect 24676 23749 24685 23783
rect 24685 23749 24719 23783
rect 24719 23749 24728 23783
rect 24676 23740 24728 23749
rect 25596 23783 25648 23792
rect 25596 23749 25605 23783
rect 25605 23749 25639 23783
rect 25639 23749 25648 23783
rect 25596 23740 25648 23749
rect 26700 23740 26752 23792
rect 27160 23783 27212 23792
rect 27160 23749 27169 23783
rect 27169 23749 27203 23783
rect 27203 23749 27212 23783
rect 27160 23740 27212 23749
rect 39948 23808 40000 23860
rect 21088 23715 21140 23724
rect 21088 23681 21097 23715
rect 21097 23681 21131 23715
rect 21131 23681 21140 23715
rect 21088 23672 21140 23681
rect 21548 23672 21600 23724
rect 20996 23604 21048 23656
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 35992 23740 36044 23792
rect 27160 23604 27212 23656
rect 28172 23715 28224 23724
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 28080 23604 28132 23656
rect 28908 23715 28960 23724
rect 28908 23681 28917 23715
rect 28917 23681 28951 23715
rect 28951 23681 28960 23715
rect 28908 23672 28960 23681
rect 29184 23672 29236 23724
rect 30472 23672 30524 23724
rect 30564 23672 30616 23724
rect 32588 23715 32640 23724
rect 32588 23681 32597 23715
rect 32597 23681 32631 23715
rect 32631 23681 32640 23715
rect 32588 23672 32640 23681
rect 21180 23536 21232 23588
rect 22192 23579 22244 23588
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 22192 23536 22244 23545
rect 24124 23579 24176 23588
rect 24124 23545 24133 23579
rect 24133 23545 24167 23579
rect 24167 23545 24176 23579
rect 24124 23536 24176 23545
rect 25320 23579 25372 23588
rect 25320 23545 25329 23579
rect 25329 23545 25363 23579
rect 25363 23545 25372 23579
rect 25320 23536 25372 23545
rect 25412 23536 25464 23588
rect 29184 23579 29236 23588
rect 29184 23545 29193 23579
rect 29193 23545 29227 23579
rect 29227 23545 29236 23579
rect 29184 23536 29236 23545
rect 22744 23468 22796 23520
rect 25044 23468 25096 23520
rect 25136 23511 25188 23520
rect 25136 23477 25145 23511
rect 25145 23477 25179 23511
rect 25179 23477 25188 23511
rect 25136 23468 25188 23477
rect 27252 23468 27304 23520
rect 28356 23468 28408 23520
rect 30104 23511 30156 23520
rect 30104 23477 30113 23511
rect 30113 23477 30147 23511
rect 30147 23477 30156 23511
rect 30104 23468 30156 23477
rect 30564 23579 30616 23588
rect 30564 23545 30573 23579
rect 30573 23545 30607 23579
rect 30607 23545 30616 23579
rect 30564 23536 30616 23545
rect 30932 23468 30984 23520
rect 31208 23647 31260 23656
rect 31208 23613 31217 23647
rect 31217 23613 31251 23647
rect 31251 23613 31260 23647
rect 31208 23604 31260 23613
rect 31300 23536 31352 23588
rect 32036 23604 32088 23656
rect 33692 23672 33744 23724
rect 33968 23672 34020 23724
rect 34060 23715 34112 23724
rect 34060 23681 34069 23715
rect 34069 23681 34103 23715
rect 34103 23681 34112 23715
rect 34060 23672 34112 23681
rect 34612 23715 34664 23724
rect 34612 23681 34621 23715
rect 34621 23681 34655 23715
rect 34655 23681 34664 23715
rect 34612 23672 34664 23681
rect 35348 23672 35400 23724
rect 35532 23672 35584 23724
rect 36452 23672 36504 23724
rect 37188 23672 37240 23724
rect 42708 23672 42760 23724
rect 35900 23604 35952 23656
rect 39028 23604 39080 23656
rect 39212 23604 39264 23656
rect 43996 23604 44048 23656
rect 35256 23536 35308 23588
rect 35348 23536 35400 23588
rect 33048 23468 33100 23520
rect 33508 23468 33560 23520
rect 34060 23468 34112 23520
rect 34612 23468 34664 23520
rect 39580 23536 39632 23588
rect 37648 23468 37700 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 10968 23264 11020 23316
rect 17316 23307 17368 23316
rect 17316 23273 17325 23307
rect 17325 23273 17359 23307
rect 17359 23273 17368 23307
rect 17316 23264 17368 23273
rect 10692 23171 10744 23180
rect 10692 23137 10701 23171
rect 10701 23137 10735 23171
rect 10735 23137 10744 23171
rect 10692 23128 10744 23137
rect 16856 23128 16908 23180
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 12256 22992 12308 23044
rect 16764 22992 16816 23044
rect 22468 23264 22520 23316
rect 24308 23264 24360 23316
rect 24768 23264 24820 23316
rect 18788 23196 18840 23248
rect 18696 23060 18748 23112
rect 20444 23128 20496 23180
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 19892 23060 19944 23112
rect 21088 23060 21140 23112
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 26608 23196 26660 23248
rect 23204 23171 23256 23180
rect 23204 23137 23213 23171
rect 23213 23137 23247 23171
rect 23247 23137 23256 23171
rect 23204 23128 23256 23137
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 26976 23128 27028 23180
rect 27436 23171 27488 23180
rect 27436 23137 27445 23171
rect 27445 23137 27479 23171
rect 27479 23137 27488 23171
rect 27436 23128 27488 23137
rect 28172 23128 28224 23180
rect 30288 23264 30340 23316
rect 31760 23264 31812 23316
rect 32496 23264 32548 23316
rect 33048 23264 33100 23316
rect 38200 23264 38252 23316
rect 30104 23196 30156 23248
rect 19248 22992 19300 23044
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 19708 22924 19760 22976
rect 19984 22924 20036 22976
rect 20352 22924 20404 22976
rect 21180 22924 21232 22976
rect 22468 23103 22520 23112
rect 22468 23069 22477 23103
rect 22477 23069 22511 23103
rect 22511 23069 22520 23103
rect 22468 23060 22520 23069
rect 22560 23103 22612 23112
rect 22560 23069 22569 23103
rect 22569 23069 22603 23103
rect 22603 23069 22612 23103
rect 22560 23060 22612 23069
rect 22376 22992 22428 23044
rect 24768 23060 24820 23112
rect 27252 23060 27304 23112
rect 30288 23105 30340 23112
rect 30288 23071 30297 23105
rect 30297 23071 30331 23105
rect 30331 23071 30340 23105
rect 35532 23128 35584 23180
rect 30288 23060 30340 23071
rect 33692 23103 33744 23112
rect 33692 23069 33701 23103
rect 33701 23069 33735 23103
rect 33735 23069 33744 23103
rect 33692 23060 33744 23069
rect 34244 23060 34296 23112
rect 35624 23103 35676 23112
rect 35624 23069 35633 23103
rect 35633 23069 35667 23103
rect 35667 23069 35676 23103
rect 35624 23060 35676 23069
rect 36084 23128 36136 23180
rect 36544 23171 36596 23180
rect 36544 23137 36553 23171
rect 36553 23137 36587 23171
rect 36587 23137 36596 23171
rect 36544 23128 36596 23137
rect 35808 23103 35860 23112
rect 35808 23069 35817 23103
rect 35817 23069 35851 23103
rect 35851 23069 35860 23103
rect 35808 23060 35860 23069
rect 36176 23060 36228 23112
rect 36636 23060 36688 23112
rect 36728 23103 36780 23112
rect 36728 23069 36737 23103
rect 36737 23069 36771 23103
rect 36771 23069 36780 23103
rect 36728 23060 36780 23069
rect 38476 23196 38528 23248
rect 37188 23128 37240 23180
rect 37648 23103 37700 23112
rect 37648 23069 37657 23103
rect 37657 23069 37691 23103
rect 37691 23069 37700 23103
rect 37648 23060 37700 23069
rect 43076 23264 43128 23316
rect 40224 23128 40276 23180
rect 25780 23035 25832 23044
rect 25780 23001 25789 23035
rect 25789 23001 25823 23035
rect 25823 23001 25832 23035
rect 25780 22992 25832 23001
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 24860 22924 24912 22976
rect 25504 22924 25556 22976
rect 28356 22992 28408 23044
rect 30840 22924 30892 22976
rect 33324 22924 33376 22976
rect 34152 22992 34204 23044
rect 38752 23060 38804 23112
rect 39028 23103 39080 23112
rect 39028 23069 39035 23103
rect 39035 23069 39080 23103
rect 39028 23060 39080 23069
rect 39396 23060 39448 23112
rect 40040 23103 40092 23112
rect 40040 23069 40049 23103
rect 40049 23069 40083 23103
rect 40083 23069 40092 23103
rect 40040 23060 40092 23069
rect 40316 23103 40368 23112
rect 40316 23069 40325 23103
rect 40325 23069 40359 23103
rect 40359 23069 40368 23103
rect 40316 23060 40368 23069
rect 42708 23171 42760 23180
rect 42708 23137 42717 23171
rect 42717 23137 42751 23171
rect 42751 23137 42760 23171
rect 42708 23128 42760 23137
rect 43260 23128 43312 23180
rect 39120 23035 39172 23044
rect 39120 23001 39129 23035
rect 39129 23001 39163 23035
rect 39163 23001 39172 23035
rect 39120 22992 39172 23001
rect 34612 22924 34664 22976
rect 37004 22967 37056 22976
rect 37004 22933 37013 22967
rect 37013 22933 37047 22967
rect 37047 22933 37056 22967
rect 37004 22924 37056 22933
rect 39028 22924 39080 22976
rect 42064 22924 42116 22976
rect 43168 22924 43220 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 15108 22720 15160 22772
rect 16948 22763 17000 22772
rect 16948 22729 16957 22763
rect 16957 22729 16991 22763
rect 16991 22729 17000 22763
rect 16948 22720 17000 22729
rect 18880 22720 18932 22772
rect 19156 22720 19208 22772
rect 20536 22720 20588 22772
rect 22560 22720 22612 22772
rect 23480 22720 23532 22772
rect 24400 22720 24452 22772
rect 27988 22720 28040 22772
rect 31392 22720 31444 22772
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 16764 22584 16816 22636
rect 18052 22652 18104 22704
rect 13636 22559 13688 22568
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 18328 22584 18380 22636
rect 22192 22652 22244 22704
rect 25320 22652 25372 22704
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 27068 22584 27120 22636
rect 27712 22627 27764 22636
rect 27712 22593 27721 22627
rect 27721 22593 27755 22627
rect 27755 22593 27764 22627
rect 27712 22584 27764 22593
rect 27896 22627 27948 22636
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 28356 22695 28408 22704
rect 28356 22661 28365 22695
rect 28365 22661 28399 22695
rect 28399 22661 28408 22695
rect 28356 22652 28408 22661
rect 33324 22652 33376 22704
rect 33692 22652 33744 22704
rect 35256 22695 35308 22704
rect 35256 22661 35265 22695
rect 35265 22661 35299 22695
rect 35299 22661 35308 22695
rect 35256 22652 35308 22661
rect 35808 22720 35860 22772
rect 36176 22763 36228 22772
rect 36176 22729 36185 22763
rect 36185 22729 36219 22763
rect 36219 22729 36228 22763
rect 36176 22720 36228 22729
rect 40316 22720 40368 22772
rect 30104 22627 30156 22636
rect 17040 22516 17092 22568
rect 20536 22559 20588 22568
rect 20536 22525 20545 22559
rect 20545 22525 20579 22559
rect 20579 22525 20588 22559
rect 20536 22516 20588 22525
rect 21180 22516 21232 22568
rect 25228 22516 25280 22568
rect 25596 22516 25648 22568
rect 26056 22516 26108 22568
rect 22008 22448 22060 22500
rect 22192 22448 22244 22500
rect 17224 22380 17276 22432
rect 17316 22380 17368 22432
rect 19892 22423 19944 22432
rect 19892 22389 19901 22423
rect 19901 22389 19935 22423
rect 19935 22389 19944 22423
rect 19892 22380 19944 22389
rect 20444 22380 20496 22432
rect 27896 22448 27948 22500
rect 24952 22380 25004 22432
rect 25596 22380 25648 22432
rect 27436 22380 27488 22432
rect 28908 22380 28960 22432
rect 29552 22448 29604 22500
rect 30104 22593 30113 22627
rect 30113 22593 30147 22627
rect 30147 22593 30156 22627
rect 30104 22584 30156 22593
rect 30288 22584 30340 22636
rect 30840 22627 30892 22636
rect 30840 22593 30849 22627
rect 30849 22593 30883 22627
rect 30883 22593 30892 22627
rect 30840 22584 30892 22593
rect 31116 22584 31168 22636
rect 32128 22584 32180 22636
rect 33784 22627 33836 22636
rect 33784 22593 33793 22627
rect 33793 22593 33827 22627
rect 33827 22593 33836 22627
rect 33784 22584 33836 22593
rect 34244 22584 34296 22636
rect 34520 22584 34572 22636
rect 35348 22627 35400 22636
rect 35348 22593 35357 22627
rect 35357 22593 35391 22627
rect 35391 22593 35400 22627
rect 35348 22584 35400 22593
rect 30380 22516 30432 22568
rect 31484 22516 31536 22568
rect 35532 22584 35584 22636
rect 31116 22491 31168 22500
rect 31116 22457 31125 22491
rect 31125 22457 31159 22491
rect 31159 22457 31168 22491
rect 31116 22448 31168 22457
rect 30104 22380 30156 22432
rect 35992 22516 36044 22568
rect 37832 22627 37884 22636
rect 37832 22593 37841 22627
rect 37841 22593 37875 22627
rect 37875 22593 37884 22627
rect 37832 22584 37884 22593
rect 38660 22584 38712 22636
rect 38844 22584 38896 22636
rect 39028 22627 39080 22636
rect 39028 22593 39038 22627
rect 39038 22593 39072 22627
rect 39072 22593 39080 22627
rect 39028 22584 39080 22593
rect 39212 22627 39264 22636
rect 39212 22593 39221 22627
rect 39221 22593 39255 22627
rect 39255 22593 39264 22627
rect 39212 22584 39264 22593
rect 39580 22584 39632 22636
rect 36544 22516 36596 22568
rect 37280 22516 37332 22568
rect 37556 22516 37608 22568
rect 34152 22491 34204 22500
rect 34152 22457 34161 22491
rect 34161 22457 34195 22491
rect 34195 22457 34204 22491
rect 34152 22448 34204 22457
rect 34244 22448 34296 22500
rect 36544 22380 36596 22432
rect 37372 22448 37424 22500
rect 39304 22516 39356 22568
rect 39212 22380 39264 22432
rect 39580 22423 39632 22432
rect 39580 22389 39589 22423
rect 39589 22389 39623 22423
rect 39623 22389 39632 22423
rect 39580 22380 39632 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 13636 22176 13688 22228
rect 20536 22176 20588 22228
rect 23848 22176 23900 22228
rect 25228 22176 25280 22228
rect 25780 22176 25832 22228
rect 20444 22108 20496 22160
rect 22100 22108 22152 22160
rect 31116 22176 31168 22228
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 10692 21972 10744 22024
rect 11980 21972 12032 22024
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 17040 22040 17092 22092
rect 18696 22040 18748 22092
rect 20352 22040 20404 22092
rect 28632 22108 28684 22160
rect 34796 22176 34848 22228
rect 35992 22176 36044 22228
rect 36636 22176 36688 22228
rect 40132 22176 40184 22228
rect 43168 22219 43220 22228
rect 43168 22185 43177 22219
rect 43177 22185 43211 22219
rect 43211 22185 43220 22219
rect 43168 22176 43220 22185
rect 15200 21972 15252 22024
rect 17316 21972 17368 22024
rect 19432 21972 19484 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 19984 22015 20036 22024
rect 19984 21981 19993 22015
rect 19993 21981 20027 22015
rect 20027 21981 20036 22015
rect 19984 21972 20036 21981
rect 20260 21972 20312 22024
rect 20628 21972 20680 22024
rect 21456 21972 21508 22024
rect 22192 22015 22244 22024
rect 22192 21981 22201 22015
rect 22201 21981 22235 22015
rect 22235 21981 22244 22015
rect 22192 21972 22244 21981
rect 15016 21904 15068 21956
rect 12164 21879 12216 21888
rect 12164 21845 12173 21879
rect 12173 21845 12207 21879
rect 12207 21845 12216 21879
rect 12164 21836 12216 21845
rect 12256 21836 12308 21888
rect 14648 21836 14700 21888
rect 15108 21879 15160 21888
rect 15108 21845 15117 21879
rect 15117 21845 15151 21879
rect 15151 21845 15160 21879
rect 15108 21836 15160 21845
rect 18696 21904 18748 21956
rect 21272 21904 21324 21956
rect 21364 21904 21416 21956
rect 22560 21972 22612 22024
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 25136 21972 25188 22024
rect 27068 21972 27120 22024
rect 23020 21904 23072 21956
rect 19984 21836 20036 21888
rect 20168 21836 20220 21888
rect 23296 21836 23348 21888
rect 24676 21879 24728 21888
rect 24676 21845 24685 21879
rect 24685 21845 24719 21879
rect 24719 21845 24728 21879
rect 24676 21836 24728 21845
rect 25596 21904 25648 21956
rect 27620 21972 27672 22024
rect 27988 22015 28040 22024
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 27988 21972 28040 21981
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 28264 21972 28316 22024
rect 30012 22083 30064 22092
rect 30012 22049 30021 22083
rect 30021 22049 30055 22083
rect 30055 22049 30064 22083
rect 30012 22040 30064 22049
rect 31208 22040 31260 22092
rect 33048 22040 33100 22092
rect 30288 22015 30340 22024
rect 30288 21981 30297 22015
rect 30297 21981 30331 22015
rect 30331 21981 30340 22015
rect 30288 21972 30340 21981
rect 25872 21836 25924 21888
rect 26976 21879 27028 21888
rect 26976 21845 26985 21879
rect 26985 21845 27019 21879
rect 27019 21845 27028 21879
rect 26976 21836 27028 21845
rect 30932 21904 30984 21956
rect 32312 21904 32364 21956
rect 33600 21972 33652 22024
rect 37924 22108 37976 22160
rect 39120 22108 39172 22160
rect 34980 22040 35032 22092
rect 40408 22040 40460 22092
rect 33416 21904 33468 21956
rect 34060 21904 34112 21956
rect 34244 21904 34296 21956
rect 34336 21904 34388 21956
rect 27712 21836 27764 21888
rect 29644 21836 29696 21888
rect 31116 21836 31168 21888
rect 33784 21836 33836 21888
rect 34428 21836 34480 21888
rect 40040 21972 40092 22024
rect 41880 21972 41932 22024
rect 42064 22015 42116 22024
rect 42064 21981 42098 22015
rect 42098 21981 42116 22015
rect 42064 21972 42116 21981
rect 35072 21879 35124 21888
rect 35072 21845 35081 21879
rect 35081 21845 35115 21879
rect 35115 21845 35124 21879
rect 35072 21836 35124 21845
rect 35348 21836 35400 21888
rect 39304 21836 39356 21888
rect 40132 21947 40184 21956
rect 40132 21913 40141 21947
rect 40141 21913 40175 21947
rect 40175 21913 40184 21947
rect 40132 21904 40184 21913
rect 39580 21836 39632 21888
rect 39764 21836 39816 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 16212 21632 16264 21684
rect 23204 21632 23256 21684
rect 24676 21632 24728 21684
rect 25596 21675 25648 21684
rect 25596 21641 25605 21675
rect 25605 21641 25639 21675
rect 25639 21641 25648 21675
rect 25596 21632 25648 21641
rect 27528 21632 27580 21684
rect 27988 21632 28040 21684
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 14648 21496 14700 21548
rect 15016 21539 15068 21548
rect 15016 21505 15025 21539
rect 15025 21505 15059 21539
rect 15059 21505 15068 21539
rect 15016 21496 15068 21505
rect 15108 21496 15160 21548
rect 20352 21607 20404 21616
rect 20352 21573 20361 21607
rect 20361 21573 20395 21607
rect 20395 21573 20404 21607
rect 20352 21564 20404 21573
rect 16120 21496 16172 21548
rect 21364 21539 21416 21548
rect 21364 21505 21373 21539
rect 21373 21505 21407 21539
rect 21407 21505 21416 21539
rect 21364 21496 21416 21505
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 13544 21428 13596 21480
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 21180 21471 21232 21480
rect 21180 21437 21189 21471
rect 21189 21437 21223 21471
rect 21223 21437 21232 21471
rect 21180 21428 21232 21437
rect 23020 21539 23072 21548
rect 23020 21505 23029 21539
rect 23029 21505 23063 21539
rect 23063 21505 23072 21539
rect 28080 21564 28132 21616
rect 23020 21496 23072 21505
rect 24860 21496 24912 21548
rect 25688 21496 25740 21548
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 27528 21496 27580 21548
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 27896 21496 27948 21548
rect 31116 21632 31168 21684
rect 31208 21607 31260 21616
rect 31208 21573 31217 21607
rect 31217 21573 31251 21607
rect 31251 21573 31260 21607
rect 31208 21564 31260 21573
rect 31300 21564 31352 21616
rect 13268 21360 13320 21412
rect 13728 21360 13780 21412
rect 15752 21335 15804 21344
rect 15752 21301 15761 21335
rect 15761 21301 15795 21335
rect 15795 21301 15804 21335
rect 15752 21292 15804 21301
rect 20168 21360 20220 21412
rect 23204 21428 23256 21480
rect 24952 21471 25004 21480
rect 24952 21437 24961 21471
rect 24961 21437 24995 21471
rect 24995 21437 25004 21471
rect 24952 21428 25004 21437
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 25596 21471 25648 21480
rect 25596 21437 25605 21471
rect 25605 21437 25639 21471
rect 25639 21437 25648 21471
rect 25596 21428 25648 21437
rect 27068 21428 27120 21480
rect 28540 21428 28592 21480
rect 30472 21428 30524 21480
rect 31116 21471 31168 21480
rect 31116 21437 31125 21471
rect 31125 21437 31159 21471
rect 31159 21437 31168 21471
rect 31116 21428 31168 21437
rect 33416 21496 33468 21548
rect 29368 21360 29420 21412
rect 32312 21471 32364 21480
rect 32312 21437 32321 21471
rect 32321 21437 32355 21471
rect 32355 21437 32364 21471
rect 32312 21428 32364 21437
rect 33600 21428 33652 21480
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 22744 21292 22796 21344
rect 24860 21292 24912 21344
rect 25596 21292 25648 21344
rect 33140 21292 33192 21344
rect 33968 21607 34020 21616
rect 33968 21573 33977 21607
rect 33977 21573 34011 21607
rect 34011 21573 34020 21607
rect 33968 21564 34020 21573
rect 34704 21632 34756 21684
rect 35624 21632 35676 21684
rect 37464 21632 37516 21684
rect 35072 21564 35124 21616
rect 37280 21564 37332 21616
rect 34152 21539 34204 21548
rect 34152 21505 34161 21539
rect 34161 21505 34195 21539
rect 34195 21505 34204 21539
rect 34152 21496 34204 21505
rect 34244 21360 34296 21412
rect 34336 21403 34388 21412
rect 34336 21369 34345 21403
rect 34345 21369 34379 21403
rect 34379 21369 34388 21403
rect 34336 21360 34388 21369
rect 34520 21428 34572 21480
rect 34704 21428 34756 21480
rect 34796 21428 34848 21480
rect 35532 21428 35584 21480
rect 36084 21428 36136 21480
rect 36268 21496 36320 21548
rect 37556 21496 37608 21548
rect 39212 21632 39264 21684
rect 39304 21632 39356 21684
rect 39948 21632 40000 21684
rect 40040 21632 40092 21684
rect 43168 21607 43220 21616
rect 43168 21573 43177 21607
rect 43177 21573 43211 21607
rect 43211 21573 43220 21607
rect 43168 21564 43220 21573
rect 38660 21539 38712 21548
rect 38660 21505 38669 21539
rect 38669 21505 38703 21539
rect 38703 21505 38712 21539
rect 38660 21496 38712 21505
rect 38752 21539 38804 21548
rect 38752 21505 38762 21539
rect 38762 21505 38796 21539
rect 38796 21505 38804 21539
rect 38752 21496 38804 21505
rect 37188 21428 37240 21480
rect 37740 21428 37792 21480
rect 39396 21496 39448 21548
rect 40592 21496 40644 21548
rect 41972 21496 42024 21548
rect 42708 21496 42760 21548
rect 37832 21360 37884 21412
rect 40316 21360 40368 21412
rect 34520 21292 34572 21344
rect 36728 21292 36780 21344
rect 38384 21292 38436 21344
rect 39396 21292 39448 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 16764 21088 16816 21140
rect 17132 21088 17184 21140
rect 18420 21088 18472 21140
rect 24768 21088 24820 21140
rect 24952 21131 25004 21140
rect 24952 21097 24961 21131
rect 24961 21097 24995 21131
rect 24995 21097 25004 21131
rect 24952 21088 25004 21097
rect 14648 21020 14700 21072
rect 16672 21020 16724 21072
rect 19340 21020 19392 21072
rect 20904 21020 20956 21072
rect 25136 21131 25188 21140
rect 25136 21097 25145 21131
rect 25145 21097 25179 21131
rect 25179 21097 25188 21131
rect 25136 21088 25188 21097
rect 25688 21131 25740 21140
rect 25688 21097 25697 21131
rect 25697 21097 25731 21131
rect 25731 21097 25740 21131
rect 25688 21088 25740 21097
rect 29000 21088 29052 21140
rect 29736 21131 29788 21140
rect 29736 21097 29745 21131
rect 29745 21097 29779 21131
rect 29779 21097 29788 21131
rect 29736 21088 29788 21097
rect 30380 21088 30432 21140
rect 32220 21088 32272 21140
rect 27436 21020 27488 21072
rect 27804 21020 27856 21072
rect 29368 21020 29420 21072
rect 29460 21020 29512 21072
rect 30288 21020 30340 21072
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 13268 20884 13320 20936
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 15108 20884 15160 20936
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 16120 20884 16172 20936
rect 16212 20927 16264 20936
rect 16212 20893 16221 20927
rect 16221 20893 16255 20927
rect 16255 20893 16264 20927
rect 16212 20884 16264 20893
rect 17132 20995 17184 21004
rect 17132 20961 17141 20995
rect 17141 20961 17175 20995
rect 17175 20961 17184 20995
rect 17132 20952 17184 20961
rect 21456 20952 21508 21004
rect 25872 20952 25924 21004
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 22192 20884 22244 20936
rect 23388 20884 23440 20936
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 20168 20816 20220 20868
rect 24860 20884 24912 20936
rect 25228 20884 25280 20936
rect 25320 20884 25372 20936
rect 26976 20884 27028 20936
rect 25872 20816 25924 20868
rect 27804 20859 27856 20868
rect 20628 20748 20680 20800
rect 21364 20748 21416 20800
rect 22836 20748 22888 20800
rect 23296 20748 23348 20800
rect 24768 20748 24820 20800
rect 27804 20825 27813 20859
rect 27813 20825 27847 20859
rect 27847 20825 27856 20859
rect 27804 20816 27856 20825
rect 28080 20859 28132 20868
rect 28080 20825 28089 20859
rect 28089 20825 28123 20859
rect 28123 20825 28132 20859
rect 28080 20816 28132 20825
rect 29644 20884 29696 20936
rect 30012 20884 30064 20936
rect 31576 21020 31628 21072
rect 31852 20952 31904 21004
rect 32404 20995 32456 21004
rect 32404 20961 32413 20995
rect 32413 20961 32447 20995
rect 32447 20961 32456 20995
rect 32404 20952 32456 20961
rect 33600 20952 33652 21004
rect 31576 20927 31628 20936
rect 31576 20893 31585 20927
rect 31585 20893 31619 20927
rect 31619 20893 31628 20927
rect 31576 20884 31628 20893
rect 31760 20884 31812 20936
rect 33692 20884 33744 20936
rect 33876 20816 33928 20868
rect 34428 20952 34480 21004
rect 34152 20927 34204 20936
rect 34152 20893 34161 20927
rect 34161 20893 34195 20927
rect 34195 20893 34204 20927
rect 34152 20884 34204 20893
rect 36728 21020 36780 21072
rect 36544 20952 36596 21004
rect 37832 20995 37884 21004
rect 37832 20961 37841 20995
rect 37841 20961 37875 20995
rect 37875 20961 37884 20995
rect 37832 20952 37884 20961
rect 27528 20748 27580 20800
rect 29920 20748 29972 20800
rect 30288 20748 30340 20800
rect 34704 20816 34756 20868
rect 35440 20927 35492 20936
rect 35440 20893 35449 20927
rect 35449 20893 35483 20927
rect 35483 20893 35492 20927
rect 35440 20884 35492 20893
rect 34796 20748 34848 20800
rect 34888 20791 34940 20800
rect 34888 20757 34897 20791
rect 34897 20757 34931 20791
rect 34931 20757 34940 20791
rect 34888 20748 34940 20757
rect 36728 20859 36780 20868
rect 36728 20825 36737 20859
rect 36737 20825 36771 20859
rect 36771 20825 36780 20859
rect 36728 20816 36780 20825
rect 37188 20884 37240 20936
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 40592 21131 40644 21140
rect 40592 21097 40601 21131
rect 40601 21097 40635 21131
rect 40635 21097 40644 21131
rect 40592 21088 40644 21097
rect 40408 21020 40460 21072
rect 39304 20952 39356 21004
rect 39396 20995 39448 21004
rect 39396 20961 39405 20995
rect 39405 20961 39439 20995
rect 39439 20961 39448 20995
rect 39396 20952 39448 20961
rect 40132 20995 40184 21004
rect 40132 20961 40141 20995
rect 40141 20961 40175 20995
rect 40175 20961 40184 20995
rect 40132 20952 40184 20961
rect 43260 20952 43312 21004
rect 37556 20816 37608 20868
rect 39764 20884 39816 20936
rect 40132 20816 40184 20868
rect 42708 20816 42760 20868
rect 37188 20748 37240 20800
rect 37648 20748 37700 20800
rect 39304 20791 39356 20800
rect 39304 20757 39313 20791
rect 39313 20757 39347 20791
rect 39347 20757 39356 20791
rect 39304 20748 39356 20757
rect 42524 20791 42576 20800
rect 42524 20757 42533 20791
rect 42533 20757 42567 20791
rect 42567 20757 42576 20791
rect 42524 20748 42576 20757
rect 42800 20748 42852 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 13268 20544 13320 20596
rect 14740 20544 14792 20596
rect 17132 20544 17184 20596
rect 27896 20544 27948 20596
rect 28724 20544 28776 20596
rect 29920 20544 29972 20596
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 15108 20408 15160 20460
rect 15200 20408 15252 20460
rect 20168 20476 20220 20528
rect 14556 20340 14608 20392
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 14924 20340 14976 20349
rect 18880 20408 18932 20460
rect 18144 20340 18196 20392
rect 20076 20408 20128 20460
rect 20352 20408 20404 20460
rect 22744 20476 22796 20528
rect 24216 20476 24268 20528
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 22100 20408 22152 20460
rect 22652 20408 22704 20460
rect 19340 20340 19392 20392
rect 23940 20408 23992 20460
rect 24860 20451 24912 20460
rect 24860 20417 24869 20451
rect 24869 20417 24903 20451
rect 24903 20417 24912 20451
rect 24860 20408 24912 20417
rect 25688 20408 25740 20460
rect 26056 20408 26108 20460
rect 27068 20408 27120 20460
rect 25320 20340 25372 20392
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 28540 20451 28592 20460
rect 28540 20417 28544 20451
rect 28544 20417 28578 20451
rect 28578 20417 28592 20451
rect 28540 20408 28592 20417
rect 27896 20340 27948 20392
rect 15292 20272 15344 20324
rect 18512 20315 18564 20324
rect 18512 20281 18521 20315
rect 18521 20281 18555 20315
rect 18555 20281 18564 20315
rect 18512 20272 18564 20281
rect 23388 20272 23440 20324
rect 24032 20272 24084 20324
rect 28724 20451 28776 20460
rect 28724 20417 28733 20451
rect 28733 20417 28767 20451
rect 28767 20417 28776 20451
rect 28724 20408 28776 20417
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 30104 20519 30156 20528
rect 30104 20485 30113 20519
rect 30113 20485 30147 20519
rect 30147 20485 30156 20519
rect 30104 20476 30156 20485
rect 30380 20544 30432 20596
rect 34060 20544 34112 20596
rect 30656 20408 30708 20460
rect 33692 20340 33744 20392
rect 34244 20451 34296 20460
rect 34244 20417 34253 20451
rect 34253 20417 34287 20451
rect 34287 20417 34296 20451
rect 34244 20408 34296 20417
rect 34888 20476 34940 20528
rect 35348 20519 35400 20528
rect 35348 20485 35357 20519
rect 35357 20485 35391 20519
rect 35391 20485 35400 20519
rect 35348 20476 35400 20485
rect 34520 20451 34572 20460
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 34796 20408 34848 20460
rect 35256 20451 35308 20460
rect 35256 20417 35265 20451
rect 35265 20417 35299 20451
rect 35299 20417 35308 20451
rect 35256 20408 35308 20417
rect 39028 20544 39080 20596
rect 42708 20544 42760 20596
rect 38844 20408 38896 20460
rect 39120 20451 39172 20460
rect 39120 20417 39130 20451
rect 39130 20417 39164 20451
rect 39164 20417 39172 20451
rect 39120 20408 39172 20417
rect 37372 20340 37424 20392
rect 37740 20340 37792 20392
rect 38752 20340 38804 20392
rect 39488 20451 39540 20460
rect 39488 20417 39502 20451
rect 39502 20417 39536 20451
rect 39536 20417 39540 20451
rect 39488 20408 39540 20417
rect 40132 20451 40184 20460
rect 40132 20417 40141 20451
rect 40141 20417 40175 20451
rect 40175 20417 40184 20451
rect 40132 20408 40184 20417
rect 40408 20451 40460 20460
rect 40408 20417 40417 20451
rect 40417 20417 40451 20451
rect 40451 20417 40460 20451
rect 40408 20408 40460 20417
rect 42708 20408 42760 20460
rect 42800 20340 42852 20392
rect 43168 20383 43220 20392
rect 43168 20349 43177 20383
rect 43177 20349 43211 20383
rect 43211 20349 43220 20383
rect 43168 20340 43220 20349
rect 23020 20204 23072 20256
rect 24952 20204 25004 20256
rect 27252 20247 27304 20256
rect 27252 20213 27261 20247
rect 27261 20213 27295 20247
rect 27295 20213 27304 20247
rect 27252 20204 27304 20213
rect 29828 20247 29880 20256
rect 29828 20213 29837 20247
rect 29837 20213 29871 20247
rect 29871 20213 29880 20247
rect 29828 20204 29880 20213
rect 32220 20204 32272 20256
rect 34704 20204 34756 20256
rect 37464 20272 37516 20324
rect 42984 20272 43036 20324
rect 37556 20204 37608 20256
rect 40132 20204 40184 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 14096 20000 14148 20052
rect 15384 20000 15436 20052
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 24860 20000 24912 20052
rect 28356 20000 28408 20052
rect 15476 19864 15528 19916
rect 16028 19864 16080 19916
rect 14832 19796 14884 19848
rect 18328 19932 18380 19984
rect 22652 19932 22704 19984
rect 24676 19932 24728 19984
rect 24768 19932 24820 19984
rect 20352 19864 20404 19916
rect 20904 19864 20956 19916
rect 23756 19907 23808 19916
rect 23756 19873 23765 19907
rect 23765 19873 23799 19907
rect 23799 19873 23808 19907
rect 23756 19864 23808 19873
rect 18420 19796 18472 19848
rect 20076 19796 20128 19848
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 25044 19864 25096 19916
rect 27804 19864 27856 19916
rect 14556 19728 14608 19780
rect 20628 19728 20680 19780
rect 23940 19839 23992 19848
rect 23940 19805 23949 19839
rect 23949 19805 23983 19839
rect 23983 19805 23992 19839
rect 23940 19796 23992 19805
rect 24216 19796 24268 19848
rect 24860 19796 24912 19848
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 25504 19796 25556 19848
rect 23388 19728 23440 19780
rect 19432 19660 19484 19712
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 22560 19660 22612 19712
rect 23112 19660 23164 19712
rect 25228 19771 25280 19780
rect 25228 19737 25237 19771
rect 25237 19737 25271 19771
rect 25271 19737 25280 19771
rect 25228 19728 25280 19737
rect 27252 19796 27304 19848
rect 28080 19839 28132 19848
rect 28080 19805 28103 19839
rect 28103 19805 28132 19839
rect 28080 19796 28132 19805
rect 28172 19839 28224 19848
rect 28172 19805 28181 19839
rect 28181 19805 28215 19839
rect 28215 19805 28224 19839
rect 28172 19796 28224 19805
rect 28448 19771 28500 19780
rect 28448 19737 28457 19771
rect 28457 19737 28491 19771
rect 28491 19737 28500 19771
rect 28448 19728 28500 19737
rect 29460 20000 29512 20052
rect 29644 20000 29696 20052
rect 30656 20043 30708 20052
rect 30656 20009 30665 20043
rect 30665 20009 30699 20043
rect 30699 20009 30708 20043
rect 30656 20000 30708 20009
rect 33692 20000 33744 20052
rect 37372 20000 37424 20052
rect 40040 20000 40092 20052
rect 41420 20000 41472 20052
rect 42800 20000 42852 20052
rect 28908 19932 28960 19984
rect 31852 19932 31904 19984
rect 37280 19932 37332 19984
rect 37924 19932 37976 19984
rect 39028 19932 39080 19984
rect 29736 19907 29788 19916
rect 29092 19796 29144 19848
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 29920 19864 29972 19916
rect 29460 19796 29512 19848
rect 30012 19839 30064 19848
rect 30012 19805 30021 19839
rect 30021 19805 30055 19839
rect 30055 19805 30064 19839
rect 30012 19796 30064 19805
rect 30104 19796 30156 19848
rect 31116 19864 31168 19916
rect 31760 19839 31812 19848
rect 31760 19805 31769 19839
rect 31769 19805 31803 19839
rect 31803 19805 31812 19839
rect 31760 19796 31812 19805
rect 31852 19839 31904 19848
rect 31852 19805 31861 19839
rect 31861 19805 31895 19839
rect 31895 19805 31904 19839
rect 31852 19796 31904 19805
rect 33876 19839 33928 19848
rect 33876 19805 33880 19839
rect 33880 19805 33914 19839
rect 33914 19805 33928 19839
rect 33876 19796 33928 19805
rect 34060 19839 34112 19848
rect 34060 19805 34069 19839
rect 34069 19805 34103 19839
rect 34103 19805 34112 19839
rect 34060 19796 34112 19805
rect 34336 19839 34388 19848
rect 34336 19805 34345 19839
rect 34345 19805 34379 19839
rect 34379 19805 34388 19839
rect 34336 19796 34388 19805
rect 36084 19796 36136 19848
rect 30380 19728 30432 19780
rect 32588 19728 32640 19780
rect 33416 19728 33468 19780
rect 34428 19728 34480 19780
rect 26056 19660 26108 19712
rect 27896 19703 27948 19712
rect 27896 19669 27905 19703
rect 27905 19669 27939 19703
rect 27939 19669 27948 19703
rect 27896 19660 27948 19669
rect 28724 19660 28776 19712
rect 33692 19703 33744 19712
rect 33692 19669 33701 19703
rect 33701 19669 33735 19703
rect 33735 19669 33744 19703
rect 33692 19660 33744 19669
rect 37188 19839 37240 19848
rect 37188 19805 37198 19839
rect 37198 19805 37232 19839
rect 37232 19805 37240 19839
rect 37188 19796 37240 19805
rect 37280 19796 37332 19848
rect 37464 19839 37516 19848
rect 37464 19805 37473 19839
rect 37473 19805 37507 19839
rect 37507 19805 37516 19839
rect 37464 19796 37516 19805
rect 37556 19839 37608 19848
rect 37556 19805 37570 19839
rect 37570 19805 37604 19839
rect 37604 19805 37608 19839
rect 37556 19796 37608 19805
rect 38752 19796 38804 19848
rect 38844 19839 38896 19848
rect 38844 19805 38853 19839
rect 38853 19805 38887 19839
rect 38887 19805 38896 19839
rect 38844 19796 38896 19805
rect 38936 19839 38988 19848
rect 38936 19805 38946 19839
rect 38946 19805 38980 19839
rect 38980 19805 38988 19839
rect 38936 19796 38988 19805
rect 39028 19796 39080 19848
rect 40132 19907 40184 19916
rect 40132 19873 40141 19907
rect 40141 19873 40175 19907
rect 40175 19873 40184 19907
rect 40132 19864 40184 19873
rect 37832 19660 37884 19712
rect 38752 19660 38804 19712
rect 39488 19796 39540 19848
rect 39672 19796 39724 19848
rect 40316 19839 40368 19848
rect 40316 19805 40325 19839
rect 40325 19805 40359 19839
rect 40359 19805 40368 19839
rect 40316 19796 40368 19805
rect 41512 19796 41564 19848
rect 42524 19796 42576 19848
rect 41604 19728 41656 19780
rect 41696 19660 41748 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 15108 19456 15160 19508
rect 19432 19456 19484 19508
rect 20260 19456 20312 19508
rect 22928 19499 22980 19508
rect 22928 19465 22937 19499
rect 22937 19465 22971 19499
rect 22971 19465 22980 19499
rect 22928 19456 22980 19465
rect 23020 19456 23072 19508
rect 23848 19456 23900 19508
rect 23940 19499 23992 19508
rect 23940 19465 23949 19499
rect 23949 19465 23983 19499
rect 23983 19465 23992 19499
rect 23940 19456 23992 19465
rect 11980 19320 12032 19372
rect 15752 19388 15804 19440
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 17224 19388 17276 19440
rect 25504 19456 25556 19508
rect 28724 19499 28776 19508
rect 28724 19465 28733 19499
rect 28733 19465 28767 19499
rect 28767 19465 28776 19499
rect 28724 19456 28776 19465
rect 28908 19456 28960 19508
rect 29920 19456 29972 19508
rect 31760 19499 31812 19508
rect 31760 19465 31769 19499
rect 31769 19465 31803 19499
rect 31803 19465 31812 19499
rect 31760 19456 31812 19465
rect 16948 19320 17000 19372
rect 14280 19252 14332 19304
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 13728 19227 13780 19236
rect 13728 19193 13737 19227
rect 13737 19193 13771 19227
rect 13771 19193 13780 19227
rect 13728 19184 13780 19193
rect 14556 19116 14608 19168
rect 15292 19116 15344 19168
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18604 19320 18656 19372
rect 19248 19252 19300 19304
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 24768 19363 24820 19372
rect 24768 19329 24777 19363
rect 24777 19329 24811 19363
rect 24811 19329 24820 19363
rect 24768 19320 24820 19329
rect 25688 19388 25740 19440
rect 29092 19388 29144 19440
rect 25044 19320 25096 19372
rect 25320 19320 25372 19372
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 26056 19320 26108 19329
rect 27804 19320 27856 19372
rect 28356 19320 28408 19372
rect 28448 19320 28500 19372
rect 28908 19320 28960 19372
rect 29644 19320 29696 19372
rect 32128 19388 32180 19440
rect 21272 19252 21324 19304
rect 29000 19252 29052 19304
rect 29092 19295 29144 19304
rect 29092 19261 29101 19295
rect 29101 19261 29135 19295
rect 29135 19261 29144 19295
rect 29092 19252 29144 19261
rect 30104 19252 30156 19304
rect 18420 19116 18472 19168
rect 19708 19116 19760 19168
rect 20904 19116 20956 19168
rect 24860 19184 24912 19236
rect 25872 19184 25924 19236
rect 34428 19456 34480 19508
rect 38844 19456 38896 19508
rect 39672 19456 39724 19508
rect 39764 19499 39816 19508
rect 39764 19465 39773 19499
rect 39773 19465 39807 19499
rect 39807 19465 39816 19499
rect 39764 19456 39816 19465
rect 41604 19499 41656 19508
rect 41604 19465 41613 19499
rect 41613 19465 41647 19499
rect 41647 19465 41656 19499
rect 41604 19456 41656 19465
rect 41696 19499 41748 19508
rect 41696 19465 41705 19499
rect 41705 19465 41739 19499
rect 41739 19465 41748 19499
rect 41696 19456 41748 19465
rect 42892 19456 42944 19508
rect 42984 19499 43036 19508
rect 42984 19465 42993 19499
rect 42993 19465 43027 19499
rect 43027 19465 43036 19499
rect 42984 19456 43036 19465
rect 35716 19388 35768 19440
rect 39304 19388 39356 19440
rect 42708 19388 42760 19440
rect 34244 19320 34296 19372
rect 37372 19320 37424 19372
rect 37648 19320 37700 19372
rect 37832 19363 37884 19372
rect 37832 19329 37841 19363
rect 37841 19329 37875 19363
rect 37875 19329 37884 19363
rect 37832 19320 37884 19329
rect 39580 19363 39632 19372
rect 39580 19329 39589 19363
rect 39589 19329 39623 19363
rect 39623 19329 39632 19363
rect 39580 19320 39632 19329
rect 34704 19252 34756 19304
rect 43260 19252 43312 19304
rect 42708 19184 42760 19236
rect 40132 19116 40184 19168
rect 41236 19159 41288 19168
rect 41236 19125 41245 19159
rect 41245 19125 41279 19159
rect 41279 19125 41288 19159
rect 41236 19116 41288 19125
rect 42616 19159 42668 19168
rect 42616 19125 42625 19159
rect 42625 19125 42659 19159
rect 42659 19125 42668 19159
rect 42616 19116 42668 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 15844 18912 15896 18964
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 15108 18751 15160 18760
rect 15108 18717 15117 18751
rect 15117 18717 15151 18751
rect 15151 18717 15160 18751
rect 15108 18708 15160 18717
rect 15752 18708 15804 18760
rect 16948 18708 17000 18760
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 18144 18708 18196 18760
rect 18420 18708 18472 18760
rect 19340 18708 19392 18760
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 19984 18708 20036 18760
rect 20628 18776 20680 18828
rect 21272 18776 21324 18828
rect 23388 18844 23440 18896
rect 25228 18955 25280 18964
rect 25228 18921 25237 18955
rect 25237 18921 25271 18955
rect 25271 18921 25280 18955
rect 25228 18912 25280 18921
rect 26056 18912 26108 18964
rect 28172 18912 28224 18964
rect 33784 18912 33836 18964
rect 35440 18912 35492 18964
rect 42984 18912 43036 18964
rect 25412 18844 25464 18896
rect 28724 18844 28776 18896
rect 34704 18844 34756 18896
rect 22652 18708 22704 18760
rect 22836 18708 22888 18760
rect 23756 18708 23808 18760
rect 25688 18751 25740 18760
rect 25688 18717 25697 18751
rect 25697 18717 25731 18751
rect 25731 18717 25740 18751
rect 25688 18708 25740 18717
rect 29000 18776 29052 18828
rect 35348 18819 35400 18828
rect 35348 18785 35357 18819
rect 35357 18785 35391 18819
rect 35391 18785 35400 18819
rect 35348 18776 35400 18785
rect 14924 18640 14976 18692
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 16672 18640 16724 18649
rect 18236 18640 18288 18692
rect 28908 18751 28960 18760
rect 28908 18717 28917 18751
rect 28917 18717 28951 18751
rect 28951 18717 28960 18751
rect 28908 18708 28960 18717
rect 33692 18708 33744 18760
rect 34796 18708 34848 18760
rect 36268 18751 36320 18760
rect 36268 18717 36277 18751
rect 36277 18717 36311 18751
rect 36311 18717 36320 18751
rect 36268 18708 36320 18717
rect 36452 18751 36504 18760
rect 36452 18717 36461 18751
rect 36461 18717 36495 18751
rect 36495 18717 36504 18751
rect 36452 18708 36504 18717
rect 29092 18640 29144 18692
rect 14832 18572 14884 18624
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 18144 18572 18196 18624
rect 18604 18572 18656 18624
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 20996 18615 21048 18624
rect 20996 18581 21005 18615
rect 21005 18581 21039 18615
rect 21039 18581 21048 18615
rect 20996 18572 21048 18581
rect 21364 18615 21416 18624
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 22928 18572 22980 18624
rect 39580 18640 39632 18692
rect 40684 18708 40736 18760
rect 41512 18708 41564 18760
rect 42616 18708 42668 18760
rect 42800 18640 42852 18692
rect 37556 18572 37608 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 15476 18368 15528 18420
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 19984 18368 20036 18420
rect 21272 18368 21324 18420
rect 22928 18411 22980 18420
rect 22928 18377 22937 18411
rect 22937 18377 22971 18411
rect 22971 18377 22980 18411
rect 22928 18368 22980 18377
rect 29000 18368 29052 18420
rect 38844 18411 38896 18420
rect 38844 18377 38853 18411
rect 38853 18377 38887 18411
rect 38887 18377 38896 18411
rect 38844 18368 38896 18377
rect 41604 18368 41656 18420
rect 17960 18300 18012 18352
rect 18236 18300 18288 18352
rect 14924 18232 14976 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 21364 18300 21416 18352
rect 23020 18343 23072 18352
rect 23020 18309 23029 18343
rect 23029 18309 23063 18343
rect 23063 18309 23072 18343
rect 23020 18300 23072 18309
rect 29092 18300 29144 18352
rect 30196 18343 30248 18352
rect 30196 18309 30205 18343
rect 30205 18309 30239 18343
rect 30239 18309 30248 18343
rect 30196 18300 30248 18309
rect 30656 18300 30708 18352
rect 35808 18300 35860 18352
rect 22652 18232 22704 18284
rect 25688 18232 25740 18284
rect 28724 18275 28776 18284
rect 28724 18241 28733 18275
rect 28733 18241 28767 18275
rect 28767 18241 28776 18275
rect 28724 18232 28776 18241
rect 33784 18232 33836 18284
rect 35716 18232 35768 18284
rect 20352 18164 20404 18216
rect 29368 18207 29420 18216
rect 29368 18173 29377 18207
rect 29377 18173 29411 18207
rect 29411 18173 29420 18207
rect 29368 18164 29420 18173
rect 35348 18164 35400 18216
rect 16948 18096 17000 18148
rect 22284 18096 22336 18148
rect 23112 18096 23164 18148
rect 28080 18096 28132 18148
rect 33692 18096 33744 18148
rect 36452 18232 36504 18284
rect 41236 18300 41288 18352
rect 43168 18343 43220 18352
rect 43168 18309 43177 18343
rect 43177 18309 43211 18343
rect 43211 18309 43220 18343
rect 43168 18300 43220 18309
rect 37556 18232 37608 18284
rect 39580 18275 39632 18284
rect 39580 18241 39589 18275
rect 39589 18241 39623 18275
rect 39623 18241 39632 18275
rect 39580 18232 39632 18241
rect 40040 18232 40092 18284
rect 40684 18275 40736 18284
rect 40684 18241 40693 18275
rect 40693 18241 40727 18275
rect 40727 18241 40736 18275
rect 40684 18232 40736 18241
rect 42892 18275 42944 18284
rect 42892 18241 42901 18275
rect 42901 18241 42935 18275
rect 42935 18241 42944 18275
rect 42892 18232 42944 18241
rect 39304 18164 39356 18216
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 23388 18028 23440 18080
rect 36544 18028 36596 18080
rect 40316 18028 40368 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15200 17824 15252 17876
rect 22744 17824 22796 17876
rect 37464 17824 37516 17876
rect 41420 17867 41472 17876
rect 41420 17833 41429 17867
rect 41429 17833 41463 17867
rect 41463 17833 41472 17867
rect 41420 17824 41472 17833
rect 14924 17756 14976 17808
rect 17776 17756 17828 17808
rect 24124 17756 24176 17808
rect 28264 17756 28316 17808
rect 33876 17756 33928 17808
rect 19340 17688 19392 17740
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 17316 17620 17368 17672
rect 16028 17552 16080 17604
rect 17132 17552 17184 17604
rect 19432 17620 19484 17672
rect 22100 17688 22152 17740
rect 22652 17688 22704 17740
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20444 17620 20496 17672
rect 22100 17552 22152 17604
rect 22744 17620 22796 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 26332 17620 26384 17672
rect 29368 17688 29420 17740
rect 31760 17688 31812 17740
rect 35716 17688 35768 17740
rect 27160 17552 27212 17604
rect 27252 17552 27304 17604
rect 28356 17595 28408 17604
rect 28356 17561 28365 17595
rect 28365 17561 28399 17595
rect 28399 17561 28408 17595
rect 28356 17552 28408 17561
rect 30012 17595 30064 17604
rect 30012 17561 30046 17595
rect 30046 17561 30064 17595
rect 30012 17552 30064 17561
rect 31760 17552 31812 17604
rect 33416 17663 33468 17672
rect 33416 17629 33425 17663
rect 33425 17629 33459 17663
rect 33459 17629 33468 17663
rect 33416 17620 33468 17629
rect 15292 17484 15344 17536
rect 18604 17484 18656 17536
rect 22008 17527 22060 17536
rect 22008 17493 22017 17527
rect 22017 17493 22051 17527
rect 22051 17493 22060 17527
rect 22008 17484 22060 17493
rect 22192 17484 22244 17536
rect 27528 17484 27580 17536
rect 31116 17527 31168 17536
rect 31116 17493 31125 17527
rect 31125 17493 31159 17527
rect 31159 17493 31168 17527
rect 31116 17484 31168 17493
rect 31852 17484 31904 17536
rect 35532 17552 35584 17604
rect 35808 17663 35860 17672
rect 35808 17629 35817 17663
rect 35817 17629 35851 17663
rect 35851 17629 35860 17663
rect 35808 17620 35860 17629
rect 36544 17663 36596 17672
rect 36544 17629 36578 17663
rect 36578 17629 36596 17663
rect 36544 17620 36596 17629
rect 40040 17663 40092 17672
rect 40040 17629 40049 17663
rect 40049 17629 40083 17663
rect 40083 17629 40092 17663
rect 40040 17620 40092 17629
rect 40316 17663 40368 17672
rect 40316 17629 40339 17663
rect 40339 17629 40368 17663
rect 40316 17620 40368 17629
rect 42800 17620 42852 17672
rect 35992 17552 36044 17604
rect 43168 17595 43220 17604
rect 43168 17561 43177 17595
rect 43177 17561 43211 17595
rect 43211 17561 43220 17595
rect 43168 17552 43220 17561
rect 37556 17484 37608 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 15384 17280 15436 17332
rect 22468 17280 22520 17332
rect 23296 17280 23348 17332
rect 23572 17280 23624 17332
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17592 17076 17644 17128
rect 19432 17144 19484 17196
rect 19984 17212 20036 17264
rect 20996 17212 21048 17264
rect 22008 17255 22060 17264
rect 22008 17221 22017 17255
rect 22017 17221 22051 17255
rect 22051 17221 22060 17255
rect 22008 17212 22060 17221
rect 22192 17255 22244 17264
rect 22192 17221 22201 17255
rect 22201 17221 22235 17255
rect 22235 17221 22244 17255
rect 22192 17212 22244 17221
rect 22284 17212 22336 17264
rect 20444 17144 20496 17196
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 22468 17144 22520 17196
rect 25780 17212 25832 17264
rect 23572 17144 23624 17196
rect 27160 17323 27212 17332
rect 27160 17289 27169 17323
rect 27169 17289 27203 17323
rect 27203 17289 27212 17323
rect 27160 17280 27212 17289
rect 27528 17323 27580 17332
rect 27528 17289 27537 17323
rect 27537 17289 27571 17323
rect 27571 17289 27580 17323
rect 27528 17280 27580 17289
rect 27712 17280 27764 17332
rect 29920 17280 29972 17332
rect 31760 17323 31812 17332
rect 31760 17289 31769 17323
rect 31769 17289 31803 17323
rect 31803 17289 31812 17323
rect 31760 17280 31812 17289
rect 36268 17280 36320 17332
rect 27436 17212 27488 17264
rect 34796 17212 34848 17264
rect 15568 17008 15620 17060
rect 16212 16940 16264 16992
rect 18788 16940 18840 16992
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 23940 17119 23992 17128
rect 23940 17085 23949 17119
rect 23949 17085 23983 17119
rect 23983 17085 23992 17119
rect 23940 17076 23992 17085
rect 31208 17119 31260 17128
rect 31208 17085 31217 17119
rect 31217 17085 31251 17119
rect 31251 17085 31260 17119
rect 31208 17076 31260 17085
rect 31852 17144 31904 17196
rect 32404 17144 32456 17196
rect 33508 17187 33560 17196
rect 33508 17153 33517 17187
rect 33517 17153 33551 17187
rect 33551 17153 33560 17187
rect 33508 17144 33560 17153
rect 33600 17144 33652 17196
rect 37280 17144 37332 17196
rect 38200 17144 38252 17196
rect 31576 17076 31628 17128
rect 35992 17076 36044 17128
rect 22008 17008 22060 17060
rect 35440 17008 35492 17060
rect 22100 16940 22152 16992
rect 22192 16940 22244 16992
rect 24676 16940 24728 16992
rect 29092 16983 29144 16992
rect 29092 16949 29101 16983
rect 29101 16949 29135 16983
rect 29135 16949 29144 16983
rect 29092 16940 29144 16949
rect 33692 16983 33744 16992
rect 33692 16949 33701 16983
rect 33701 16949 33735 16983
rect 33735 16949 33744 16983
rect 33692 16940 33744 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 17316 16736 17368 16788
rect 17592 16779 17644 16788
rect 17592 16745 17601 16779
rect 17601 16745 17635 16779
rect 17635 16745 17644 16779
rect 17592 16736 17644 16745
rect 23572 16779 23624 16788
rect 23572 16745 23581 16779
rect 23581 16745 23615 16779
rect 23615 16745 23624 16779
rect 23572 16736 23624 16745
rect 23940 16736 23992 16788
rect 22100 16711 22152 16720
rect 22100 16677 22109 16711
rect 22109 16677 22143 16711
rect 22143 16677 22152 16711
rect 22100 16668 22152 16677
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 18604 16600 18656 16652
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 20996 16532 21048 16584
rect 20812 16507 20864 16516
rect 20812 16473 20821 16507
rect 20821 16473 20855 16507
rect 20855 16473 20864 16507
rect 20812 16464 20864 16473
rect 20904 16507 20956 16516
rect 20904 16473 20913 16507
rect 20913 16473 20947 16507
rect 20947 16473 20956 16507
rect 20904 16464 20956 16473
rect 22192 16532 22244 16584
rect 22284 16532 22336 16584
rect 22468 16532 22520 16584
rect 26332 16736 26384 16788
rect 26976 16736 27028 16788
rect 28356 16736 28408 16788
rect 28632 16779 28684 16788
rect 28632 16745 28641 16779
rect 28641 16745 28675 16779
rect 28675 16745 28684 16779
rect 28632 16736 28684 16745
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 24676 16532 24728 16584
rect 27620 16600 27672 16652
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 28540 16600 28592 16652
rect 31116 16600 31168 16652
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 38200 16600 38252 16652
rect 38384 16643 38436 16652
rect 38384 16609 38393 16643
rect 38393 16609 38427 16643
rect 38427 16609 38436 16643
rect 38384 16600 38436 16609
rect 41512 16643 41564 16652
rect 41512 16609 41521 16643
rect 41521 16609 41555 16643
rect 41555 16609 41564 16643
rect 41512 16600 41564 16609
rect 22652 16396 22704 16448
rect 27528 16532 27580 16584
rect 30656 16575 30708 16584
rect 30656 16541 30665 16575
rect 30665 16541 30699 16575
rect 30699 16541 30708 16575
rect 30656 16532 30708 16541
rect 31760 16532 31812 16584
rect 32036 16575 32088 16584
rect 32036 16541 32045 16575
rect 32045 16541 32079 16575
rect 32079 16541 32088 16575
rect 32036 16532 32088 16541
rect 32404 16575 32456 16584
rect 32404 16541 32413 16575
rect 32413 16541 32447 16575
rect 32447 16541 32456 16575
rect 32404 16532 32456 16541
rect 34520 16532 34572 16584
rect 35808 16575 35860 16584
rect 35808 16541 35817 16575
rect 35817 16541 35851 16575
rect 35851 16541 35860 16575
rect 35808 16532 35860 16541
rect 35900 16575 35952 16584
rect 35900 16541 35909 16575
rect 35909 16541 35943 16575
rect 35943 16541 35952 16575
rect 35900 16532 35952 16541
rect 36360 16532 36412 16584
rect 29092 16464 29144 16516
rect 30196 16464 30248 16516
rect 31668 16464 31720 16516
rect 38476 16464 38528 16516
rect 40500 16464 40552 16516
rect 27068 16396 27120 16448
rect 28172 16439 28224 16448
rect 28172 16405 28181 16439
rect 28181 16405 28215 16439
rect 28215 16405 28224 16439
rect 28172 16396 28224 16405
rect 37464 16396 37516 16448
rect 37740 16396 37792 16448
rect 40132 16439 40184 16448
rect 40132 16405 40141 16439
rect 40141 16405 40175 16439
rect 40175 16405 40184 16439
rect 40132 16396 40184 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 23572 16192 23624 16244
rect 27436 16192 27488 16244
rect 30012 16192 30064 16244
rect 31116 16192 31168 16244
rect 31760 16235 31812 16244
rect 31760 16201 31769 16235
rect 31769 16201 31803 16235
rect 31803 16201 31812 16235
rect 31760 16192 31812 16201
rect 37556 16235 37608 16244
rect 37556 16201 37565 16235
rect 37565 16201 37599 16235
rect 37599 16201 37608 16235
rect 37556 16192 37608 16201
rect 38200 16192 38252 16244
rect 40500 16235 40552 16244
rect 40500 16201 40509 16235
rect 40509 16201 40543 16235
rect 40543 16201 40552 16235
rect 40500 16192 40552 16201
rect 22192 16167 22244 16176
rect 22192 16133 22201 16167
rect 22201 16133 22235 16167
rect 22235 16133 22244 16167
rect 22192 16124 22244 16133
rect 22376 16167 22428 16176
rect 22376 16133 22401 16167
rect 22401 16133 22428 16167
rect 22376 16124 22428 16133
rect 22652 16124 22704 16176
rect 23388 16167 23440 16176
rect 23388 16133 23397 16167
rect 23397 16133 23431 16167
rect 23431 16133 23440 16167
rect 23388 16124 23440 16133
rect 29460 16124 29512 16176
rect 30196 16124 30248 16176
rect 18420 16056 18472 16108
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 19984 16056 20036 16108
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20812 16056 20864 16108
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 30288 16056 30340 16108
rect 29920 15988 29972 16040
rect 31116 16099 31168 16108
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 31116 16056 31168 16065
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 33324 16099 33376 16108
rect 33324 16065 33358 16099
rect 33358 16065 33376 16099
rect 30104 15920 30156 15972
rect 33324 16056 33376 16065
rect 35716 16124 35768 16176
rect 35256 16099 35308 16108
rect 35256 16065 35290 16099
rect 35290 16065 35308 16099
rect 35256 16056 35308 16065
rect 37464 16099 37516 16108
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 40132 16099 40184 16108
rect 40132 16065 40141 16099
rect 40141 16065 40175 16099
rect 40175 16065 40184 16099
rect 40132 16056 40184 16065
rect 33048 16031 33100 16040
rect 33048 15997 33057 16031
rect 33057 15997 33091 16031
rect 33091 15997 33100 16031
rect 33048 15988 33100 15997
rect 38476 16031 38528 16040
rect 38476 15997 38485 16031
rect 38485 15997 38519 16031
rect 38519 15997 38528 16031
rect 38476 15988 38528 15997
rect 38660 16031 38712 16040
rect 38660 15997 38669 16031
rect 38669 15997 38703 16031
rect 38703 15997 38712 16031
rect 38660 15988 38712 15997
rect 38844 15988 38896 16040
rect 20904 15852 20956 15904
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 22284 15852 22336 15904
rect 22744 15852 22796 15904
rect 27160 15895 27212 15904
rect 27160 15861 27169 15895
rect 27169 15861 27203 15895
rect 27203 15861 27212 15895
rect 27160 15852 27212 15861
rect 34428 15895 34480 15904
rect 34428 15861 34437 15895
rect 34437 15861 34471 15895
rect 34471 15861 34480 15895
rect 34428 15852 34480 15861
rect 36360 15895 36412 15904
rect 36360 15861 36369 15895
rect 36369 15861 36403 15895
rect 36403 15861 36412 15895
rect 36360 15852 36412 15861
rect 43352 15895 43404 15904
rect 43352 15861 43361 15895
rect 43361 15861 43395 15895
rect 43395 15861 43404 15895
rect 43352 15852 43404 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 22376 15648 22428 15700
rect 27528 15648 27580 15700
rect 34520 15648 34572 15700
rect 35348 15648 35400 15700
rect 38476 15648 38528 15700
rect 20904 15580 20956 15632
rect 24124 15580 24176 15632
rect 29000 15512 29052 15564
rect 29920 15512 29972 15564
rect 30472 15512 30524 15564
rect 18512 15444 18564 15496
rect 18604 15444 18656 15496
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 20352 15444 20404 15496
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 22744 15487 22796 15496
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 23388 15444 23440 15496
rect 26332 15444 26384 15496
rect 28724 15444 28776 15496
rect 30104 15487 30156 15496
rect 30104 15453 30113 15487
rect 30113 15453 30147 15487
rect 30147 15453 30156 15487
rect 30104 15444 30156 15453
rect 22100 15419 22152 15428
rect 22100 15385 22109 15419
rect 22109 15385 22143 15419
rect 22143 15385 22152 15419
rect 22100 15376 22152 15385
rect 24308 15376 24360 15428
rect 25320 15376 25372 15428
rect 27160 15376 27212 15428
rect 19432 15308 19484 15360
rect 31392 15376 31444 15428
rect 35348 15512 35400 15564
rect 35716 15512 35768 15564
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 34428 15444 34480 15496
rect 35532 15444 35584 15496
rect 37740 15487 37792 15496
rect 37740 15453 37774 15487
rect 37774 15453 37792 15487
rect 37740 15444 37792 15453
rect 33968 15419 34020 15428
rect 33968 15385 33977 15419
rect 33977 15385 34011 15419
rect 34011 15385 34020 15419
rect 33968 15376 34020 15385
rect 36360 15376 36412 15428
rect 29736 15351 29788 15360
rect 29736 15317 29745 15351
rect 29745 15317 29779 15351
rect 29779 15317 29788 15351
rect 29736 15308 29788 15317
rect 32036 15351 32088 15360
rect 32036 15317 32045 15351
rect 32045 15317 32079 15351
rect 32079 15317 32088 15351
rect 32036 15308 32088 15317
rect 33140 15308 33192 15360
rect 38200 15308 38252 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 18052 15104 18104 15156
rect 22284 15104 22336 15156
rect 30104 15104 30156 15156
rect 31116 15104 31168 15156
rect 33048 15104 33100 15156
rect 35532 15104 35584 15156
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 18420 14900 18472 14952
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 23296 15036 23348 15088
rect 23664 15036 23716 15088
rect 20720 14968 20772 15020
rect 21088 14968 21140 15020
rect 22100 14968 22152 15020
rect 19432 14900 19484 14952
rect 22560 14968 22612 15020
rect 23112 14968 23164 15020
rect 29736 15036 29788 15088
rect 34428 15036 34480 15088
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 20352 14875 20404 14884
rect 20352 14841 20361 14875
rect 20361 14841 20395 14875
rect 20395 14841 20404 14875
rect 20352 14832 20404 14841
rect 18880 14764 18932 14816
rect 20168 14764 20220 14816
rect 29736 14900 29788 14952
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 31668 14968 31720 15020
rect 33140 14968 33192 15020
rect 34520 14968 34572 15020
rect 35808 15011 35860 15020
rect 35808 14977 35817 15011
rect 35817 14977 35851 15011
rect 35851 14977 35860 15011
rect 35808 14968 35860 14977
rect 35900 15011 35952 15020
rect 35900 14977 35909 15011
rect 35909 14977 35943 15011
rect 35943 14977 35952 15011
rect 35900 14968 35952 14977
rect 32312 14943 32364 14952
rect 32312 14909 32321 14943
rect 32321 14909 32355 14943
rect 32355 14909 32364 14943
rect 32312 14900 32364 14909
rect 38016 15011 38068 15020
rect 38016 14977 38025 15011
rect 38025 14977 38059 15011
rect 38059 14977 38068 15011
rect 38016 14968 38068 14977
rect 38292 15011 38344 15020
rect 23388 14832 23440 14884
rect 32036 14832 32088 14884
rect 23940 14807 23992 14816
rect 23940 14773 23949 14807
rect 23949 14773 23983 14807
rect 23983 14773 23992 14807
rect 23940 14764 23992 14773
rect 28816 14764 28868 14816
rect 31208 14764 31260 14816
rect 33140 14764 33192 14816
rect 33324 14875 33376 14884
rect 33324 14841 33333 14875
rect 33333 14841 33367 14875
rect 33367 14841 33376 14875
rect 33324 14832 33376 14841
rect 33416 14832 33468 14884
rect 35900 14832 35952 14884
rect 38292 14977 38301 15011
rect 38301 14977 38335 15011
rect 38335 14977 38344 15011
rect 38292 14968 38344 14977
rect 38660 15011 38712 15020
rect 38660 14977 38669 15011
rect 38669 14977 38703 15011
rect 38703 14977 38712 15011
rect 38660 14968 38712 14977
rect 39120 15036 39172 15088
rect 39488 14968 39540 15020
rect 38476 14943 38528 14952
rect 38476 14909 38485 14943
rect 38485 14909 38519 14943
rect 38519 14909 38528 14943
rect 38476 14900 38528 14909
rect 39764 14943 39816 14952
rect 39764 14909 39773 14943
rect 39773 14909 39807 14943
rect 39807 14909 39816 14943
rect 39764 14900 39816 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 18420 14603 18472 14612
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 27804 14560 27856 14612
rect 20352 14492 20404 14544
rect 27068 14492 27120 14544
rect 27344 14492 27396 14544
rect 33324 14560 33376 14612
rect 33784 14560 33836 14612
rect 39488 14603 39540 14612
rect 39488 14569 39497 14603
rect 39497 14569 39531 14603
rect 39531 14569 39540 14603
rect 39488 14560 39540 14569
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 22008 14467 22060 14476
rect 22008 14433 22017 14467
rect 22017 14433 22051 14467
rect 22051 14433 22060 14467
rect 22008 14424 22060 14433
rect 25596 14424 25648 14476
rect 19432 14356 19484 14408
rect 20720 14356 20772 14408
rect 21272 14288 21324 14340
rect 23848 14356 23900 14408
rect 26148 14356 26200 14408
rect 27068 14399 27120 14408
rect 27068 14365 27077 14399
rect 27077 14365 27111 14399
rect 27111 14365 27120 14399
rect 27068 14356 27120 14365
rect 27804 14356 27856 14408
rect 30564 14424 30616 14476
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 25136 14288 25188 14340
rect 23664 14220 23716 14272
rect 26976 14288 27028 14340
rect 29000 14288 29052 14340
rect 25504 14220 25556 14272
rect 26608 14220 26660 14272
rect 27988 14220 28040 14272
rect 29920 14331 29972 14340
rect 29920 14297 29929 14331
rect 29929 14297 29963 14331
rect 29963 14297 29972 14331
rect 29920 14288 29972 14297
rect 30196 14288 30248 14340
rect 30472 14331 30524 14340
rect 30472 14297 30481 14331
rect 30481 14297 30515 14331
rect 30515 14297 30524 14331
rect 30472 14288 30524 14297
rect 29184 14263 29236 14272
rect 29184 14229 29193 14263
rect 29193 14229 29227 14263
rect 29227 14229 29236 14263
rect 29184 14220 29236 14229
rect 31668 14356 31720 14408
rect 33048 14356 33100 14408
rect 33140 14356 33192 14408
rect 35716 14424 35768 14476
rect 38844 14467 38896 14476
rect 38844 14433 38853 14467
rect 38853 14433 38887 14467
rect 38887 14433 38896 14467
rect 38844 14424 38896 14433
rect 31576 14288 31628 14340
rect 31392 14220 31444 14272
rect 32772 14288 32824 14340
rect 35992 14356 36044 14408
rect 39120 14399 39172 14408
rect 39120 14365 39129 14399
rect 39129 14365 39163 14399
rect 39163 14365 39172 14399
rect 39120 14356 39172 14365
rect 39764 14356 39816 14408
rect 43352 14399 43404 14408
rect 43352 14365 43361 14399
rect 43361 14365 43395 14399
rect 43395 14365 43404 14399
rect 43352 14356 43404 14365
rect 34428 14288 34480 14340
rect 35440 14220 35492 14272
rect 35900 14263 35952 14272
rect 35900 14229 35909 14263
rect 35909 14229 35943 14263
rect 35943 14229 35952 14263
rect 35900 14220 35952 14229
rect 39948 14288 40000 14340
rect 40408 14288 40460 14340
rect 41420 14263 41472 14272
rect 41420 14229 41429 14263
rect 41429 14229 41463 14263
rect 41463 14229 41472 14263
rect 41420 14220 41472 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 20168 14016 20220 14068
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 27068 14016 27120 14068
rect 27528 14059 27580 14068
rect 27528 14025 27537 14059
rect 27537 14025 27571 14059
rect 27571 14025 27580 14059
rect 27528 14016 27580 14025
rect 30564 14016 30616 14068
rect 32772 14059 32824 14068
rect 32772 14025 32781 14059
rect 32781 14025 32815 14059
rect 32815 14025 32824 14059
rect 32772 14016 32824 14025
rect 33232 14059 33284 14068
rect 33232 14025 33241 14059
rect 33241 14025 33275 14059
rect 33275 14025 33284 14059
rect 33232 14016 33284 14025
rect 34428 14016 34480 14068
rect 34520 14059 34572 14068
rect 34520 14025 34529 14059
rect 34529 14025 34563 14059
rect 34563 14025 34572 14059
rect 34520 14016 34572 14025
rect 23388 13948 23440 14000
rect 19984 13880 20036 13932
rect 20720 13880 20772 13932
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 24768 13880 24820 13932
rect 28172 13948 28224 14000
rect 29184 13948 29236 14000
rect 30288 13948 30340 14000
rect 27436 13880 27488 13932
rect 19432 13812 19484 13864
rect 25136 13744 25188 13796
rect 26608 13855 26660 13864
rect 26608 13821 26617 13855
rect 26617 13821 26651 13855
rect 26651 13821 26660 13855
rect 26608 13812 26660 13821
rect 27344 13812 27396 13864
rect 28724 13855 28776 13864
rect 28724 13821 28733 13855
rect 28733 13821 28767 13855
rect 28767 13821 28776 13855
rect 28724 13812 28776 13821
rect 33784 13948 33836 14000
rect 31668 13923 31720 13932
rect 31668 13889 31677 13923
rect 31677 13889 31711 13923
rect 31711 13889 31720 13923
rect 31668 13880 31720 13889
rect 32036 13880 32088 13932
rect 33324 13855 33376 13864
rect 33324 13821 33333 13855
rect 33333 13821 33367 13855
rect 33367 13821 33376 13855
rect 33324 13812 33376 13821
rect 33968 13880 34020 13932
rect 34796 13880 34848 13932
rect 35532 13948 35584 14000
rect 35900 14016 35952 14068
rect 38476 14016 38528 14068
rect 38384 13948 38436 14000
rect 39948 13991 40000 14000
rect 39948 13957 39957 13991
rect 39957 13957 39991 13991
rect 39991 13957 40000 13991
rect 39948 13948 40000 13957
rect 40408 14059 40460 14068
rect 40408 14025 40417 14059
rect 40417 14025 40451 14059
rect 40451 14025 40460 14059
rect 40408 14016 40460 14025
rect 41420 13948 41472 14000
rect 35440 13923 35492 13932
rect 35440 13889 35474 13923
rect 35474 13889 35492 13923
rect 35440 13880 35492 13889
rect 26424 13787 26476 13796
rect 26424 13753 26433 13787
rect 26433 13753 26467 13787
rect 26467 13753 26476 13787
rect 26424 13744 26476 13753
rect 27252 13744 27304 13796
rect 40224 13744 40276 13796
rect 24676 13676 24728 13728
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 28540 13676 28592 13728
rect 29000 13676 29052 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 23480 13472 23532 13524
rect 27528 13515 27580 13524
rect 27528 13481 27537 13515
rect 27537 13481 27571 13515
rect 27571 13481 27580 13515
rect 27528 13472 27580 13481
rect 23664 13404 23716 13456
rect 32312 13404 32364 13456
rect 38660 13404 38712 13456
rect 25320 13379 25372 13388
rect 25320 13345 25329 13379
rect 25329 13345 25363 13379
rect 25363 13345 25372 13379
rect 25320 13336 25372 13345
rect 23940 13268 23992 13320
rect 26148 13311 26200 13320
rect 26148 13277 26157 13311
rect 26157 13277 26191 13311
rect 26191 13277 26200 13311
rect 26148 13268 26200 13277
rect 28540 13268 28592 13320
rect 29736 13268 29788 13320
rect 33968 13336 34020 13388
rect 37280 13336 37332 13388
rect 38844 13404 38896 13456
rect 32956 13268 33008 13320
rect 23204 13243 23256 13252
rect 23204 13209 23213 13243
rect 23213 13209 23247 13243
rect 23247 13209 23256 13243
rect 23204 13200 23256 13209
rect 27160 13200 27212 13252
rect 29920 13200 29972 13252
rect 34704 13268 34756 13320
rect 35808 13311 35860 13320
rect 35808 13277 35817 13311
rect 35817 13277 35851 13311
rect 35851 13277 35860 13311
rect 35808 13268 35860 13277
rect 35900 13311 35952 13320
rect 35900 13277 35909 13311
rect 35909 13277 35943 13311
rect 35943 13277 35952 13311
rect 35900 13268 35952 13277
rect 36084 13268 36136 13320
rect 38292 13311 38344 13320
rect 38292 13277 38301 13311
rect 38301 13277 38335 13311
rect 38335 13277 38344 13311
rect 38292 13268 38344 13277
rect 41144 13268 41196 13320
rect 39948 13200 40000 13252
rect 40132 13200 40184 13252
rect 23112 13132 23164 13184
rect 25596 13132 25648 13184
rect 32312 13132 32364 13184
rect 40040 13175 40092 13184
rect 40040 13141 40049 13175
rect 40049 13141 40083 13175
rect 40083 13141 40092 13175
rect 40040 13132 40092 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 22652 12792 22704 12844
rect 24676 12835 24728 12844
rect 24676 12801 24685 12835
rect 24685 12801 24719 12835
rect 24719 12801 24728 12835
rect 24676 12792 24728 12801
rect 24860 12792 24912 12844
rect 29920 12928 29972 12980
rect 34704 12971 34756 12980
rect 34704 12937 34713 12971
rect 34713 12937 34747 12971
rect 34747 12937 34756 12971
rect 34704 12928 34756 12937
rect 35624 12928 35676 12980
rect 36452 12928 36504 12980
rect 41144 12971 41196 12980
rect 41144 12937 41153 12971
rect 41153 12937 41187 12971
rect 41187 12937 41196 12971
rect 41144 12928 41196 12937
rect 26976 12792 27028 12844
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 29736 12860 29788 12912
rect 31484 12860 31536 12912
rect 29552 12792 29604 12844
rect 30656 12835 30708 12844
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 31576 12792 31628 12844
rect 32404 12792 32456 12844
rect 33048 12860 33100 12912
rect 35348 12860 35400 12912
rect 40040 12903 40092 12912
rect 32772 12835 32824 12844
rect 32772 12801 32806 12835
rect 32806 12801 32824 12835
rect 32772 12792 32824 12801
rect 33968 12792 34020 12844
rect 34152 12792 34204 12844
rect 30564 12767 30616 12776
rect 30564 12733 30573 12767
rect 30573 12733 30607 12767
rect 30607 12733 30616 12767
rect 30564 12724 30616 12733
rect 34704 12792 34756 12844
rect 35624 12835 35676 12844
rect 35624 12801 35633 12835
rect 35633 12801 35667 12835
rect 35667 12801 35676 12835
rect 35624 12792 35676 12801
rect 23664 12656 23716 12708
rect 25688 12656 25740 12708
rect 35808 12724 35860 12776
rect 38292 12835 38344 12844
rect 38292 12801 38301 12835
rect 38301 12801 38335 12835
rect 38335 12801 38344 12835
rect 38292 12792 38344 12801
rect 38660 12835 38712 12844
rect 38660 12801 38669 12835
rect 38669 12801 38703 12835
rect 38703 12801 38712 12835
rect 38660 12792 38712 12801
rect 38936 12835 38988 12844
rect 38936 12801 38945 12835
rect 38945 12801 38979 12835
rect 38979 12801 38988 12835
rect 38936 12792 38988 12801
rect 40040 12869 40074 12903
rect 40074 12869 40092 12903
rect 40040 12860 40092 12869
rect 38476 12767 38528 12776
rect 38476 12733 38485 12767
rect 38485 12733 38519 12767
rect 38519 12733 38528 12767
rect 38476 12724 38528 12733
rect 39764 12767 39816 12776
rect 39764 12733 39773 12767
rect 39773 12733 39807 12767
rect 39807 12733 39816 12767
rect 39764 12724 39816 12733
rect 43168 12767 43220 12776
rect 43168 12733 43177 12767
rect 43177 12733 43211 12767
rect 43211 12733 43220 12767
rect 43168 12724 43220 12733
rect 25136 12588 25188 12640
rect 30472 12588 30524 12640
rect 33876 12631 33928 12640
rect 33876 12597 33885 12631
rect 33885 12597 33919 12631
rect 33919 12597 33928 12631
rect 33876 12588 33928 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 24860 12384 24912 12436
rect 30564 12384 30616 12436
rect 30656 12384 30708 12436
rect 32772 12384 32824 12436
rect 39948 12384 40000 12436
rect 24768 12316 24820 12368
rect 26424 12316 26476 12368
rect 33324 12316 33376 12368
rect 23388 12180 23440 12232
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 31300 12248 31352 12300
rect 32588 12248 32640 12300
rect 25320 12180 25372 12232
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 25688 12223 25740 12232
rect 25688 12189 25697 12223
rect 25697 12189 25731 12223
rect 25731 12189 25740 12223
rect 25688 12180 25740 12189
rect 26608 12180 26660 12232
rect 26792 12223 26844 12232
rect 26792 12189 26801 12223
rect 26801 12189 26835 12223
rect 26835 12189 26844 12223
rect 26792 12180 26844 12189
rect 28816 12180 28868 12232
rect 28632 12112 28684 12164
rect 28908 12112 28960 12164
rect 35716 12248 35768 12300
rect 33876 12180 33928 12232
rect 37556 12180 37608 12232
rect 39764 12180 39816 12232
rect 40132 12112 40184 12164
rect 40592 12112 40644 12164
rect 23112 12087 23164 12096
rect 23112 12053 23121 12087
rect 23121 12053 23155 12087
rect 23155 12053 23164 12087
rect 23112 12044 23164 12053
rect 28816 12087 28868 12096
rect 28816 12053 28825 12087
rect 28825 12053 28859 12087
rect 28859 12053 28868 12087
rect 28816 12044 28868 12053
rect 31208 12087 31260 12096
rect 31208 12053 31217 12087
rect 31217 12053 31251 12087
rect 31251 12053 31260 12087
rect 31208 12044 31260 12053
rect 31300 12087 31352 12096
rect 31300 12053 31309 12087
rect 31309 12053 31343 12087
rect 31343 12053 31352 12087
rect 31300 12044 31352 12053
rect 35532 12087 35584 12096
rect 35532 12053 35541 12087
rect 35541 12053 35575 12087
rect 35575 12053 35584 12087
rect 35532 12044 35584 12053
rect 36084 12044 36136 12096
rect 36544 12044 36596 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 23204 11840 23256 11892
rect 23112 11704 23164 11756
rect 27896 11840 27948 11892
rect 28816 11840 28868 11892
rect 29828 11840 29880 11892
rect 30932 11883 30984 11892
rect 30932 11849 30941 11883
rect 30941 11849 30975 11883
rect 30975 11849 30984 11883
rect 30932 11840 30984 11849
rect 34704 11840 34756 11892
rect 36544 11883 36596 11892
rect 36544 11849 36553 11883
rect 36553 11849 36587 11883
rect 36587 11849 36596 11883
rect 36544 11840 36596 11849
rect 36820 11840 36872 11892
rect 26792 11772 26844 11824
rect 28540 11815 28592 11824
rect 28540 11781 28549 11815
rect 28549 11781 28583 11815
rect 28583 11781 28592 11815
rect 28540 11772 28592 11781
rect 34060 11772 34112 11824
rect 35532 11772 35584 11824
rect 38292 11772 38344 11824
rect 26608 11704 26660 11756
rect 25136 11679 25188 11688
rect 25136 11645 25145 11679
rect 25145 11645 25179 11679
rect 25179 11645 25188 11679
rect 25136 11636 25188 11645
rect 27344 11636 27396 11688
rect 30288 11636 30340 11688
rect 31300 11704 31352 11756
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 34796 11704 34848 11756
rect 38476 11704 38528 11756
rect 39948 11840 40000 11892
rect 40592 11883 40644 11892
rect 40592 11849 40601 11883
rect 40601 11849 40635 11883
rect 40635 11849 40644 11883
rect 40592 11840 40644 11849
rect 40132 11815 40184 11824
rect 40132 11781 40141 11815
rect 40141 11781 40175 11815
rect 40175 11781 40184 11815
rect 40132 11772 40184 11781
rect 38384 11679 38436 11688
rect 38384 11645 38393 11679
rect 38393 11645 38427 11679
rect 38427 11645 38436 11679
rect 38384 11636 38436 11645
rect 40224 11636 40276 11688
rect 43168 11679 43220 11688
rect 43168 11645 43177 11679
rect 43177 11645 43211 11679
rect 43211 11645 43220 11679
rect 43168 11636 43220 11645
rect 22744 11543 22796 11552
rect 22744 11509 22753 11543
rect 22753 11509 22787 11543
rect 22787 11509 22796 11543
rect 22744 11500 22796 11509
rect 24676 11500 24728 11552
rect 25872 11543 25924 11552
rect 25872 11509 25881 11543
rect 25881 11509 25915 11543
rect 25915 11509 25924 11543
rect 25872 11500 25924 11509
rect 28080 11543 28132 11552
rect 28080 11509 28089 11543
rect 28089 11509 28123 11543
rect 28123 11509 28132 11543
rect 28080 11500 28132 11509
rect 30380 11500 30432 11552
rect 37832 11500 37884 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 23204 11339 23256 11348
rect 23204 11305 23213 11339
rect 23213 11305 23247 11339
rect 23247 11305 23256 11339
rect 23204 11296 23256 11305
rect 26792 11296 26844 11348
rect 28816 11296 28868 11348
rect 31300 11296 31352 11348
rect 33968 11296 34020 11348
rect 35624 11296 35676 11348
rect 38476 11296 38528 11348
rect 26148 11160 26200 11212
rect 29000 11160 29052 11212
rect 30104 11203 30156 11212
rect 30104 11169 30113 11203
rect 30113 11169 30147 11203
rect 30147 11169 30156 11203
rect 30104 11160 30156 11169
rect 32404 11203 32456 11212
rect 32404 11169 32413 11203
rect 32413 11169 32447 11203
rect 32447 11169 32456 11203
rect 32404 11160 32456 11169
rect 34796 11160 34848 11212
rect 21916 11092 21968 11144
rect 24676 11092 24728 11144
rect 28080 11092 28132 11144
rect 30380 11135 30432 11144
rect 30380 11101 30414 11135
rect 30414 11101 30432 11135
rect 30380 11092 30432 11101
rect 37556 11135 37608 11144
rect 37556 11101 37565 11135
rect 37565 11101 37599 11135
rect 37599 11101 37608 11135
rect 37556 11092 37608 11101
rect 37832 11135 37884 11144
rect 37832 11101 37866 11135
rect 37866 11101 37884 11135
rect 37832 11092 37884 11101
rect 22744 11024 22796 11076
rect 32864 11024 32916 11076
rect 35164 11067 35216 11076
rect 35164 11033 35198 11067
rect 35198 11033 35216 11067
rect 35164 11024 35216 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 26608 10795 26660 10804
rect 26608 10761 26617 10795
rect 26617 10761 26651 10795
rect 26651 10761 26660 10795
rect 26608 10752 26660 10761
rect 28908 10752 28960 10804
rect 31208 10752 31260 10804
rect 32864 10795 32916 10804
rect 32864 10761 32873 10795
rect 32873 10761 32907 10795
rect 32907 10761 32916 10795
rect 32864 10752 32916 10761
rect 33968 10752 34020 10804
rect 35164 10752 35216 10804
rect 35624 10752 35676 10804
rect 38936 10795 38988 10804
rect 38936 10761 38945 10795
rect 38945 10761 38979 10795
rect 38979 10761 38988 10795
rect 38936 10752 38988 10761
rect 26148 10684 26200 10736
rect 25872 10616 25924 10668
rect 28724 10684 28776 10736
rect 31024 10684 31076 10736
rect 38292 10684 38344 10736
rect 28264 10616 28316 10668
rect 30104 10659 30156 10668
rect 30104 10625 30113 10659
rect 30113 10625 30147 10659
rect 30147 10625 30156 10659
rect 30104 10616 30156 10625
rect 30380 10659 30432 10668
rect 30380 10625 30414 10659
rect 30414 10625 30432 10659
rect 30380 10616 30432 10625
rect 37556 10659 37608 10668
rect 37556 10625 37565 10659
rect 37565 10625 37599 10659
rect 37599 10625 37608 10659
rect 37556 10616 37608 10625
rect 37832 10659 37884 10668
rect 37832 10625 37866 10659
rect 37866 10625 37884 10659
rect 37832 10616 37884 10625
rect 33324 10548 33376 10600
rect 35624 10591 35676 10600
rect 35624 10557 35633 10591
rect 35633 10557 35667 10591
rect 35667 10557 35676 10591
rect 35624 10548 35676 10557
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 28264 10251 28316 10260
rect 28264 10217 28273 10251
rect 28273 10217 28307 10251
rect 28307 10217 28316 10251
rect 28264 10208 28316 10217
rect 30380 10208 30432 10260
rect 37832 10251 37884 10260
rect 37832 10217 37841 10251
rect 37841 10217 37875 10251
rect 37875 10217 37884 10251
rect 37832 10208 37884 10217
rect 28632 10140 28684 10192
rect 28540 10072 28592 10124
rect 30564 10140 30616 10192
rect 30932 10115 30984 10124
rect 30932 10081 30941 10115
rect 30941 10081 30975 10115
rect 30975 10081 30984 10115
rect 30932 10072 30984 10081
rect 35624 10140 35676 10192
rect 36912 10140 36964 10192
rect 38292 10115 38344 10124
rect 38292 10081 38301 10115
rect 38301 10081 38335 10115
rect 38335 10081 38344 10115
rect 38292 10072 38344 10081
rect 38844 10072 38896 10124
rect 28908 10004 28960 10056
rect 31208 10004 31260 10056
rect 38936 10004 38988 10056
rect 43168 9979 43220 9988
rect 43168 9945 43177 9979
rect 43177 9945 43211 9979
rect 43211 9945 43220 9979
rect 43168 9936 43220 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 33784 8440 33836 8492
rect 43996 8372 44048 8424
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 33692 6740 33744 6792
rect 43168 6715 43220 6724
rect 43168 6681 43177 6715
rect 43177 6681 43211 6715
rect 43211 6681 43220 6715
rect 43168 6672 43220 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 42800 5652 42852 5704
rect 43996 5584 44048 5636
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 37004 4088 37056 4140
rect 43168 4063 43220 4072
rect 43168 4029 43177 4063
rect 43177 4029 43211 4063
rect 43211 4029 43220 4063
rect 43168 4020 43220 4029
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 34704 2388 34756 2440
rect 43168 2363 43220 2372
rect 43168 2329 43177 2363
rect 43177 2329 43211 2363
rect 43211 2329 43220 2363
rect 43168 2320 43220 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 2226 44200 2282 45000
rect 5906 44200 5962 45000
rect 9586 44200 9642 45000
rect 13266 44200 13322 45000
rect 16946 44200 17002 45000
rect 20626 44200 20682 45000
rect 24306 44200 24362 45000
rect 27986 44200 28042 45000
rect 31666 44200 31722 45000
rect 35346 44200 35402 45000
rect 39026 44200 39082 45000
rect 42706 44200 42762 45000
rect 2240 42226 2268 44200
rect 5920 42226 5948 44200
rect 9600 44146 9628 44200
rect 9600 44118 9720 44146
rect 7196 42288 7248 42294
rect 7196 42230 7248 42236
rect 2228 42220 2280 42226
rect 2228 42162 2280 42168
rect 5908 42220 5960 42226
rect 5908 42162 5960 42168
rect 5632 42152 5684 42158
rect 5632 42094 5684 42100
rect 7012 42152 7064 42158
rect 7012 42094 7064 42100
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 5540 41608 5592 41614
rect 5540 41550 5592 41556
rect 5552 41206 5580 41550
rect 5540 41200 5592 41206
rect 5540 41142 5592 41148
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 5264 40384 5316 40390
rect 5264 40326 5316 40332
rect 5276 40118 5304 40326
rect 5264 40112 5316 40118
rect 5264 40054 5316 40060
rect 5552 39846 5580 41142
rect 5644 40526 5672 42094
rect 6552 42016 6604 42022
rect 6552 41958 6604 41964
rect 6564 41614 6592 41958
rect 7024 41818 7052 42094
rect 7012 41812 7064 41818
rect 7012 41754 7064 41760
rect 6552 41608 6604 41614
rect 6552 41550 6604 41556
rect 6828 41268 6880 41274
rect 6828 41210 6880 41216
rect 6840 40526 6868 41210
rect 5632 40520 5684 40526
rect 5632 40462 5684 40468
rect 6828 40520 6880 40526
rect 6828 40462 6880 40468
rect 6000 40384 6052 40390
rect 6000 40326 6052 40332
rect 6644 40384 6696 40390
rect 6644 40326 6696 40332
rect 6012 40186 6040 40326
rect 6000 40180 6052 40186
rect 6000 40122 6052 40128
rect 4620 39840 4672 39846
rect 4620 39782 4672 39788
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 6552 39840 6604 39846
rect 6552 39782 6604 39788
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4632 37942 4660 39782
rect 6564 38962 6592 39782
rect 6656 39438 6684 40326
rect 6840 40118 6868 40462
rect 7024 40458 7052 41754
rect 7104 40588 7156 40594
rect 7104 40530 7156 40536
rect 7012 40452 7064 40458
rect 7012 40394 7064 40400
rect 6828 40112 6880 40118
rect 6828 40054 6880 40060
rect 7116 39982 7144 40530
rect 7208 40390 7236 42230
rect 9692 42226 9720 44118
rect 13280 42226 13308 44200
rect 16960 44130 16988 44200
rect 20640 44146 20668 44200
rect 16948 44124 17000 44130
rect 16948 44066 17000 44072
rect 18144 44124 18196 44130
rect 20640 44118 20760 44146
rect 18144 44066 18196 44072
rect 14372 42288 14424 42294
rect 14372 42230 14424 42236
rect 9680 42220 9732 42226
rect 9680 42162 9732 42168
rect 13268 42220 13320 42226
rect 13268 42162 13320 42168
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 9220 42152 9272 42158
rect 9220 42094 9272 42100
rect 10324 42152 10376 42158
rect 10324 42094 10376 42100
rect 13636 42152 13688 42158
rect 13636 42094 13688 42100
rect 9128 41608 9180 41614
rect 9128 41550 9180 41556
rect 9140 41206 9168 41550
rect 9128 41200 9180 41206
rect 9128 41142 9180 41148
rect 8392 41132 8444 41138
rect 8392 41074 8444 41080
rect 7196 40384 7248 40390
rect 7196 40326 7248 40332
rect 7208 40089 7236 40326
rect 8404 40186 8432 41074
rect 9036 40928 9088 40934
rect 9036 40870 9088 40876
rect 8944 40656 8996 40662
rect 8944 40598 8996 40604
rect 8760 40452 8812 40458
rect 8760 40394 8812 40400
rect 8392 40180 8444 40186
rect 8392 40122 8444 40128
rect 7194 40080 7250 40089
rect 7194 40015 7250 40024
rect 7104 39976 7156 39982
rect 7104 39918 7156 39924
rect 6736 39500 6788 39506
rect 6736 39442 6788 39448
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6748 39030 6776 39442
rect 7380 39432 7432 39438
rect 7380 39374 7432 39380
rect 7104 39364 7156 39370
rect 7104 39306 7156 39312
rect 6736 39024 6788 39030
rect 6736 38966 6788 38972
rect 5816 38956 5868 38962
rect 5816 38898 5868 38904
rect 5908 38956 5960 38962
rect 5908 38898 5960 38904
rect 6552 38956 6604 38962
rect 6552 38898 6604 38904
rect 5828 38350 5856 38898
rect 5920 38350 5948 38898
rect 6736 38888 6788 38894
rect 6736 38830 6788 38836
rect 5816 38344 5868 38350
rect 5816 38286 5868 38292
rect 5908 38344 5960 38350
rect 5908 38286 5960 38292
rect 6184 38276 6236 38282
rect 6184 38218 6236 38224
rect 4620 37936 4672 37942
rect 4620 37878 4672 37884
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 37878
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4908 37466 4936 37810
rect 5540 37664 5592 37670
rect 5540 37606 5592 37612
rect 4896 37460 4948 37466
rect 4896 37402 4948 37408
rect 5356 37324 5408 37330
rect 5356 37266 5408 37272
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 34678 4660 36110
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 5000 35834 5028 36042
rect 4988 35828 5040 35834
rect 4988 35770 5040 35776
rect 5368 35630 5396 37266
rect 5552 37194 5580 37606
rect 6196 37330 6224 38218
rect 6184 37324 6236 37330
rect 6184 37266 6236 37272
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5552 36281 5580 37130
rect 5538 36272 5594 36281
rect 5538 36207 5594 36216
rect 5540 36032 5592 36038
rect 5538 36000 5540 36009
rect 5592 36000 5594 36009
rect 5594 35958 5672 35986
rect 5538 35935 5594 35944
rect 5172 35624 5224 35630
rect 5172 35566 5224 35572
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 5448 35624 5500 35630
rect 5448 35566 5500 35572
rect 5184 35222 5212 35566
rect 5172 35216 5224 35222
rect 5172 35158 5224 35164
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5368 33810 5396 35566
rect 5460 35290 5488 35566
rect 5448 35284 5500 35290
rect 5448 35226 5500 35232
rect 5538 35184 5594 35193
rect 5538 35119 5594 35128
rect 5552 35086 5580 35119
rect 5644 35086 5672 35958
rect 5540 35080 5592 35086
rect 5540 35022 5592 35028
rect 5632 35080 5684 35086
rect 5632 35022 5684 35028
rect 5816 34604 5868 34610
rect 5816 34546 5868 34552
rect 5828 34202 5856 34546
rect 5816 34196 5868 34202
rect 5816 34138 5868 34144
rect 5276 33782 5396 33810
rect 5276 33318 5304 33782
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 5264 33312 5316 33318
rect 5264 33254 5316 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4908 32910 4936 33254
rect 4160 32904 4212 32910
rect 4160 32846 4212 32852
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4172 32230 4200 32846
rect 4712 32428 4764 32434
rect 4712 32370 4764 32376
rect 4160 32224 4212 32230
rect 4160 32166 4212 32172
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30870 4660 32166
rect 4724 32026 4752 32370
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 5276 31890 5304 33254
rect 5368 33046 5396 33390
rect 5356 33040 5408 33046
rect 5356 32982 5408 32988
rect 5356 32292 5408 32298
rect 5356 32234 5408 32240
rect 5264 31884 5316 31890
rect 5264 31826 5316 31832
rect 5368 31754 5396 32234
rect 5356 31748 5408 31754
rect 5356 31690 5408 31696
rect 6196 31210 6224 37266
rect 6748 36582 6776 38830
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 7024 38350 7052 38694
rect 7116 38654 7144 39306
rect 7392 38962 7420 39374
rect 8772 39030 8800 40394
rect 8956 39982 8984 40598
rect 9048 40390 9076 40870
rect 9140 40594 9168 41142
rect 9232 41002 9260 42094
rect 9588 41540 9640 41546
rect 9588 41482 9640 41488
rect 9600 41274 9628 41482
rect 10048 41472 10100 41478
rect 10048 41414 10100 41420
rect 9588 41268 9640 41274
rect 9588 41210 9640 41216
rect 10060 41070 10088 41414
rect 10336 41138 10364 42094
rect 12992 42016 13044 42022
rect 12992 41958 13044 41964
rect 13004 41614 13032 41958
rect 12072 41608 12124 41614
rect 12072 41550 12124 41556
rect 12992 41608 13044 41614
rect 12992 41550 13044 41556
rect 10324 41132 10376 41138
rect 10324 41074 10376 41080
rect 11980 41132 12032 41138
rect 11980 41074 12032 41080
rect 10048 41064 10100 41070
rect 10048 41006 10100 41012
rect 9220 40996 9272 41002
rect 9220 40938 9272 40944
rect 9232 40662 9260 40938
rect 9220 40656 9272 40662
rect 9220 40598 9272 40604
rect 9128 40588 9180 40594
rect 9128 40530 9180 40536
rect 9588 40520 9640 40526
rect 9640 40468 9720 40474
rect 9588 40462 9720 40468
rect 9600 40446 9720 40462
rect 9036 40384 9088 40390
rect 9036 40326 9088 40332
rect 9048 40186 9076 40326
rect 9036 40180 9088 40186
rect 9036 40122 9088 40128
rect 9692 40050 9720 40446
rect 9864 40384 9916 40390
rect 9864 40326 9916 40332
rect 9876 40118 9904 40326
rect 10060 40118 10088 41006
rect 9864 40112 9916 40118
rect 9864 40054 9916 40060
rect 10048 40112 10100 40118
rect 10048 40054 10100 40060
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 8944 39976 8996 39982
rect 8944 39918 8996 39924
rect 9956 39976 10008 39982
rect 10336 39953 10364 41074
rect 11704 40928 11756 40934
rect 11704 40870 11756 40876
rect 11716 40458 11744 40870
rect 11704 40452 11756 40458
rect 11704 40394 11756 40400
rect 11992 40186 12020 41074
rect 12084 41002 12112 41550
rect 12164 41268 12216 41274
rect 12164 41210 12216 41216
rect 12072 40996 12124 41002
rect 12072 40938 12124 40944
rect 12084 40526 12112 40938
rect 12176 40730 12204 41210
rect 13648 41070 13676 42094
rect 13740 41478 13768 42162
rect 14280 42016 14332 42022
rect 14280 41958 14332 41964
rect 13728 41472 13780 41478
rect 13728 41414 13780 41420
rect 13636 41064 13688 41070
rect 13636 41006 13688 41012
rect 12164 40724 12216 40730
rect 12164 40666 12216 40672
rect 12072 40520 12124 40526
rect 12072 40462 12124 40468
rect 11980 40180 12032 40186
rect 11980 40122 12032 40128
rect 10692 39976 10744 39982
rect 9956 39918 10008 39924
rect 10322 39944 10378 39953
rect 9968 39506 9996 39918
rect 10322 39879 10378 39888
rect 10690 39944 10692 39953
rect 10744 39944 10746 39953
rect 10690 39879 10746 39888
rect 11796 39840 11848 39846
rect 11796 39782 11848 39788
rect 9956 39500 10008 39506
rect 9956 39442 10008 39448
rect 8760 39024 8812 39030
rect 8760 38966 8812 38972
rect 7380 38956 7432 38962
rect 7380 38898 7432 38904
rect 7288 38752 7340 38758
rect 7288 38694 7340 38700
rect 7116 38626 7236 38654
rect 7208 38350 7236 38626
rect 7012 38344 7064 38350
rect 7012 38286 7064 38292
rect 7196 38344 7248 38350
rect 7196 38286 7248 38292
rect 7024 37942 7052 38286
rect 7012 37936 7064 37942
rect 7012 37878 7064 37884
rect 7024 37262 7052 37878
rect 7208 37874 7236 38286
rect 7196 37868 7248 37874
rect 7196 37810 7248 37816
rect 7300 37754 7328 38694
rect 7208 37726 7328 37754
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 6920 37188 6972 37194
rect 6920 37130 6972 37136
rect 6828 37120 6880 37126
rect 6828 37062 6880 37068
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6748 36378 6776 36518
rect 6736 36372 6788 36378
rect 6736 36314 6788 36320
rect 6644 36032 6696 36038
rect 6644 35974 6696 35980
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6380 33998 6408 34342
rect 6656 34066 6684 35974
rect 6748 35714 6776 36314
rect 6840 36174 6868 37062
rect 6932 36174 6960 37130
rect 7208 36174 7236 37726
rect 7392 37670 7420 38898
rect 8772 38350 8800 38966
rect 9968 38962 9996 39442
rect 10416 39432 10468 39438
rect 10416 39374 10468 39380
rect 11336 39432 11388 39438
rect 11336 39374 11388 39380
rect 10232 39364 10284 39370
rect 10232 39306 10284 39312
rect 9956 38956 10008 38962
rect 9956 38898 10008 38904
rect 9036 38752 9088 38758
rect 9036 38694 9088 38700
rect 7932 38344 7984 38350
rect 7932 38286 7984 38292
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 8760 38344 8812 38350
rect 8760 38286 8812 38292
rect 7840 37868 7892 37874
rect 7840 37810 7892 37816
rect 7380 37664 7432 37670
rect 7380 37606 7432 37612
rect 7852 37194 7880 37810
rect 7944 37330 7972 38286
rect 8128 37874 8156 38286
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 8116 37868 8168 37874
rect 8116 37810 8168 37816
rect 7932 37324 7984 37330
rect 7932 37266 7984 37272
rect 7840 37188 7892 37194
rect 7840 37130 7892 37136
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 6828 36168 6880 36174
rect 6828 36110 6880 36116
rect 6920 36168 6972 36174
rect 6920 36110 6972 36116
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 6840 35834 6868 36110
rect 6828 35828 6880 35834
rect 6828 35770 6880 35776
rect 7208 35766 7236 36110
rect 7196 35760 7248 35766
rect 6748 35686 6868 35714
rect 7196 35702 7248 35708
rect 6644 34060 6696 34066
rect 6644 34002 6696 34008
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6460 33992 6512 33998
rect 6460 33934 6512 33940
rect 6380 33590 6408 33934
rect 6368 33584 6420 33590
rect 6368 33526 6420 33532
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 6288 33114 6316 33458
rect 6276 33108 6328 33114
rect 6276 33050 6328 33056
rect 6276 31748 6328 31754
rect 6276 31690 6328 31696
rect 6184 31204 6236 31210
rect 6184 31146 6236 31152
rect 4620 30864 4672 30870
rect 4620 30806 4672 30812
rect 4632 30326 4660 30806
rect 6288 30734 6316 31690
rect 6472 30802 6500 33934
rect 6736 33924 6788 33930
rect 6736 33866 6788 33872
rect 6644 33448 6696 33454
rect 6644 33390 6696 33396
rect 6656 32570 6684 33390
rect 6748 32910 6776 33866
rect 6840 33522 6868 35686
rect 7012 35556 7064 35562
rect 7012 35498 7064 35504
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6644 32564 6696 32570
rect 6564 32524 6644 32552
rect 6564 31822 6592 32524
rect 6644 32506 6696 32512
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6276 30728 6328 30734
rect 6276 30670 6328 30676
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 4620 30320 4672 30326
rect 4620 30262 4672 30268
rect 4816 30258 4844 30534
rect 5552 30394 5580 30534
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 6932 29866 6960 34342
rect 7024 33998 7052 35498
rect 7104 35488 7156 35494
rect 7104 35430 7156 35436
rect 7116 34610 7144 35430
rect 7104 34604 7156 34610
rect 7104 34546 7156 34552
rect 7116 34134 7144 34546
rect 7104 34128 7156 34134
rect 7104 34070 7156 34076
rect 7012 33992 7064 33998
rect 7064 33940 7144 33946
rect 7012 33934 7144 33940
rect 7024 33918 7144 33934
rect 7012 33856 7064 33862
rect 7012 33798 7064 33804
rect 7024 33522 7052 33798
rect 7012 33516 7064 33522
rect 7012 33458 7064 33464
rect 7024 32978 7052 33458
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 7024 32366 7052 32778
rect 7012 32360 7064 32366
rect 7012 32302 7064 32308
rect 7116 31822 7144 33918
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7024 30938 7052 31758
rect 7208 31278 7236 35702
rect 7300 35086 7328 36518
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 7288 34604 7340 34610
rect 7288 34546 7340 34552
rect 7300 32434 7328 34546
rect 7288 32428 7340 32434
rect 7288 32370 7340 32376
rect 7300 31346 7328 32370
rect 7392 31890 7420 37062
rect 7852 36786 7880 37130
rect 7840 36780 7892 36786
rect 7840 36722 7892 36728
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 7576 36106 7604 36518
rect 7564 36100 7616 36106
rect 7564 36042 7616 36048
rect 7576 35154 7604 36042
rect 7852 35698 7880 36722
rect 7840 35692 7892 35698
rect 7840 35634 7892 35640
rect 7944 35154 7972 37266
rect 8128 37194 8156 37810
rect 8220 37262 8248 38150
rect 9048 37874 9076 38694
rect 10140 38412 10192 38418
rect 10140 38354 10192 38360
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 9036 37868 9088 37874
rect 9036 37810 9088 37816
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 8116 37188 8168 37194
rect 8116 37130 8168 37136
rect 8116 36916 8168 36922
rect 8116 36858 8168 36864
rect 8024 36780 8076 36786
rect 8024 36722 8076 36728
rect 8036 36310 8064 36722
rect 8024 36304 8076 36310
rect 8024 36246 8076 36252
rect 7564 35148 7616 35154
rect 7564 35090 7616 35096
rect 7932 35148 7984 35154
rect 7932 35090 7984 35096
rect 7656 35080 7708 35086
rect 7656 35022 7708 35028
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7576 34678 7604 34886
rect 7564 34672 7616 34678
rect 7564 34614 7616 34620
rect 7564 34468 7616 34474
rect 7564 34410 7616 34416
rect 7472 34400 7524 34406
rect 7472 34342 7524 34348
rect 7484 34202 7512 34342
rect 7472 34196 7524 34202
rect 7472 34138 7524 34144
rect 7576 33386 7604 34410
rect 7564 33380 7616 33386
rect 7564 33322 7616 33328
rect 7576 33114 7604 33322
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7576 32994 7604 33050
rect 7484 32966 7604 32994
rect 7484 31890 7512 32966
rect 7668 32842 7696 35022
rect 7932 35012 7984 35018
rect 7932 34954 7984 34960
rect 7944 33930 7972 34954
rect 7840 33924 7892 33930
rect 7840 33866 7892 33872
rect 7932 33924 7984 33930
rect 7932 33866 7984 33872
rect 7852 33114 7880 33866
rect 7944 33386 7972 33866
rect 8036 33538 8064 36246
rect 8128 36174 8156 36858
rect 8220 36718 8248 37198
rect 8944 36780 8996 36786
rect 8944 36722 8996 36728
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 8852 36644 8904 36650
rect 8852 36586 8904 36592
rect 8116 36168 8168 36174
rect 8116 36110 8168 36116
rect 8128 35494 8156 36110
rect 8864 36106 8892 36586
rect 8852 36100 8904 36106
rect 8852 36042 8904 36048
rect 8300 36032 8352 36038
rect 8300 35974 8352 35980
rect 8576 36032 8628 36038
rect 8576 35974 8628 35980
rect 8208 35828 8260 35834
rect 8312 35816 8340 35974
rect 8260 35788 8340 35816
rect 8208 35770 8260 35776
rect 8392 35556 8444 35562
rect 8392 35498 8444 35504
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8404 34542 8432 35498
rect 8484 35012 8536 35018
rect 8484 34954 8536 34960
rect 8496 34610 8524 34954
rect 8484 34604 8536 34610
rect 8484 34546 8536 34552
rect 8392 34536 8444 34542
rect 8392 34478 8444 34484
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 8128 33658 8156 34138
rect 8116 33652 8168 33658
rect 8116 33594 8168 33600
rect 8036 33510 8156 33538
rect 7932 33380 7984 33386
rect 7932 33322 7984 33328
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 7656 32836 7708 32842
rect 7656 32778 7708 32784
rect 7668 32434 7696 32778
rect 7748 32768 7800 32774
rect 7748 32710 7800 32716
rect 7760 32570 7788 32710
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7656 32428 7708 32434
rect 7656 32370 7708 32376
rect 7564 32360 7616 32366
rect 7564 32302 7616 32308
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7472 31884 7524 31890
rect 7472 31826 7524 31832
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 7196 31272 7248 31278
rect 7116 31220 7196 31226
rect 7116 31214 7248 31220
rect 7116 31198 7236 31214
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 7116 30734 7144 31198
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 6932 29838 7052 29866
rect 6644 29504 6696 29510
rect 6644 29446 6696 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5552 27402 5580 27814
rect 5644 27402 5672 28494
rect 6656 28490 6684 29446
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6828 28552 6880 28558
rect 6932 28540 6960 29106
rect 6880 28512 6960 28540
rect 6828 28494 6880 28500
rect 6644 28484 6696 28490
rect 6644 28426 6696 28432
rect 7024 28218 7052 29838
rect 7116 29714 7144 30670
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 7208 29646 7236 31078
rect 7300 30938 7328 31282
rect 7392 31090 7420 31826
rect 7576 31482 7604 32302
rect 7564 31476 7616 31482
rect 7564 31418 7616 31424
rect 7392 31062 7604 31090
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 7380 30796 7432 30802
rect 7380 30738 7432 30744
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 7392 29578 7420 30738
rect 7484 30394 7512 30874
rect 7576 30666 7604 31062
rect 7564 30660 7616 30666
rect 7564 30602 7616 30608
rect 7472 30388 7524 30394
rect 7472 30330 7524 30336
rect 7944 29594 7972 33322
rect 8128 32910 8156 33510
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8036 32230 8064 32846
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 8024 31952 8076 31958
rect 8024 31894 8076 31900
rect 8036 31414 8064 31894
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8128 30734 8156 31078
rect 8220 30734 8248 31826
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8312 31346 8340 31622
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8404 31226 8432 34478
rect 8496 34066 8524 34546
rect 8588 34066 8616 35974
rect 8864 35698 8892 36042
rect 8956 35834 8984 36722
rect 8944 35828 8996 35834
rect 8944 35770 8996 35776
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8772 35222 8800 35634
rect 8760 35216 8812 35222
rect 8760 35158 8812 35164
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 8576 34060 8628 34066
rect 8576 34002 8628 34008
rect 8772 33538 8800 35158
rect 8864 34542 8892 35634
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8772 33510 8892 33538
rect 8864 33318 8892 33510
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8852 33312 8904 33318
rect 8852 33254 8904 33260
rect 8668 32768 8720 32774
rect 8668 32710 8720 32716
rect 8576 32428 8628 32434
rect 8680 32416 8708 32710
rect 8628 32388 8708 32416
rect 8576 32370 8628 32376
rect 8312 31210 8432 31226
rect 8680 31210 8708 32388
rect 8772 31822 8800 33254
rect 8760 31816 8812 31822
rect 8760 31758 8812 31764
rect 8300 31204 8432 31210
rect 8352 31198 8432 31204
rect 8668 31204 8720 31210
rect 8300 31146 8352 31152
rect 8668 31146 8720 31152
rect 8312 30802 8340 31146
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8772 30734 8800 31758
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 8116 29776 8168 29782
rect 8116 29718 8168 29724
rect 7104 29572 7156 29578
rect 7104 29514 7156 29520
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7840 29572 7892 29578
rect 7944 29566 8064 29594
rect 7840 29514 7892 29520
rect 7116 28694 7144 29514
rect 7104 28688 7156 28694
rect 7104 28630 7156 28636
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7852 28082 7880 29514
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 7944 28762 7972 29106
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 6932 27402 6960 28018
rect 8036 27470 8064 29566
rect 8128 28762 8156 29718
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 8128 28558 8156 28698
rect 8220 28694 8248 29106
rect 8208 28688 8260 28694
rect 8208 28630 8260 28636
rect 8312 28558 8340 29242
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8128 27470 8156 28494
rect 8404 28490 8432 29446
rect 8588 28558 8616 30534
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8956 28082 8984 34682
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 8220 27538 8248 27814
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 5540 27396 5592 27402
rect 5540 27338 5592 27344
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7760 26994 7788 27270
rect 8128 27130 8156 27406
rect 8392 27396 8444 27402
rect 8392 27338 8444 27344
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 8128 26382 8156 27066
rect 8404 26858 8432 27338
rect 9048 26994 9076 37810
rect 9496 37800 9548 37806
rect 9496 37742 9548 37748
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9232 34542 9260 35634
rect 9508 35086 9536 37742
rect 9600 35290 9628 37946
rect 9864 37936 9916 37942
rect 9864 37878 9916 37884
rect 9680 37732 9732 37738
rect 9680 37674 9732 37680
rect 9692 37262 9720 37674
rect 9876 37670 9904 37878
rect 9864 37664 9916 37670
rect 9864 37606 9916 37612
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9692 35698 9720 36722
rect 9772 36644 9824 36650
rect 9772 36586 9824 36592
rect 9784 36174 9812 36586
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 9680 35692 9732 35698
rect 9680 35634 9732 35640
rect 9680 35556 9732 35562
rect 9680 35498 9732 35504
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9496 35080 9548 35086
rect 9496 35022 9548 35028
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9416 34610 9444 34682
rect 9404 34604 9456 34610
rect 9404 34546 9456 34552
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 9416 33998 9444 34546
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9496 33584 9548 33590
rect 9496 33526 9548 33532
rect 9312 33516 9364 33522
rect 9312 33458 9364 33464
rect 9324 33114 9352 33458
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9404 32904 9456 32910
rect 9404 32846 9456 32852
rect 9416 32570 9444 32846
rect 9404 32564 9456 32570
rect 9404 32506 9456 32512
rect 9312 32496 9364 32502
rect 9312 32438 9364 32444
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9232 31414 9260 31622
rect 9324 31482 9352 32438
rect 9508 32434 9536 33526
rect 9600 32502 9628 35226
rect 9692 34678 9720 35498
rect 9784 35018 9812 35770
rect 9772 35012 9824 35018
rect 9772 34954 9824 34960
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 9680 34400 9732 34406
rect 9680 34342 9732 34348
rect 9692 33930 9720 34342
rect 9680 33924 9732 33930
rect 9680 33866 9732 33872
rect 9784 33522 9812 34954
rect 9876 34746 9904 37606
rect 10048 37256 10100 37262
rect 9968 37204 10048 37210
rect 9968 37198 10100 37204
rect 9968 37182 10088 37198
rect 9968 36922 9996 37182
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 9968 36378 9996 36858
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 9956 36372 10008 36378
rect 9956 36314 10008 36320
rect 10060 35766 10088 36654
rect 10048 35760 10100 35766
rect 10048 35702 10100 35708
rect 10152 35698 10180 38354
rect 10244 37942 10272 39306
rect 10428 38962 10456 39374
rect 10416 38956 10468 38962
rect 10416 38898 10468 38904
rect 10232 37936 10284 37942
rect 10232 37878 10284 37884
rect 10244 36786 10272 37878
rect 10428 37874 10456 38898
rect 11152 38344 11204 38350
rect 11152 38286 11204 38292
rect 10416 37868 10468 37874
rect 10416 37810 10468 37816
rect 10508 37868 10560 37874
rect 10508 37810 10560 37816
rect 11060 37868 11112 37874
rect 11060 37810 11112 37816
rect 10324 37256 10376 37262
rect 10322 37224 10324 37233
rect 10376 37224 10378 37233
rect 10322 37159 10378 37168
rect 10428 36786 10456 37810
rect 10520 37738 10548 37810
rect 10692 37800 10744 37806
rect 10692 37742 10744 37748
rect 10508 37732 10560 37738
rect 10508 37674 10560 37680
rect 10704 37670 10732 37742
rect 10692 37664 10744 37670
rect 10692 37606 10744 37612
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 10704 36854 10732 37062
rect 10692 36848 10744 36854
rect 10692 36790 10744 36796
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10416 36780 10468 36786
rect 10416 36722 10468 36728
rect 10508 36712 10560 36718
rect 10508 36654 10560 36660
rect 10520 36310 10548 36654
rect 10876 36576 10928 36582
rect 10876 36518 10928 36524
rect 10968 36576 11020 36582
rect 10968 36518 11020 36524
rect 10888 36417 10916 36518
rect 10874 36408 10930 36417
rect 10874 36343 10930 36352
rect 10232 36304 10284 36310
rect 10232 36246 10284 36252
rect 10508 36304 10560 36310
rect 10508 36246 10560 36252
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9784 32978 9812 33254
rect 9772 32972 9824 32978
rect 9772 32914 9824 32920
rect 9588 32496 9640 32502
rect 9588 32438 9640 32444
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9508 31754 9536 32370
rect 9692 32026 9720 32370
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9876 31822 9904 33798
rect 9968 32842 9996 35634
rect 10244 35086 10272 36246
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 10336 35834 10364 36110
rect 10520 36038 10548 36246
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 10324 35828 10376 35834
rect 10324 35770 10376 35776
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 9956 32836 10008 32842
rect 9956 32778 10008 32784
rect 10060 32774 10088 34546
rect 10324 34536 10376 34542
rect 10324 34478 10376 34484
rect 10232 34468 10284 34474
rect 10232 34410 10284 34416
rect 10244 34066 10272 34410
rect 10336 34066 10364 34478
rect 10232 34060 10284 34066
rect 10232 34002 10284 34008
rect 10324 34060 10376 34066
rect 10324 34002 10376 34008
rect 10244 33658 10272 34002
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10336 33402 10364 34002
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10152 33374 10364 33402
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9416 31726 9536 31754
rect 9312 31476 9364 31482
rect 9312 31418 9364 31424
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 9220 29844 9272 29850
rect 9220 29786 9272 29792
rect 9232 29306 9260 29786
rect 9324 29646 9352 31282
rect 9416 30326 9444 31726
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9508 30802 9536 31418
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9772 30796 9824 30802
rect 9772 30738 9824 30744
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9128 29232 9180 29238
rect 9128 29174 9180 29180
rect 9140 28558 9168 29174
rect 9416 28558 9444 30262
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9140 27470 9168 28494
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 27062 9168 27406
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8392 26852 8444 26858
rect 8392 26794 8444 26800
rect 9036 26512 9088 26518
rect 9036 26454 9088 26460
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 9048 24818 9076 26454
rect 9508 26382 9536 30534
rect 9784 30258 9812 30738
rect 9876 30734 9904 31146
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26382 9720 26726
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 8312 24410 8340 24550
rect 9416 24410 9444 26250
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 10152 24274 10180 33374
rect 10428 33266 10456 33458
rect 10336 33238 10456 33266
rect 10336 32774 10364 33238
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 10324 32768 10376 32774
rect 10324 32710 10376 32716
rect 10336 32230 10364 32710
rect 10324 32224 10376 32230
rect 10324 32166 10376 32172
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10336 31686 10364 31962
rect 10324 31680 10376 31686
rect 10324 31622 10376 31628
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 10244 26926 10272 31418
rect 10428 31346 10456 33050
rect 10520 31346 10548 35974
rect 10600 35692 10652 35698
rect 10600 35634 10652 35640
rect 10612 34678 10640 35634
rect 10980 35562 11008 36518
rect 11072 36310 11100 37810
rect 11164 37398 11192 38286
rect 11152 37392 11204 37398
rect 11152 37334 11204 37340
rect 11348 37194 11376 39374
rect 11808 38962 11836 39782
rect 11888 39364 11940 39370
rect 11888 39306 11940 39312
rect 11796 38956 11848 38962
rect 11796 38898 11848 38904
rect 11428 38820 11480 38826
rect 11428 38762 11480 38768
rect 11440 37806 11468 38762
rect 11428 37800 11480 37806
rect 11428 37742 11480 37748
rect 11336 37188 11388 37194
rect 11336 37130 11388 37136
rect 11060 36304 11112 36310
rect 11060 36246 11112 36252
rect 11072 36174 11100 36246
rect 11348 36174 11376 37130
rect 11440 37074 11468 37742
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11612 37664 11664 37670
rect 11612 37606 11664 37612
rect 11532 37398 11560 37606
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 11624 37262 11652 37606
rect 11704 37460 11756 37466
rect 11704 37402 11756 37408
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 11440 37046 11652 37074
rect 11428 36780 11480 36786
rect 11428 36722 11480 36728
rect 11440 36650 11468 36722
rect 11428 36644 11480 36650
rect 11428 36586 11480 36592
rect 11520 36372 11572 36378
rect 11520 36314 11572 36320
rect 11532 36174 11560 36314
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 11336 36168 11388 36174
rect 11336 36110 11388 36116
rect 11520 36168 11572 36174
rect 11520 36110 11572 36116
rect 11532 36038 11560 36110
rect 11244 36032 11296 36038
rect 11244 35974 11296 35980
rect 11520 36032 11572 36038
rect 11520 35974 11572 35980
rect 10968 35556 11020 35562
rect 10968 35498 11020 35504
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10600 34672 10652 34678
rect 10600 34614 10652 34620
rect 10612 33114 10640 34614
rect 10796 34134 10824 35022
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 10784 34128 10836 34134
rect 10784 34070 10836 34076
rect 10968 34060 11020 34066
rect 10968 34002 11020 34008
rect 10692 33584 10744 33590
rect 10692 33526 10744 33532
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10704 32842 10732 33526
rect 10980 33522 11008 34002
rect 11072 33930 11100 34886
rect 11152 34128 11204 34134
rect 11152 34070 11204 34076
rect 11164 33930 11192 34070
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 11152 33924 11204 33930
rect 11152 33866 11204 33872
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10968 33516 11020 33522
rect 10968 33458 11020 33464
rect 10692 32836 10744 32842
rect 10692 32778 10744 32784
rect 10796 32502 10824 33458
rect 10980 33114 11008 33458
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 11072 32994 11100 33866
rect 11072 32966 11192 32994
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10796 32366 10824 32438
rect 10784 32360 10836 32366
rect 10784 32302 10836 32308
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10612 31482 10640 31758
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10600 31476 10652 31482
rect 10600 31418 10652 31424
rect 10416 31340 10468 31346
rect 10416 31282 10468 31288
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 10428 30802 10456 31282
rect 10704 31226 10732 31622
rect 10520 31198 10732 31226
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10520 30734 10548 31198
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10508 30728 10560 30734
rect 10508 30670 10560 30676
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 10336 27130 10364 27338
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10520 27010 10548 30670
rect 10704 30666 10732 31078
rect 10796 30802 10824 32302
rect 10876 31952 10928 31958
rect 10876 31894 10928 31900
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 10704 30258 10732 30602
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10704 29578 10732 29990
rect 10692 29572 10744 29578
rect 10692 29514 10744 29520
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 27130 10732 27270
rect 10888 27130 10916 31894
rect 10980 30734 11008 32846
rect 11164 32026 11192 32966
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 11256 31958 11284 35974
rect 11624 35698 11652 37046
rect 11716 36378 11744 37402
rect 11808 37126 11836 38898
rect 11900 37262 11928 39306
rect 11980 39296 12032 39302
rect 11980 39238 12032 39244
rect 11992 38282 12020 39238
rect 11980 38276 12032 38282
rect 11980 38218 12032 38224
rect 11992 37466 12020 38218
rect 11980 37460 12032 37466
rect 11980 37402 12032 37408
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 11796 37120 11848 37126
rect 11796 37062 11848 37068
rect 11704 36372 11756 36378
rect 11704 36314 11756 36320
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 11348 33862 11376 34886
rect 11428 34128 11480 34134
rect 11428 34070 11480 34076
rect 11336 33856 11388 33862
rect 11336 33798 11388 33804
rect 11348 32774 11376 33798
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11348 32570 11376 32710
rect 11336 32564 11388 32570
rect 11336 32506 11388 32512
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 11440 31686 11468 34070
rect 11624 32230 11652 35634
rect 11716 35222 11744 36314
rect 11888 36168 11940 36174
rect 11888 36110 11940 36116
rect 11900 35766 11928 36110
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 11992 35834 12020 36042
rect 11980 35828 12032 35834
rect 11980 35770 12032 35776
rect 11888 35760 11940 35766
rect 11888 35702 11940 35708
rect 11704 35216 11756 35222
rect 11756 35164 11836 35170
rect 11704 35158 11836 35164
rect 11716 35142 11836 35158
rect 11808 35086 11836 35142
rect 11704 35080 11756 35086
rect 11704 35022 11756 35028
rect 11796 35080 11848 35086
rect 11796 35022 11848 35028
rect 11716 34610 11744 35022
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 12084 33590 12112 40462
rect 12176 40186 12204 40666
rect 12164 40180 12216 40186
rect 12164 40122 12216 40128
rect 13740 40050 13768 41414
rect 14292 41206 14320 41958
rect 14280 41200 14332 41206
rect 14280 41142 14332 41148
rect 14280 40452 14332 40458
rect 14280 40394 14332 40400
rect 13728 40044 13780 40050
rect 13728 39986 13780 39992
rect 14292 39982 14320 40394
rect 14384 40186 14412 42230
rect 18156 42226 18184 44066
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 20732 42226 20760 44118
rect 23388 42356 23440 42362
rect 23388 42298 23440 42304
rect 14556 42220 14608 42226
rect 14556 42162 14608 42168
rect 15108 42220 15160 42226
rect 15108 42162 15160 42168
rect 17224 42220 17276 42226
rect 17224 42162 17276 42168
rect 18144 42220 18196 42226
rect 18144 42162 18196 42168
rect 20720 42220 20772 42226
rect 20720 42162 20772 42168
rect 14568 42090 14596 42162
rect 14556 42084 14608 42090
rect 14556 42026 14608 42032
rect 14568 41414 14596 42026
rect 14568 41386 14780 41414
rect 14556 41200 14608 41206
rect 14556 41142 14608 41148
rect 14568 40458 14596 41142
rect 14648 40928 14700 40934
rect 14648 40870 14700 40876
rect 14660 40458 14688 40870
rect 14752 40458 14780 41386
rect 15016 40996 15068 41002
rect 15016 40938 15068 40944
rect 14556 40452 14608 40458
rect 14556 40394 14608 40400
rect 14648 40452 14700 40458
rect 14648 40394 14700 40400
rect 14740 40452 14792 40458
rect 14740 40394 14792 40400
rect 14924 40452 14976 40458
rect 14924 40394 14976 40400
rect 14372 40180 14424 40186
rect 14372 40122 14424 40128
rect 12440 39976 12492 39982
rect 12440 39918 12492 39924
rect 14280 39976 14332 39982
rect 14280 39918 14332 39924
rect 12452 38826 12480 39918
rect 14740 39364 14792 39370
rect 14740 39306 14792 39312
rect 12992 39024 13044 39030
rect 12992 38966 13044 38972
rect 12808 38956 12860 38962
rect 12808 38898 12860 38904
rect 12440 38820 12492 38826
rect 12440 38762 12492 38768
rect 12348 38548 12400 38554
rect 12348 38490 12400 38496
rect 12360 37874 12388 38490
rect 12348 37868 12400 37874
rect 12348 37810 12400 37816
rect 12256 37664 12308 37670
rect 12256 37606 12308 37612
rect 12268 37330 12296 37606
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 12176 34134 12204 37198
rect 12360 36922 12388 37810
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12360 36689 12388 36858
rect 12346 36680 12402 36689
rect 12346 36615 12402 36624
rect 12452 36394 12480 38762
rect 12820 38298 12848 38898
rect 12820 38282 12940 38298
rect 12624 38276 12676 38282
rect 12624 38218 12676 38224
rect 12820 38276 12952 38282
rect 12820 38270 12900 38276
rect 12636 38010 12664 38218
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 12532 37188 12584 37194
rect 12532 37130 12584 37136
rect 12360 36366 12480 36394
rect 12360 36020 12388 36366
rect 12544 36174 12572 37130
rect 12636 36786 12664 37946
rect 12820 37874 12848 38270
rect 12900 38218 12952 38224
rect 12808 37868 12860 37874
rect 12808 37810 12860 37816
rect 12716 37732 12768 37738
rect 12716 37674 12768 37680
rect 12728 37398 12756 37674
rect 12716 37392 12768 37398
rect 12716 37334 12768 37340
rect 12820 37210 12848 37810
rect 13004 37670 13032 38966
rect 14004 38956 14056 38962
rect 14004 38898 14056 38904
rect 13084 38888 13136 38894
rect 13084 38830 13136 38836
rect 13096 38214 13124 38830
rect 13452 38344 13504 38350
rect 13452 38286 13504 38292
rect 13084 38208 13136 38214
rect 13084 38150 13136 38156
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 13360 38208 13412 38214
rect 13360 38150 13412 38156
rect 13096 37874 13124 38150
rect 13084 37868 13136 37874
rect 13084 37810 13136 37816
rect 12992 37664 13044 37670
rect 12992 37606 13044 37612
rect 13096 37330 13124 37810
rect 13280 37466 13308 38150
rect 13268 37460 13320 37466
rect 13268 37402 13320 37408
rect 13372 37398 13400 38150
rect 13360 37392 13412 37398
rect 13464 37369 13492 38286
rect 13820 38208 13872 38214
rect 13820 38150 13872 38156
rect 13832 37874 13860 38150
rect 14016 38010 14044 38898
rect 14752 38826 14780 39306
rect 14740 38820 14792 38826
rect 14740 38762 14792 38768
rect 14188 38752 14240 38758
rect 14188 38694 14240 38700
rect 14096 38412 14148 38418
rect 14096 38354 14148 38360
rect 14004 38004 14056 38010
rect 14004 37946 14056 37952
rect 14108 37874 14136 38354
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 14096 37868 14148 37874
rect 14096 37810 14148 37816
rect 13360 37334 13412 37340
rect 13450 37360 13506 37369
rect 13084 37324 13136 37330
rect 13084 37266 13136 37272
rect 13372 37233 13400 37334
rect 13450 37295 13506 37304
rect 13728 37324 13780 37330
rect 13780 37284 13860 37312
rect 13728 37266 13780 37272
rect 12728 37182 12848 37210
rect 13358 37224 13414 37233
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12622 36680 12678 36689
rect 12622 36615 12678 36624
rect 12532 36168 12584 36174
rect 12532 36110 12584 36116
rect 12360 35992 12480 36020
rect 12256 35284 12308 35290
rect 12256 35226 12308 35232
rect 12164 34128 12216 34134
rect 12164 34070 12216 34076
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11716 32366 11744 32846
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11704 32360 11756 32366
rect 11704 32302 11756 32308
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11428 31680 11480 31686
rect 11428 31622 11480 31628
rect 11440 31278 11468 31622
rect 11716 31346 11744 32302
rect 11992 31890 12020 32778
rect 12072 32360 12124 32366
rect 12072 32302 12124 32308
rect 11980 31884 12032 31890
rect 11980 31826 12032 31832
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11428 31272 11480 31278
rect 11428 31214 11480 31220
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 11520 30728 11572 30734
rect 11572 30676 11744 30682
rect 11520 30670 11744 30676
rect 10980 30274 11008 30670
rect 11532 30654 11744 30670
rect 11716 30598 11744 30654
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 10980 30258 11192 30274
rect 10980 30252 11204 30258
rect 10980 30246 11152 30252
rect 11152 30194 11204 30200
rect 11164 28762 11192 30194
rect 11612 30184 11664 30190
rect 11612 30126 11664 30132
rect 11624 30054 11652 30126
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11518 29880 11574 29889
rect 11624 29850 11652 29990
rect 11518 29815 11520 29824
rect 11572 29815 11574 29824
rect 11612 29844 11664 29850
rect 11520 29786 11572 29792
rect 11612 29786 11664 29792
rect 11704 29640 11756 29646
rect 11704 29582 11756 29588
rect 11716 29170 11744 29582
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 11716 27538 11744 29106
rect 12084 28218 12112 32302
rect 12176 30734 12204 33866
rect 12268 33114 12296 35226
rect 12452 34678 12480 35992
rect 12544 35086 12572 36110
rect 12636 35290 12664 36615
rect 12728 36038 12756 37182
rect 13358 37159 13414 37168
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 13636 36780 13688 36786
rect 13636 36722 13688 36728
rect 12992 36576 13044 36582
rect 13096 36564 13124 36722
rect 13648 36689 13676 36722
rect 13634 36680 13690 36689
rect 13634 36615 13690 36624
rect 13096 36536 13216 36564
rect 12992 36518 13044 36524
rect 12808 36304 12860 36310
rect 12808 36246 12860 36252
rect 12716 36032 12768 36038
rect 12716 35974 12768 35980
rect 12728 35766 12756 35974
rect 12820 35834 12848 36246
rect 12900 36168 12952 36174
rect 12900 36110 12952 36116
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 12716 35760 12768 35766
rect 12716 35702 12768 35708
rect 12716 35556 12768 35562
rect 12716 35498 12768 35504
rect 12624 35284 12676 35290
rect 12624 35226 12676 35232
rect 12532 35080 12584 35086
rect 12532 35022 12584 35028
rect 12440 34672 12492 34678
rect 12440 34614 12492 34620
rect 12728 34610 12756 35498
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12256 33108 12308 33114
rect 12256 33050 12308 33056
rect 12256 32904 12308 32910
rect 12256 32846 12308 32852
rect 12268 32298 12296 32846
rect 12728 32570 12756 34546
rect 12912 34474 12940 36110
rect 13004 35698 13032 36518
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 12992 35692 13044 35698
rect 12992 35634 13044 35640
rect 12900 34468 12952 34474
rect 12900 34410 12952 34416
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 12912 33590 12940 33866
rect 12900 33584 12952 33590
rect 12900 33526 12952 33532
rect 13004 33436 13032 35634
rect 13096 34678 13124 36110
rect 13084 34672 13136 34678
rect 13084 34614 13136 34620
rect 13188 34105 13216 36536
rect 13648 36378 13676 36615
rect 13636 36372 13688 36378
rect 13636 36314 13688 36320
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13372 35193 13400 35770
rect 13544 35760 13596 35766
rect 13544 35702 13596 35708
rect 13358 35184 13414 35193
rect 13358 35119 13414 35128
rect 13174 34096 13230 34105
rect 13174 34031 13230 34040
rect 13372 33454 13400 35119
rect 13556 34610 13584 35702
rect 13728 34672 13780 34678
rect 13728 34614 13780 34620
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13544 34468 13596 34474
rect 13544 34410 13596 34416
rect 13556 33522 13584 34410
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13740 33454 13768 34614
rect 13832 34610 13860 37284
rect 14016 36922 14044 37810
rect 14108 37466 14136 37810
rect 14200 37806 14228 38694
rect 14280 38480 14332 38486
rect 14280 38422 14332 38428
rect 14188 37800 14240 37806
rect 14188 37742 14240 37748
rect 14096 37460 14148 37466
rect 14096 37402 14148 37408
rect 14188 37188 14240 37194
rect 14188 37130 14240 37136
rect 14004 36916 14056 36922
rect 14004 36858 14056 36864
rect 14200 36174 14228 37130
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 14292 35494 14320 38422
rect 14752 38350 14780 38762
rect 14832 38752 14884 38758
rect 14832 38694 14884 38700
rect 14740 38344 14792 38350
rect 14740 38286 14792 38292
rect 14752 37754 14780 38286
rect 14844 37874 14872 38694
rect 14832 37868 14884 37874
rect 14832 37810 14884 37816
rect 14752 37726 14872 37754
rect 14372 37664 14424 37670
rect 14372 37606 14424 37612
rect 14384 35630 14412 37606
rect 14740 37460 14792 37466
rect 14740 37402 14792 37408
rect 14464 37256 14516 37262
rect 14464 37198 14516 37204
rect 14476 35766 14504 37198
rect 14648 36780 14700 36786
rect 14648 36722 14700 36728
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 36378 14596 36518
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14660 36242 14688 36722
rect 14752 36718 14780 37402
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 14648 36236 14700 36242
rect 14648 36178 14700 36184
rect 14464 35760 14516 35766
rect 14464 35702 14516 35708
rect 14372 35624 14424 35630
rect 14372 35566 14424 35572
rect 14280 35488 14332 35494
rect 14280 35430 14332 35436
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13832 33998 13860 34546
rect 14292 34406 14320 35430
rect 14384 35154 14412 35566
rect 14372 35148 14424 35154
rect 14372 35090 14424 35096
rect 14280 34400 14332 34406
rect 14280 34342 14332 34348
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 14292 33930 14320 34342
rect 14280 33924 14332 33930
rect 14280 33866 14332 33872
rect 14188 33516 14240 33522
rect 14384 33504 14412 35090
rect 14476 35086 14504 35702
rect 14844 35698 14872 37726
rect 14556 35692 14608 35698
rect 14556 35634 14608 35640
rect 14832 35692 14884 35698
rect 14832 35634 14884 35640
rect 14568 35086 14596 35634
rect 14464 35080 14516 35086
rect 14464 35022 14516 35028
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14476 34542 14504 35022
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14568 33522 14596 35022
rect 14240 33476 14412 33504
rect 14556 33516 14608 33522
rect 14188 33458 14240 33464
rect 14556 33458 14608 33464
rect 12912 33408 13032 33436
rect 13360 33448 13412 33454
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12716 32564 12768 32570
rect 12716 32506 12768 32512
rect 12440 32496 12492 32502
rect 12440 32438 12492 32444
rect 12256 32292 12308 32298
rect 12256 32234 12308 32240
rect 12452 31754 12480 32438
rect 12820 32434 12848 32710
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12820 32314 12848 32370
rect 12728 32286 12848 32314
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12360 29646 12388 30194
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12360 28762 12388 29582
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 12360 28082 12388 28698
rect 12728 28558 12756 32286
rect 12912 31754 12940 33408
rect 13728 33448 13780 33454
rect 13412 33408 13492 33436
rect 13360 33390 13412 33396
rect 12992 33312 13044 33318
rect 12992 33254 13044 33260
rect 12820 31726 12940 31754
rect 12820 31142 12848 31726
rect 12808 31136 12860 31142
rect 12808 31078 12860 31084
rect 12820 29646 12848 31078
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12452 28014 12480 28426
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10520 26982 10732 27010
rect 10980 26994 11008 27406
rect 11716 26994 11744 27474
rect 12164 27396 12216 27402
rect 12164 27338 12216 27344
rect 10232 26920 10284 26926
rect 10232 26862 10284 26868
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 10244 24954 10272 25162
rect 10612 24954 10640 25434
rect 10704 25226 10732 26982
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10888 25430 10916 26862
rect 10980 26450 11008 26930
rect 12176 26586 12204 27338
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26586 12296 26726
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12452 26450 12480 27950
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 12544 27062 12572 27814
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 10692 25220 10744 25226
rect 10692 25162 10744 25168
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10704 24818 10732 25162
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10888 24750 10916 25366
rect 10980 25294 11008 26386
rect 12728 26382 12756 28494
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12636 25974 12664 26182
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 11888 25832 11940 25838
rect 11888 25774 11940 25780
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10888 24274 10916 24686
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 11072 24206 11100 24618
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 9876 23730 9904 24006
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 10244 23662 10272 24006
rect 11072 23798 11100 24142
rect 11716 24138 11744 25094
rect 11900 24750 11928 25774
rect 13004 25294 13032 33254
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 13096 32026 13124 32370
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 13372 31958 13400 32506
rect 13360 31952 13412 31958
rect 13360 31894 13412 31900
rect 13372 31482 13400 31894
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13268 30252 13320 30258
rect 13464 30240 13492 33408
rect 13728 33390 13780 33396
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 13912 33312 13964 33318
rect 13912 33254 13964 33260
rect 13556 32280 13584 33254
rect 13636 32564 13688 32570
rect 13636 32506 13688 32512
rect 13648 32434 13676 32506
rect 13924 32434 13952 33254
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 13636 32428 13688 32434
rect 13636 32370 13688 32376
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 13556 32252 13676 32280
rect 13648 31754 13676 32252
rect 13912 31952 13964 31958
rect 13912 31894 13964 31900
rect 13636 31748 13688 31754
rect 13636 31690 13688 31696
rect 13820 31680 13872 31686
rect 13820 31622 13872 31628
rect 13832 31142 13860 31622
rect 13924 31414 13952 31894
rect 14200 31890 14228 32710
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14292 31890 14320 32302
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 13912 31408 13964 31414
rect 13912 31350 13964 31356
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13832 30326 13860 31078
rect 13820 30320 13872 30326
rect 13820 30262 13872 30268
rect 13924 30258 13952 31350
rect 13320 30212 13492 30240
rect 13912 30252 13964 30258
rect 13268 30194 13320 30200
rect 14200 30240 14228 31826
rect 14292 30734 14320 31826
rect 14568 31822 14596 32166
rect 14556 31816 14608 31822
rect 14556 31758 14608 31764
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 14476 30326 14504 30534
rect 14660 30394 14688 30602
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14464 30320 14516 30326
rect 14464 30262 14516 30268
rect 14372 30252 14424 30258
rect 14200 30212 14372 30240
rect 13912 30194 13964 30200
rect 14372 30194 14424 30200
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 13188 29102 13216 30058
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13096 26790 13124 27270
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 26314 13124 26726
rect 13280 26518 13308 30194
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13372 28490 13400 29446
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13648 28762 13676 29106
rect 14004 28960 14056 28966
rect 14004 28902 14056 28908
rect 13636 28756 13688 28762
rect 13636 28698 13688 28704
rect 14016 28558 14044 28902
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13372 28082 13400 28426
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 11900 24206 11928 24686
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 12728 24070 12756 25230
rect 13372 25226 13400 28018
rect 13464 27130 13492 28086
rect 13832 27946 13860 28426
rect 14292 28218 14320 28494
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 13820 27940 13872 27946
rect 13820 27882 13872 27888
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13464 26926 13492 27066
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 14384 25294 14412 30194
rect 14464 29028 14516 29034
rect 14464 28970 14516 28976
rect 14476 28626 14504 28970
rect 14648 28960 14700 28966
rect 14752 28914 14780 32370
rect 14700 28908 14780 28914
rect 14648 28902 14780 28908
rect 14660 28886 14780 28902
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14752 28558 14780 28886
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14464 28484 14516 28490
rect 14464 28426 14516 28432
rect 14476 28082 14504 28426
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14752 26994 14780 28494
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14844 28150 14872 28358
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14936 27130 14964 40394
rect 15028 36922 15056 40938
rect 15120 40934 15148 42162
rect 16580 42016 16632 42022
rect 16580 41958 16632 41964
rect 16592 41614 16620 41958
rect 16580 41608 16632 41614
rect 16580 41550 16632 41556
rect 17132 41608 17184 41614
rect 17132 41550 17184 41556
rect 15844 41132 15896 41138
rect 15844 41074 15896 41080
rect 15108 40928 15160 40934
rect 15108 40870 15160 40876
rect 15856 40730 15884 41074
rect 16488 41064 16540 41070
rect 16488 41006 16540 41012
rect 15200 40724 15252 40730
rect 15200 40666 15252 40672
rect 15844 40724 15896 40730
rect 15844 40666 15896 40672
rect 15108 40656 15160 40662
rect 15108 40598 15160 40604
rect 15120 38962 15148 40598
rect 15108 38956 15160 38962
rect 15108 38898 15160 38904
rect 15120 38418 15148 38898
rect 15108 38412 15160 38418
rect 15108 38354 15160 38360
rect 15108 37732 15160 37738
rect 15108 37674 15160 37680
rect 15016 36916 15068 36922
rect 15016 36858 15068 36864
rect 15120 36582 15148 37674
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 15108 36576 15160 36582
rect 15108 36518 15160 36524
rect 15028 36106 15056 36518
rect 15120 36174 15148 36518
rect 15108 36168 15160 36174
rect 15108 36110 15160 36116
rect 15016 36100 15068 36106
rect 15016 36042 15068 36048
rect 15212 35834 15240 40666
rect 16500 39438 16528 41006
rect 17144 41002 17172 41550
rect 17236 41206 17264 42162
rect 17316 42152 17368 42158
rect 17316 42094 17368 42100
rect 17776 42152 17828 42158
rect 17776 42094 17828 42100
rect 18696 42152 18748 42158
rect 18696 42094 18748 42100
rect 17328 41478 17356 42094
rect 17408 41540 17460 41546
rect 17408 41482 17460 41488
rect 17316 41472 17368 41478
rect 17316 41414 17368 41420
rect 17224 41200 17276 41206
rect 17224 41142 17276 41148
rect 17132 40996 17184 41002
rect 17132 40938 17184 40944
rect 17144 40610 17172 40938
rect 17144 40594 17264 40610
rect 17144 40588 17276 40594
rect 17144 40582 17224 40588
rect 17224 40530 17276 40536
rect 17132 40520 17184 40526
rect 17132 40462 17184 40468
rect 17144 39914 17172 40462
rect 17132 39908 17184 39914
rect 17132 39850 17184 39856
rect 16856 39500 16908 39506
rect 16856 39442 16908 39448
rect 15752 39432 15804 39438
rect 15752 39374 15804 39380
rect 16488 39432 16540 39438
rect 16488 39374 16540 39380
rect 15764 37738 15792 39374
rect 16304 39296 16356 39302
rect 16304 39238 16356 39244
rect 16316 38826 16344 39238
rect 16304 38820 16356 38826
rect 16304 38762 16356 38768
rect 16500 38457 16528 39374
rect 16868 38962 16896 39442
rect 16948 39364 17000 39370
rect 16948 39306 17000 39312
rect 16960 39098 16988 39306
rect 16948 39092 17000 39098
rect 16948 39034 17000 39040
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16580 38888 16632 38894
rect 16580 38830 16632 38836
rect 16486 38448 16542 38457
rect 16486 38383 16542 38392
rect 16396 38344 16448 38350
rect 16396 38286 16448 38292
rect 16488 38344 16540 38350
rect 16488 38286 16540 38292
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 15752 37732 15804 37738
rect 15752 37674 15804 37680
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15580 36786 15608 37130
rect 15764 37126 15792 37674
rect 15948 37330 15976 37810
rect 16304 37664 16356 37670
rect 16304 37606 16356 37612
rect 15936 37324 15988 37330
rect 15936 37266 15988 37272
rect 15752 37120 15804 37126
rect 15752 37062 15804 37068
rect 15476 36780 15528 36786
rect 15476 36722 15528 36728
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15488 36689 15516 36722
rect 15474 36680 15530 36689
rect 15474 36615 15530 36624
rect 15752 36644 15804 36650
rect 15752 36586 15804 36592
rect 15844 36644 15896 36650
rect 15844 36586 15896 36592
rect 15568 36576 15620 36582
rect 15568 36518 15620 36524
rect 15580 36310 15608 36518
rect 15658 36408 15714 36417
rect 15658 36343 15714 36352
rect 15672 36310 15700 36343
rect 15568 36304 15620 36310
rect 15568 36246 15620 36252
rect 15660 36304 15712 36310
rect 15660 36246 15712 36252
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15764 35698 15792 36586
rect 15856 36378 15884 36586
rect 15844 36372 15896 36378
rect 15844 36314 15896 36320
rect 15948 36310 15976 37266
rect 16316 36689 16344 37606
rect 16302 36680 16358 36689
rect 16302 36615 16358 36624
rect 16408 36582 16436 38286
rect 16500 37806 16528 38286
rect 16592 37874 16620 38830
rect 16868 38418 16896 38898
rect 16856 38412 16908 38418
rect 16856 38354 16908 38360
rect 17132 38412 17184 38418
rect 17132 38354 17184 38360
rect 16856 38276 16908 38282
rect 16856 38218 16908 38224
rect 16672 38208 16724 38214
rect 16672 38150 16724 38156
rect 16684 37942 16712 38150
rect 16672 37936 16724 37942
rect 16672 37878 16724 37884
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16868 37856 16896 38218
rect 16948 37868 17000 37874
rect 16868 37828 16948 37856
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16500 36854 16528 37742
rect 16592 36854 16620 37810
rect 16764 37664 16816 37670
rect 16764 37606 16816 37612
rect 16776 37262 16804 37606
rect 16764 37256 16816 37262
rect 16764 37198 16816 37204
rect 16488 36848 16540 36854
rect 16488 36790 16540 36796
rect 16580 36848 16632 36854
rect 16580 36790 16632 36796
rect 16868 36786 16896 37828
rect 16948 37810 17000 37816
rect 17144 37330 17172 38354
rect 17132 37324 17184 37330
rect 16960 37284 17132 37312
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 16396 36576 16448 36582
rect 16396 36518 16448 36524
rect 16028 36372 16080 36378
rect 16028 36314 16080 36320
rect 15936 36304 15988 36310
rect 15936 36246 15988 36252
rect 16040 35834 16068 36314
rect 16960 36174 16988 37284
rect 17132 37266 17184 37272
rect 17038 37224 17094 37233
rect 17038 37159 17040 37168
rect 17092 37159 17094 37168
rect 17040 37130 17092 37136
rect 17132 36916 17184 36922
rect 17132 36858 17184 36864
rect 17040 36780 17092 36786
rect 17040 36722 17092 36728
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 16028 35828 16080 35834
rect 16028 35770 16080 35776
rect 16960 35698 16988 36110
rect 17052 36020 17080 36722
rect 17144 36378 17172 36858
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17132 36032 17184 36038
rect 17052 35992 17132 36020
rect 17132 35974 17184 35980
rect 17040 35760 17092 35766
rect 17040 35702 17092 35708
rect 15384 35692 15436 35698
rect 15384 35634 15436 35640
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 16948 35692 17000 35698
rect 16948 35634 17000 35640
rect 15396 34950 15424 35634
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15672 35290 15700 35566
rect 15660 35284 15712 35290
rect 15660 35226 15712 35232
rect 15476 35012 15528 35018
rect 15476 34954 15528 34960
rect 15384 34944 15436 34950
rect 15384 34886 15436 34892
rect 15488 34542 15516 34954
rect 17052 34678 17080 35702
rect 17144 35698 17172 35974
rect 17132 35692 17184 35698
rect 17132 35634 17184 35640
rect 17236 35018 17264 40530
rect 17420 39098 17448 41482
rect 17592 41472 17644 41478
rect 17592 41414 17644 41420
rect 17604 41274 17632 41414
rect 17592 41268 17644 41274
rect 17592 41210 17644 41216
rect 17788 40050 17816 42094
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 18052 41132 18104 41138
rect 18052 41074 18104 41080
rect 17972 40662 18000 41074
rect 17960 40656 18012 40662
rect 17960 40598 18012 40604
rect 17776 40044 17828 40050
rect 17776 39986 17828 39992
rect 17684 39500 17736 39506
rect 17684 39442 17736 39448
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 17696 38350 17724 39442
rect 17972 39438 18000 40598
rect 17960 39432 18012 39438
rect 17960 39374 18012 39380
rect 18064 39302 18092 41074
rect 18420 41064 18472 41070
rect 18420 41006 18472 41012
rect 18236 40112 18288 40118
rect 18236 40054 18288 40060
rect 18248 39914 18276 40054
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 18236 39908 18288 39914
rect 18236 39850 18288 39856
rect 18340 39642 18368 39918
rect 18328 39636 18380 39642
rect 18328 39578 18380 39584
rect 18432 39438 18460 41006
rect 18708 40934 18736 42094
rect 23400 41614 23428 42298
rect 24320 42226 24348 44200
rect 28000 42226 28028 44200
rect 31680 44146 31708 44200
rect 31680 44118 31800 44146
rect 31772 42294 31800 44118
rect 35360 42294 35388 44200
rect 28356 42288 28408 42294
rect 28356 42230 28408 42236
rect 31760 42288 31812 42294
rect 31760 42230 31812 42236
rect 35348 42288 35400 42294
rect 35348 42230 35400 42236
rect 24308 42220 24360 42226
rect 24308 42162 24360 42168
rect 27252 42220 27304 42226
rect 27252 42162 27304 42168
rect 27988 42220 28040 42226
rect 27988 42162 28040 42168
rect 24952 42152 25004 42158
rect 24952 42094 25004 42100
rect 20260 41608 20312 41614
rect 20260 41550 20312 41556
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 23388 41608 23440 41614
rect 23388 41550 23440 41556
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19984 41200 20036 41206
rect 19984 41142 20036 41148
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18420 39432 18472 39438
rect 18708 39409 18736 40870
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 18880 39840 18932 39846
rect 18880 39782 18932 39788
rect 18420 39374 18472 39380
rect 18694 39400 18750 39409
rect 18694 39335 18750 39344
rect 18052 39296 18104 39302
rect 18052 39238 18104 39244
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17972 37874 18000 38490
rect 18064 37874 18092 39238
rect 18892 38962 18920 39782
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19996 38962 20024 41142
rect 20272 40526 20300 41550
rect 20352 41200 20404 41206
rect 20352 41142 20404 41148
rect 20364 40730 20392 41142
rect 21100 40934 21128 41550
rect 21180 41540 21232 41546
rect 21180 41482 21232 41488
rect 22284 41540 22336 41546
rect 22284 41482 22336 41488
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 20352 40724 20404 40730
rect 20352 40666 20404 40672
rect 21100 40594 21128 40870
rect 21088 40588 21140 40594
rect 21088 40530 21140 40536
rect 20260 40520 20312 40526
rect 20260 40462 20312 40468
rect 20272 40118 20300 40462
rect 20260 40112 20312 40118
rect 20260 40054 20312 40060
rect 21192 39642 21220 41482
rect 22296 41274 22324 41482
rect 22560 41472 22612 41478
rect 22560 41414 22612 41420
rect 22284 41268 22336 41274
rect 22284 41210 22336 41216
rect 22284 41132 22336 41138
rect 22284 41074 22336 41080
rect 22296 40610 22324 41074
rect 22468 40724 22520 40730
rect 22468 40666 22520 40672
rect 22296 40594 22416 40610
rect 22284 40588 22416 40594
rect 22336 40582 22416 40588
rect 22284 40530 22336 40536
rect 21548 40520 21600 40526
rect 21548 40462 21600 40468
rect 21180 39636 21232 39642
rect 21180 39578 21232 39584
rect 20168 39568 20220 39574
rect 20168 39510 20220 39516
rect 20076 39432 20128 39438
rect 20076 39374 20128 39380
rect 20088 39098 20116 39374
rect 20076 39092 20128 39098
rect 20076 39034 20128 39040
rect 18788 38956 18840 38962
rect 18788 38898 18840 38904
rect 18880 38956 18932 38962
rect 18880 38898 18932 38904
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 18326 38448 18382 38457
rect 18326 38383 18382 38392
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 18052 37868 18104 37874
rect 18052 37810 18104 37816
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 17696 36378 17724 37198
rect 17868 36848 17920 36854
rect 17868 36790 17920 36796
rect 17776 36712 17828 36718
rect 17776 36654 17828 36660
rect 17788 36378 17816 36654
rect 17880 36378 17908 36790
rect 17684 36372 17736 36378
rect 17684 36314 17736 36320
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17868 36372 17920 36378
rect 17868 36314 17920 36320
rect 17880 36258 17908 36314
rect 17316 36236 17368 36242
rect 17316 36178 17368 36184
rect 17604 36230 17908 36258
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 17040 34672 17092 34678
rect 17040 34614 17092 34620
rect 15476 34536 15528 34542
rect 15476 34478 15528 34484
rect 15108 33856 15160 33862
rect 15108 33798 15160 33804
rect 15120 32978 15148 33798
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15488 32842 15516 34478
rect 16948 33992 17000 33998
rect 16948 33934 17000 33940
rect 16960 33522 16988 33934
rect 16948 33516 17000 33522
rect 17052 33504 17080 34614
rect 17236 34610 17264 34954
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17132 33516 17184 33522
rect 17052 33476 17132 33504
rect 16948 33458 17000 33464
rect 17132 33458 17184 33464
rect 16488 33380 16540 33386
rect 16488 33322 16540 33328
rect 16500 32910 16528 33322
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 15476 32836 15528 32842
rect 15476 32778 15528 32784
rect 16408 32570 16436 32846
rect 16396 32564 16448 32570
rect 16396 32506 16448 32512
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16304 32224 16356 32230
rect 16304 32166 16356 32172
rect 16224 32026 16252 32166
rect 16212 32020 16264 32026
rect 16212 31962 16264 31968
rect 16316 31958 16344 32166
rect 16304 31952 16356 31958
rect 16304 31894 16356 31900
rect 17328 31754 17356 36178
rect 17604 36009 17632 36230
rect 17684 36168 17736 36174
rect 17960 36168 18012 36174
rect 17736 36128 17960 36156
rect 17684 36110 17736 36116
rect 17960 36110 18012 36116
rect 17590 36000 17646 36009
rect 17590 35935 17646 35944
rect 17500 35012 17552 35018
rect 17500 34954 17552 34960
rect 17512 33930 17540 34954
rect 17408 33924 17460 33930
rect 17408 33866 17460 33872
rect 17500 33924 17552 33930
rect 17500 33866 17552 33872
rect 17420 33114 17448 33866
rect 17512 33590 17540 33866
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17328 31726 17448 31754
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 14924 27124 14976 27130
rect 14924 27066 14976 27072
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 15028 25294 15056 31078
rect 15936 30592 15988 30598
rect 15936 30534 15988 30540
rect 15948 30190 15976 30534
rect 15936 30184 15988 30190
rect 15936 30126 15988 30132
rect 15948 29170 15976 30126
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 16212 29504 16264 29510
rect 16212 29446 16264 29452
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15212 28082 15240 28494
rect 16224 28490 16252 29446
rect 16592 28694 16620 29446
rect 16868 29306 16896 29446
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 17236 29238 17264 29786
rect 17224 29232 17276 29238
rect 17222 29200 17224 29209
rect 17276 29200 17278 29209
rect 17222 29135 17278 29144
rect 17420 29102 17448 31726
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 16580 28688 16632 28694
rect 16580 28630 16632 28636
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 17328 28218 17356 29038
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16500 27062 16528 27406
rect 16488 27056 16540 27062
rect 16488 26998 16540 27004
rect 16592 26790 16620 27406
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15212 25906 15240 26318
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15212 25294 15240 25842
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24886 12848 25094
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 13924 24614 13952 25230
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14752 24818 14780 25094
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13924 24342 13952 24550
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 11072 23338 11100 23734
rect 10980 23322 11100 23338
rect 10968 23316 11100 23322
rect 11020 23310 11100 23316
rect 10968 23258 11020 23264
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 10704 22030 10732 23122
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 11992 20942 12020 21966
rect 12084 21554 12112 22918
rect 12268 21894 12296 22986
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12176 21486 12204 21830
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 13280 21418 13308 21966
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13372 21146 13400 22034
rect 13556 21486 13584 22578
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13648 22234 13676 22510
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 14568 21876 14596 24346
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14752 23866 14780 24142
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15120 22778 15148 25162
rect 15764 24682 15792 26318
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15856 26042 15884 26250
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15856 24614 15884 25094
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 14648 21888 14700 21894
rect 14568 21848 14648 21876
rect 14648 21830 14700 21836
rect 14660 21554 14688 21830
rect 15028 21554 15056 21898
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15120 21554 15148 21830
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 11992 19378 12020 20878
rect 13280 20602 13308 20878
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 13740 19242 13768 21354
rect 14660 21078 14688 21490
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 15120 20942 15148 21490
rect 15212 21486 15240 21966
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20602 14780 20742
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 20058 14136 20402
rect 14936 20398 14964 20878
rect 15120 20466 15148 20878
rect 15212 20466 15240 20878
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14568 19786 14596 20334
rect 15304 20330 15332 20878
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15396 20058 15424 24210
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 14292 18970 14320 19246
rect 14568 19174 14596 19722
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14568 18766 14596 19110
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14844 18630 14872 19790
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 18698 14964 19314
rect 15120 18766 15148 19450
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14936 18290 14964 18634
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 14936 17814 14964 18226
rect 15212 17882 15240 18226
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 15304 17678 15332 19110
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 17542 15332 17614
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15396 17338 15424 19994
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15488 18426 15516 19858
rect 15764 19446 15792 21286
rect 16040 19922 16068 23054
rect 16224 21690 16252 23598
rect 16684 22094 16712 27950
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16868 25838 16896 26726
rect 16960 26489 16988 26930
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 16946 26480 17002 26489
rect 17052 26450 17080 26862
rect 16946 26415 16948 26424
rect 17000 26415 17002 26424
rect 17040 26444 17092 26450
rect 16948 26386 17000 26392
rect 17040 26386 17092 26392
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 17052 25294 17080 26386
rect 17144 26382 17172 27270
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17236 27033 17264 27066
rect 17222 27024 17278 27033
rect 17222 26959 17278 26968
rect 17420 26926 17448 29038
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17408 26920 17460 26926
rect 17408 26862 17460 26868
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17328 26314 17356 26862
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17420 26586 17448 26726
rect 17512 26586 17540 33526
rect 17604 30802 17632 35935
rect 17868 35692 17920 35698
rect 17972 35680 18000 36110
rect 18144 35760 18196 35766
rect 18144 35702 18196 35708
rect 18052 35692 18104 35698
rect 17972 35652 18052 35680
rect 17868 35634 17920 35640
rect 18052 35634 18104 35640
rect 17880 35290 17908 35634
rect 17868 35284 17920 35290
rect 18156 35272 18184 35702
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 17868 35226 17920 35232
rect 17972 35244 18184 35272
rect 17972 34746 18000 35244
rect 17960 34740 18012 34746
rect 17960 34682 18012 34688
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17880 32842 17908 33798
rect 17868 32836 17920 32842
rect 17868 32778 17920 32784
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17604 29646 17632 30534
rect 17972 30258 18000 34682
rect 18248 34678 18276 35430
rect 18236 34672 18288 34678
rect 18236 34614 18288 34620
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18064 32978 18092 33050
rect 18052 32972 18104 32978
rect 18052 32914 18104 32920
rect 18340 32910 18368 38383
rect 18696 38344 18748 38350
rect 18800 38332 18828 38898
rect 18878 38448 18934 38457
rect 18878 38383 18934 38392
rect 18892 38350 18920 38383
rect 18748 38304 18828 38332
rect 18880 38344 18932 38350
rect 18696 38286 18748 38292
rect 18880 38286 18932 38292
rect 18708 38010 18736 38286
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19352 38010 19380 38150
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19444 37942 19472 38898
rect 19536 38554 19564 38898
rect 19798 38584 19854 38593
rect 19524 38548 19576 38554
rect 19798 38519 19854 38528
rect 19892 38548 19944 38554
rect 19524 38490 19576 38496
rect 19812 38350 19840 38519
rect 19892 38490 19944 38496
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 19800 38344 19852 38350
rect 19800 38286 19852 38292
rect 19904 38282 19932 38490
rect 19892 38276 19944 38282
rect 19892 38218 19944 38224
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 19892 37868 19944 37874
rect 19996 37856 20024 38490
rect 20076 38276 20128 38282
rect 20076 38218 20128 38224
rect 19944 37828 20024 37856
rect 19892 37810 19944 37816
rect 19154 37360 19210 37369
rect 19154 37295 19210 37304
rect 19168 36786 19196 37295
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 18880 36644 18932 36650
rect 18880 36586 18932 36592
rect 18510 36272 18566 36281
rect 18510 36207 18566 36216
rect 18524 36174 18552 36207
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18892 35698 18920 36586
rect 19064 36372 19116 36378
rect 19064 36314 19116 36320
rect 19076 36174 19104 36314
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18696 33108 18748 33114
rect 18696 33050 18748 33056
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18156 31822 18184 32370
rect 18340 32366 18368 32846
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18432 32366 18460 32710
rect 18328 32360 18380 32366
rect 18328 32302 18380 32308
rect 18420 32360 18472 32366
rect 18420 32302 18472 32308
rect 18144 31816 18196 31822
rect 18144 31758 18196 31764
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18248 30666 18276 31282
rect 18340 30802 18368 32302
rect 18708 31754 18736 33050
rect 18616 31726 18736 31754
rect 18328 30796 18380 30802
rect 18328 30738 18380 30744
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 18248 30054 18276 30602
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 29714 18276 29990
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17776 29640 17828 29646
rect 17828 29600 18000 29628
rect 17776 29582 17828 29588
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17592 29096 17644 29102
rect 17592 29038 17644 29044
rect 17604 27470 17632 29038
rect 17880 29034 17908 29106
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 17972 28506 18000 29600
rect 18064 29306 18092 29650
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 18144 28552 18196 28558
rect 17972 28478 18092 28506
rect 18144 28494 18196 28500
rect 17684 28416 17736 28422
rect 17684 28358 17736 28364
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17696 28218 17724 28358
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 17972 27606 18000 28358
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 18064 27130 18092 28478
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17684 26852 17736 26858
rect 17684 26794 17736 26800
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17512 25974 17540 26522
rect 17696 26382 17724 26794
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 17774 26480 17830 26489
rect 17774 26415 17830 26424
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17500 25968 17552 25974
rect 17500 25910 17552 25916
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17328 24954 17356 25230
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16868 24206 16896 24686
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16868 23186 16896 24142
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 22642 16804 22986
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16684 22066 16804 22094
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16132 20942 16160 21490
rect 16224 20942 16252 21626
rect 16776 21146 16804 22066
rect 16868 21486 16896 23122
rect 16960 22778 16988 23598
rect 17328 23322 17356 24890
rect 17512 24886 17540 25910
rect 17788 25226 17816 26415
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 25770 17908 26250
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 18064 25158 18092 26726
rect 18156 26246 18184 28494
rect 18248 28014 18276 29446
rect 18432 29170 18460 30126
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18432 28626 18460 29106
rect 18524 28762 18552 29106
rect 18512 28756 18564 28762
rect 18512 28698 18564 28704
rect 18420 28620 18472 28626
rect 18420 28562 18472 28568
rect 18432 28218 18460 28562
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18340 26518 18368 27066
rect 18432 26994 18460 28154
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18328 26512 18380 26518
rect 18432 26489 18460 26930
rect 18328 26454 18380 26460
rect 18418 26480 18474 26489
rect 18418 26415 18474 26424
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18156 25974 18184 26182
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 18236 25764 18288 25770
rect 18236 25706 18288 25712
rect 18248 25294 18276 25706
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 18064 22710 18092 23462
rect 18340 23100 18368 26250
rect 18156 23072 18368 23100
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 17052 22098 17080 22510
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15764 18766 15792 19382
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15856 18970 15884 19246
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 16684 18698 16712 21014
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15580 17066 15608 17614
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 16040 17202 16068 17546
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 16224 16998 16252 17138
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 16868 15026 16896 21422
rect 17144 21146 17172 21422
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17144 20602 17172 20946
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17236 19446 17264 22374
rect 17328 22030 17356 22374
rect 18156 22094 18184 23072
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18064 22066 18184 22094
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16960 18766 16988 19314
rect 17236 19174 17264 19382
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 16960 17678 16988 18090
rect 17328 17678 17356 18702
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18358 18000 18566
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 16960 16590 16988 17614
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17144 17202 17172 17546
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17328 16794 17356 17614
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17604 16794 17632 17070
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17788 16590 17816 17750
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 18064 15162 18092 22066
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 20058 18184 20334
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18340 19990 18368 22578
rect 18420 21344 18472 21350
rect 18524 21332 18552 28358
rect 18616 26353 18644 31726
rect 18880 30592 18932 30598
rect 18880 30534 18932 30540
rect 18892 30326 18920 30534
rect 18880 30320 18932 30326
rect 18880 30262 18932 30268
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18786 29880 18842 29889
rect 18786 29815 18788 29824
rect 18840 29815 18842 29824
rect 18788 29786 18840 29792
rect 18984 29714 19012 30194
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 19076 29034 19104 36110
rect 19168 34542 19196 36722
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19444 36174 19472 36654
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19904 36174 19932 36314
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19156 34536 19208 34542
rect 19156 34478 19208 34484
rect 19168 33114 19196 34478
rect 19248 33924 19300 33930
rect 19248 33866 19300 33872
rect 19260 33454 19288 33866
rect 19248 33448 19300 33454
rect 19248 33390 19300 33396
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19260 32434 19288 33390
rect 19352 33114 19380 35770
rect 19444 34626 19472 36110
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19892 35828 19944 35834
rect 19892 35770 19944 35776
rect 19904 35222 19932 35770
rect 19996 35714 20024 37828
rect 20088 35834 20116 38218
rect 20180 37874 20208 39510
rect 20812 39432 20864 39438
rect 20812 39374 20864 39380
rect 21088 39432 21140 39438
rect 21088 39374 21140 39380
rect 20260 39296 20312 39302
rect 20260 39238 20312 39244
rect 20272 38758 20300 39238
rect 20260 38752 20312 38758
rect 20260 38694 20312 38700
rect 20824 38554 20852 39374
rect 21100 39098 21128 39374
rect 21560 39098 21588 40462
rect 22284 40452 22336 40458
rect 22284 40394 22336 40400
rect 22296 40050 22324 40394
rect 22388 40050 22416 40582
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22376 40044 22428 40050
rect 22376 39986 22428 39992
rect 21088 39092 21140 39098
rect 21088 39034 21140 39040
rect 21548 39092 21600 39098
rect 21548 39034 21600 39040
rect 20996 39024 21048 39030
rect 20996 38966 21048 38972
rect 20904 38888 20956 38894
rect 20904 38830 20956 38836
rect 20812 38548 20864 38554
rect 20812 38490 20864 38496
rect 20352 38412 20404 38418
rect 20352 38354 20404 38360
rect 20260 38344 20312 38350
rect 20260 38286 20312 38292
rect 20272 37942 20300 38286
rect 20260 37936 20312 37942
rect 20260 37878 20312 37884
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20364 36378 20392 38354
rect 20628 38344 20680 38350
rect 20628 38286 20680 38292
rect 20640 38214 20668 38286
rect 20628 38208 20680 38214
rect 20628 38150 20680 38156
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20352 36372 20404 36378
rect 20352 36314 20404 36320
rect 20076 35828 20128 35834
rect 20076 35770 20128 35776
rect 19996 35686 20208 35714
rect 19892 35216 19944 35222
rect 19892 35158 19944 35164
rect 19904 35034 19932 35158
rect 19904 35006 20116 35034
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19444 34610 19564 34626
rect 19444 34604 19576 34610
rect 19444 34598 19524 34604
rect 19524 34546 19576 34552
rect 19536 33998 19564 34546
rect 19524 33992 19576 33998
rect 19524 33934 19576 33940
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33590 20024 33798
rect 19984 33584 20036 33590
rect 19984 33526 20036 33532
rect 20088 33402 20116 35006
rect 20180 33658 20208 35686
rect 20456 35494 20484 37402
rect 20536 37188 20588 37194
rect 20536 37130 20588 37136
rect 20548 36718 20576 37130
rect 20640 36922 20668 38150
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20628 36916 20680 36922
rect 20628 36858 20680 36864
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 20548 36378 20576 36654
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20732 35834 20760 37810
rect 20916 37126 20944 38830
rect 21008 38593 21036 38966
rect 21100 38962 21220 38978
rect 21100 38956 21232 38962
rect 21100 38950 21180 38956
rect 20994 38584 21050 38593
rect 20994 38519 21050 38528
rect 21100 37806 21128 38950
rect 21180 38898 21232 38904
rect 21180 38820 21232 38826
rect 21180 38762 21232 38768
rect 21192 38554 21220 38762
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 21364 38548 21416 38554
rect 21364 38490 21416 38496
rect 21088 37800 21140 37806
rect 21088 37742 21140 37748
rect 21272 37664 21324 37670
rect 21272 37606 21324 37612
rect 20904 37120 20956 37126
rect 20904 37062 20956 37068
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20824 36174 20852 36654
rect 21284 36174 21312 37606
rect 21376 37194 21404 38490
rect 22480 38026 22508 40666
rect 22572 40594 22600 41414
rect 22848 41138 22876 41550
rect 24032 41540 24084 41546
rect 24032 41482 24084 41488
rect 23848 41472 23900 41478
rect 23848 41414 23900 41420
rect 23860 41138 23888 41414
rect 22836 41132 22888 41138
rect 22836 41074 22888 41080
rect 23848 41132 23900 41138
rect 23848 41074 23900 41080
rect 23480 40928 23532 40934
rect 23480 40870 23532 40876
rect 23848 40928 23900 40934
rect 23848 40870 23900 40876
rect 23388 40656 23440 40662
rect 23388 40598 23440 40604
rect 22560 40588 22612 40594
rect 22560 40530 22612 40536
rect 23400 40526 23428 40598
rect 23388 40520 23440 40526
rect 23388 40462 23440 40468
rect 23400 40050 23428 40462
rect 23492 40458 23520 40870
rect 23480 40452 23532 40458
rect 23480 40394 23532 40400
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 23388 40044 23440 40050
rect 23388 39986 23440 39992
rect 22558 38040 22614 38049
rect 22480 37998 22558 38026
rect 22558 37975 22614 37984
rect 22572 37874 22600 37975
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 22376 37800 22428 37806
rect 22376 37742 22428 37748
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22192 37732 22244 37738
rect 22192 37674 22244 37680
rect 21364 37188 21416 37194
rect 21364 37130 21416 37136
rect 22008 36848 22060 36854
rect 22008 36790 22060 36796
rect 22098 36816 22154 36825
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21100 35834 21128 36110
rect 21916 36032 21968 36038
rect 22020 36009 22048 36790
rect 22098 36751 22100 36760
rect 22152 36751 22154 36760
rect 22100 36722 22152 36728
rect 22112 36310 22140 36722
rect 22100 36304 22152 36310
rect 22100 36246 22152 36252
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 21916 35974 21968 35980
rect 22006 36000 22062 36009
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 20444 35488 20496 35494
rect 20444 35430 20496 35436
rect 20456 35290 20484 35430
rect 20444 35284 20496 35290
rect 20444 35226 20496 35232
rect 20352 34060 20404 34066
rect 20352 34002 20404 34008
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19904 33374 20116 33402
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19904 32910 19932 33374
rect 20076 33312 20128 33318
rect 20076 33254 20128 33260
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 19996 32910 20024 33050
rect 19892 32904 19944 32910
rect 19892 32846 19944 32852
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19340 32836 19392 32842
rect 19392 32796 19472 32824
rect 19340 32778 19392 32784
rect 19444 32502 19472 32796
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19260 30326 19288 32370
rect 19996 32230 20024 32710
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31482 20024 32166
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19352 30274 19380 31078
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 30394 19472 30670
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19352 30258 19748 30274
rect 19352 30252 19760 30258
rect 19352 30246 19708 30252
rect 19708 30194 19760 30200
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19248 30116 19300 30122
rect 19248 30058 19300 30064
rect 19260 29850 19288 30058
rect 19248 29844 19300 29850
rect 19248 29786 19300 29792
rect 19720 29628 19748 30194
rect 19812 30054 19840 30194
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19892 30048 19944 30054
rect 19892 29990 19944 29996
rect 19904 29646 19932 29990
rect 19800 29640 19852 29646
rect 19720 29600 19800 29628
rect 19800 29582 19852 29588
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19352 29306 19380 29514
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 19352 29050 19380 29242
rect 19444 29170 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19996 29170 20024 30806
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19064 29028 19116 29034
rect 19064 28970 19116 28976
rect 19076 28082 19104 28970
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18602 26344 18658 26353
rect 18708 26314 18736 27270
rect 18800 26382 18828 27406
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18602 26279 18658 26288
rect 18696 26308 18748 26314
rect 18616 25498 18644 26279
rect 18696 26250 18748 26256
rect 18604 25492 18656 25498
rect 18604 25434 18656 25440
rect 18800 25226 18828 26318
rect 18984 25838 19012 26726
rect 18972 25832 19024 25838
rect 18972 25774 19024 25780
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19076 25498 19104 25774
rect 19064 25492 19116 25498
rect 19064 25434 19116 25440
rect 18788 25220 18840 25226
rect 18788 25162 18840 25168
rect 18788 23248 18840 23254
rect 18788 23190 18840 23196
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18708 22098 18736 23054
rect 18800 22642 18828 23190
rect 19168 22778 19196 29038
rect 19352 29022 19472 29050
rect 19340 26784 19392 26790
rect 19444 26772 19472 29022
rect 19524 28688 19576 28694
rect 19524 28630 19576 28636
rect 19536 28422 19564 28630
rect 20088 28490 20116 33254
rect 20272 32570 20300 33934
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20272 30734 20300 30874
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20180 26790 20208 30602
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 20272 29714 20300 30534
rect 20260 29708 20312 29714
rect 20260 29650 20312 29656
rect 20364 27470 20392 34002
rect 20628 33380 20680 33386
rect 20628 33322 20680 33328
rect 20444 32836 20496 32842
rect 20444 32778 20496 32784
rect 20456 32434 20484 32778
rect 20640 32570 20668 33322
rect 21180 32768 21232 32774
rect 21180 32710 21232 32716
rect 21192 32570 21220 32710
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 20824 30394 20852 30602
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 20824 30258 20852 30330
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20824 28490 20852 29582
rect 20916 28762 20944 31758
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 21008 30734 21036 31690
rect 20996 30728 21048 30734
rect 20996 30670 21048 30676
rect 21008 30054 21036 30670
rect 21284 30297 21312 35634
rect 21928 35630 21956 35974
rect 22006 35935 22062 35944
rect 21916 35624 21968 35630
rect 21916 35566 21968 35572
rect 22112 35578 22140 36110
rect 22204 36009 22232 37674
rect 22388 37466 22416 37742
rect 22376 37460 22428 37466
rect 22376 37402 22428 37408
rect 22480 37398 22508 37742
rect 22468 37392 22520 37398
rect 22468 37334 22520 37340
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22296 36106 22324 36722
rect 22468 36576 22520 36582
rect 22468 36518 22520 36524
rect 22480 36378 22508 36518
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22572 36258 22600 37810
rect 22756 37777 22784 37810
rect 22742 37768 22798 37777
rect 22742 37703 22798 37712
rect 22388 36230 22600 36258
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22190 36000 22246 36009
rect 22190 35935 22246 35944
rect 22204 35698 22232 35935
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22112 35562 22232 35578
rect 22112 35556 22244 35562
rect 22112 35550 22192 35556
rect 22192 35498 22244 35504
rect 22296 35290 22324 36042
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22100 35216 22152 35222
rect 22100 35158 22152 35164
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21376 32910 21404 33050
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 21914 32328 21970 32337
rect 21914 32263 21970 32272
rect 21928 31822 21956 32263
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 22008 31816 22060 31822
rect 22112 31804 22140 35158
rect 22388 33946 22416 36230
rect 22468 36168 22520 36174
rect 22520 36128 22600 36156
rect 22468 36110 22520 36116
rect 22572 35698 22600 36128
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22480 35086 22508 35566
rect 22572 35494 22600 35634
rect 22560 35488 22612 35494
rect 22560 35430 22612 35436
rect 22572 35222 22600 35430
rect 22560 35216 22612 35222
rect 22560 35158 22612 35164
rect 22468 35080 22520 35086
rect 22848 35034 22876 39986
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 23112 39432 23164 39438
rect 23112 39374 23164 39380
rect 22940 38350 22968 39374
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 23032 38418 23060 39238
rect 23124 39001 23152 39374
rect 23110 38992 23166 39001
rect 23110 38927 23166 38936
rect 23400 38894 23428 39986
rect 23492 38962 23520 40394
rect 23860 40390 23888 40870
rect 23848 40384 23900 40390
rect 23848 40326 23900 40332
rect 23848 40180 23900 40186
rect 23848 40122 23900 40128
rect 23756 39432 23808 39438
rect 23756 39374 23808 39380
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23204 38820 23256 38826
rect 23204 38762 23256 38768
rect 23020 38412 23072 38418
rect 23020 38354 23072 38360
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 23216 36156 23244 38762
rect 23480 38004 23532 38010
rect 23480 37946 23532 37952
rect 23492 37874 23520 37946
rect 23388 37868 23440 37874
rect 23388 37810 23440 37816
rect 23480 37868 23532 37874
rect 23480 37810 23532 37816
rect 23400 37262 23428 37810
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23400 36310 23428 37198
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23388 36304 23440 36310
rect 23388 36246 23440 36252
rect 23676 36174 23704 36518
rect 23768 36378 23796 39374
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23664 36168 23716 36174
rect 23216 36128 23428 36156
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 23308 35154 23336 35634
rect 23400 35562 23428 36128
rect 23664 36110 23716 36116
rect 23480 36100 23532 36106
rect 23480 36042 23532 36048
rect 23492 35834 23520 36042
rect 23860 35834 23888 40122
rect 23940 39976 23992 39982
rect 23940 39918 23992 39924
rect 23952 38554 23980 39918
rect 24044 39642 24072 41482
rect 24400 41268 24452 41274
rect 24400 41210 24452 41216
rect 24124 41132 24176 41138
rect 24124 41074 24176 41080
rect 24136 40769 24164 41074
rect 24122 40760 24178 40769
rect 24122 40695 24178 40704
rect 24124 40384 24176 40390
rect 24124 40326 24176 40332
rect 24216 40384 24268 40390
rect 24216 40326 24268 40332
rect 24136 40186 24164 40326
rect 24124 40180 24176 40186
rect 24124 40122 24176 40128
rect 24032 39636 24084 39642
rect 24032 39578 24084 39584
rect 23940 38548 23992 38554
rect 23940 38490 23992 38496
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23848 35828 23900 35834
rect 23848 35770 23900 35776
rect 23388 35556 23440 35562
rect 23388 35498 23440 35504
rect 23400 35154 23428 35498
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 22468 35022 22520 35028
rect 22480 34610 22508 35022
rect 22572 35006 22876 35034
rect 23020 35080 23072 35086
rect 23020 35022 23072 35028
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22204 33918 22416 33946
rect 22204 32434 22232 33918
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22296 33522 22324 33798
rect 22284 33516 22336 33522
rect 22284 33458 22336 33464
rect 22480 33454 22508 33798
rect 22468 33448 22520 33454
rect 22468 33390 22520 33396
rect 22376 33380 22428 33386
rect 22376 33322 22428 33328
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22060 31776 22140 31804
rect 22008 31758 22060 31764
rect 21270 30288 21326 30297
rect 21270 30223 21272 30232
rect 21324 30223 21326 30232
rect 21456 30252 21508 30258
rect 21272 30194 21324 30200
rect 21456 30194 21508 30200
rect 21468 30054 21496 30194
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 19616 26784 19668 26790
rect 19444 26744 19616 26772
rect 19340 26726 19392 26732
rect 19616 26726 19668 26732
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 19352 26450 19380 26726
rect 20088 26602 20116 26726
rect 20088 26574 20208 26602
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19444 26314 19564 26330
rect 19444 26308 19576 26314
rect 19444 26302 19524 26308
rect 19444 26042 19472 26302
rect 19524 26250 19576 26256
rect 20076 26240 20128 26246
rect 20076 26182 20128 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 20088 25974 20116 26182
rect 20076 25968 20128 25974
rect 20076 25910 20128 25916
rect 20180 25906 20208 26574
rect 20456 26246 20484 28426
rect 20824 27946 20852 28426
rect 20916 28218 20944 28426
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 20812 27940 20864 27946
rect 20812 27882 20864 27888
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27470 20760 27814
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20810 27432 20866 27441
rect 20640 26382 20668 27406
rect 20810 27367 20866 27376
rect 20824 27334 20852 27367
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20812 26988 20864 26994
rect 20916 26976 20944 28154
rect 20864 26948 20944 26976
rect 21008 26976 21036 29990
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21100 28082 21128 28358
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21100 27334 21128 28018
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 21192 26994 21220 27338
rect 21270 27160 21326 27169
rect 21376 27130 21404 27950
rect 21270 27095 21272 27104
rect 21324 27095 21326 27104
rect 21364 27124 21416 27130
rect 21272 27066 21324 27072
rect 21364 27066 21416 27072
rect 21088 26988 21140 26994
rect 21008 26948 21088 26976
rect 20812 26930 20864 26936
rect 21088 26930 21140 26936
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21272 26988 21324 26994
rect 21324 26948 21404 26976
rect 21272 26930 21324 26936
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 19996 25498 20024 25842
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 20088 25430 20116 25774
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 20364 25294 20392 25638
rect 20640 25362 20668 26318
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 21100 24818 21128 26930
rect 21376 26897 21404 26948
rect 21362 26888 21418 26897
rect 21180 26852 21232 26858
rect 21232 26812 21312 26840
rect 21362 26823 21418 26832
rect 21456 26852 21508 26858
rect 21180 26794 21232 26800
rect 21284 26738 21312 26812
rect 21456 26794 21508 26800
rect 21468 26738 21496 26794
rect 21284 26710 21496 26738
rect 21560 26382 21588 28494
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 21652 27169 21680 27474
rect 21638 27160 21694 27169
rect 21638 27095 21694 27104
rect 21652 26994 21680 27095
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18472 21304 18552 21332
rect 18420 21286 18472 21292
rect 18432 21146 18460 21286
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18156 18630 18184 18702
rect 18248 18698 18276 19314
rect 18432 19174 18460 19790
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18766 18460 19110
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18248 18358 18276 18634
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18432 18290 18460 18702
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16114 18460 16594
rect 18524 16114 18552 20266
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18616 18630 18644 19314
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18708 18426 18736 21898
rect 18892 20466 18920 22714
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 19260 19310 19288 22986
rect 19352 21162 19380 24550
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 19984 24268 20036 24274
rect 20168 24268 20220 24274
rect 20036 24228 20168 24256
rect 19984 24210 20036 24216
rect 20168 24210 20220 24216
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23730 19472 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20272 23730 20300 23802
rect 20548 23730 20576 24142
rect 21100 24070 21128 24278
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 23730 21128 24006
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 19444 22030 19472 23666
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19708 22976 19760 22982
rect 19904 22964 19932 23054
rect 19760 22936 19932 22964
rect 19984 22976 20036 22982
rect 19708 22918 19760 22924
rect 19984 22918 20036 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19904 22030 19932 22374
rect 19996 22030 20024 22918
rect 20272 22030 20300 23666
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20364 22098 20392 22918
rect 20456 22438 20484 23122
rect 20548 22778 20576 23666
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21008 23186 21036 23598
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21100 23118 21128 23666
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21192 23118 21220 23530
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21100 22964 21128 23054
rect 21180 22976 21232 22982
rect 21100 22936 21180 22964
rect 21180 22918 21232 22924
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 21192 22574 21220 22918
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20456 22166 20484 22374
rect 20548 22234 20576 22510
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20444 22160 20496 22166
rect 20444 22102 20496 22108
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19352 21134 19472 21162
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19352 20398 19380 21014
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19444 19718 19472 21134
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19514 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18766 19748 19110
rect 19996 18850 20024 21830
rect 20180 21418 20208 21830
rect 20364 21622 20392 22034
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 20466 20116 21286
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20534 20208 20810
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20088 19854 20116 20402
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20180 19718 20208 20470
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20364 19922 20392 20402
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 19996 18822 20116 18850
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 19352 17746 19380 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18702
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19444 17678 19472 18022
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19984 17672 20036 17678
rect 20088 17660 20116 18822
rect 20036 17632 20116 17660
rect 19984 17614 20036 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 16658 18644 17478
rect 19444 17202 19472 17614
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 17270 20024 17614
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15502 18552 16050
rect 18616 15502 18644 16594
rect 18800 16590 18828 16934
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 15502 18828 16526
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 19444 14958 19472 15302
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15026 20024 16050
rect 20272 15502 20300 19450
rect 20456 18714 20484 22102
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20640 20806 20668 21966
rect 21192 21486 21220 22510
rect 21284 21962 21312 25978
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 23730 21588 25434
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 22020 23798 22048 24278
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 22020 22506 22048 23734
rect 22204 23594 22232 25366
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22204 22710 22232 22918
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22008 22500 22060 22506
rect 22008 22442 22060 22448
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20640 19786 20668 20742
rect 20916 20466 20944 21014
rect 21284 20942 21312 21898
rect 21376 21554 21404 21898
rect 21468 21554 21496 21966
rect 22112 21554 22140 22102
rect 22204 22030 22232 22442
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21468 21010 21496 21490
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 22204 20942 22232 21966
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20916 19922 20944 20402
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20640 18834 20668 19722
rect 21284 19310 21312 20878
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20364 18686 20484 18714
rect 20364 18222 20392 18686
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20456 17678 20484 18566
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20456 17202 20484 17614
rect 20916 17202 20944 19110
rect 21284 18834 21312 19246
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 17270 21036 18566
rect 21284 18426 21312 18770
rect 21376 18630 21404 20742
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21376 18358 21404 18566
rect 21364 18352 21416 18358
rect 21364 18294 21416 18300
rect 22112 17746 22140 20402
rect 22296 18154 22324 33254
rect 22388 30802 22416 33322
rect 22480 32842 22508 33390
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22388 29578 22416 30738
rect 22376 29572 22428 29578
rect 22376 29514 22428 29520
rect 22388 24818 22416 29514
rect 22572 28966 22600 35006
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22652 32972 22704 32978
rect 22652 32914 22704 32920
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22572 25906 22600 27610
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 24206 22416 24550
rect 22480 24410 22508 24754
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23798 22508 24006
rect 22468 23792 22520 23798
rect 22388 23752 22468 23780
rect 22388 23050 22416 23752
rect 22468 23734 22520 23740
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22480 23225 22508 23258
rect 22466 23216 22522 23225
rect 22466 23151 22522 23160
rect 22480 23118 22508 23151
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22376 23044 22428 23050
rect 22376 22986 22428 22992
rect 22572 22778 22600 23054
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22572 22030 22600 22714
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22664 21706 22692 32914
rect 22756 32026 22784 34682
rect 23032 34134 23060 35022
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23124 34474 23152 34954
rect 23112 34468 23164 34474
rect 23112 34410 23164 34416
rect 23020 34128 23072 34134
rect 23020 34070 23072 34076
rect 23032 33998 23060 34070
rect 23124 34066 23152 34410
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22928 33924 22980 33930
rect 22928 33866 22980 33872
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22848 32570 22876 32846
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22940 32434 22968 33866
rect 23216 33114 23244 34954
rect 23204 33108 23256 33114
rect 23204 33050 23256 33056
rect 23216 32434 23244 33050
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23020 32360 23072 32366
rect 23020 32302 23072 32308
rect 22744 32020 22796 32026
rect 22744 31962 22796 31968
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22940 31346 22968 31622
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22848 28762 22876 29786
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 22940 29238 22968 29650
rect 22928 29232 22980 29238
rect 22928 29174 22980 29180
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 23032 28558 23060 32302
rect 23112 32224 23164 32230
rect 23112 32166 23164 32172
rect 23124 31822 23152 32166
rect 23308 31822 23336 35090
rect 23400 34610 23428 35090
rect 23952 35086 23980 38490
rect 24032 35692 24084 35698
rect 24032 35634 24084 35640
rect 23940 35080 23992 35086
rect 23940 35022 23992 35028
rect 23952 34610 23980 35022
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 23848 33924 23900 33930
rect 23848 33866 23900 33872
rect 23860 33590 23888 33866
rect 23848 33584 23900 33590
rect 23848 33526 23900 33532
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 23676 33046 23704 33390
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23676 32910 23704 32982
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23388 32768 23440 32774
rect 23388 32710 23440 32716
rect 23400 32434 23428 32710
rect 23860 32434 23888 33526
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23848 32428 23900 32434
rect 23848 32370 23900 32376
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23400 31890 23428 31962
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 23492 31822 23520 32166
rect 23112 31816 23164 31822
rect 23296 31816 23348 31822
rect 23112 31758 23164 31764
rect 23294 31784 23296 31793
rect 23480 31816 23532 31822
rect 23348 31784 23350 31793
rect 23124 31414 23152 31758
rect 23480 31758 23532 31764
rect 23676 31754 23704 32370
rect 23756 32224 23808 32230
rect 23756 32166 23808 32172
rect 23294 31719 23350 31728
rect 23584 31726 23704 31754
rect 23112 31408 23164 31414
rect 23112 31350 23164 31356
rect 23584 31142 23612 31726
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23584 30938 23612 31078
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23676 30802 23704 31078
rect 23664 30796 23716 30802
rect 23664 30738 23716 30744
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23216 29714 23244 30534
rect 23584 30394 23612 30534
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23584 29850 23612 30126
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23204 29708 23256 29714
rect 23204 29650 23256 29656
rect 23202 29608 23258 29617
rect 23202 29543 23258 29552
rect 23216 29510 23244 29543
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 23020 28552 23072 28558
rect 22940 28512 23020 28540
rect 22940 28150 22968 28512
rect 23020 28494 23072 28500
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23112 28484 23164 28490
rect 23112 28426 23164 28432
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 23032 27470 23060 28358
rect 23020 27464 23072 27470
rect 22940 27412 23020 27418
rect 22940 27406 23072 27412
rect 22940 27390 23060 27406
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26858 22784 27270
rect 22940 26994 22968 27390
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22744 26852 22796 26858
rect 22744 26794 22796 26800
rect 23032 26450 23060 27270
rect 23124 27130 23152 28426
rect 23216 27674 23244 28494
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23296 28008 23348 28014
rect 23296 27950 23348 27956
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23216 26926 23244 27270
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23020 26444 23072 26450
rect 23020 26386 23072 26392
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 22928 26240 22980 26246
rect 22928 26182 22980 26188
rect 22940 25974 22968 26182
rect 23216 25974 23244 26318
rect 22928 25968 22980 25974
rect 22928 25910 22980 25916
rect 23204 25968 23256 25974
rect 23204 25910 23256 25916
rect 23308 25226 23336 27950
rect 23584 27606 23612 28018
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23768 26994 23796 32166
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23860 30802 23888 31282
rect 23848 30796 23900 30802
rect 23848 30738 23900 30744
rect 24044 30122 24072 35634
rect 24136 32978 24164 40122
rect 24228 40050 24256 40326
rect 24216 40044 24268 40050
rect 24216 39986 24268 39992
rect 24228 38758 24256 39986
rect 24216 38752 24268 38758
rect 24216 38694 24268 38700
rect 24228 35698 24256 38694
rect 24308 38344 24360 38350
rect 24308 38286 24360 38292
rect 24216 35692 24268 35698
rect 24216 35634 24268 35640
rect 24216 35488 24268 35494
rect 24320 35476 24348 38286
rect 24268 35448 24348 35476
rect 24216 35430 24268 35436
rect 24320 34610 24348 35448
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24320 33522 24348 34546
rect 24308 33516 24360 33522
rect 24308 33458 24360 33464
rect 24124 32972 24176 32978
rect 24124 32914 24176 32920
rect 24320 32910 24348 33458
rect 24308 32904 24360 32910
rect 24308 32846 24360 32852
rect 24124 31136 24176 31142
rect 24124 31078 24176 31084
rect 24136 30870 24164 31078
rect 24124 30864 24176 30870
rect 24124 30806 24176 30812
rect 24308 30252 24360 30258
rect 24308 30194 24360 30200
rect 24032 30116 24084 30122
rect 24032 30058 24084 30064
rect 24320 30054 24348 30194
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24320 29850 24348 29990
rect 24308 29844 24360 29850
rect 24308 29786 24360 29792
rect 24124 28484 24176 28490
rect 24124 28426 24176 28432
rect 24136 28218 24164 28426
rect 24124 28212 24176 28218
rect 24124 28154 24176 28160
rect 24032 28008 24084 28014
rect 24032 27950 24084 27956
rect 24044 27062 24072 27950
rect 24136 27878 24164 28154
rect 24124 27872 24176 27878
rect 24124 27814 24176 27820
rect 24032 27056 24084 27062
rect 24032 26998 24084 27004
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 23756 26988 23808 26994
rect 23756 26930 23808 26936
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23400 26382 23428 26726
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 25220 23348 25226
rect 23296 25162 23348 25168
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22756 24206 22784 24686
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22848 24410 22876 24618
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22756 23526 22784 24142
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 22480 21678 22692 21706
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22112 17610 22140 17682
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22020 17270 22048 17478
rect 22204 17270 22232 17478
rect 22480 17338 22508 21678
rect 23032 21554 23060 21898
rect 23216 21690 23244 23122
rect 23308 21894 23336 25162
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23492 24206 23520 24686
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23492 22778 23520 23666
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22664 20466 22692 21490
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22756 20534 22784 21286
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22664 19990 22692 20402
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20548 16114 20576 17070
rect 20916 16522 20944 17138
rect 21008 16590 21036 17206
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20824 16114 20852 16458
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20916 15638 20944 15846
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 20916 15502 20944 15574
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 18432 14618 18460 14894
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18892 14482 18920 14758
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 19444 14414 19472 14894
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19444 13870 19472 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 13938 20024 14962
rect 20364 14890 20392 15438
rect 21100 15026 21128 15846
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20180 14074 20208 14758
rect 20364 14550 20392 14826
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20732 14414 20760 14962
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20732 13938 20760 14350
rect 21284 14346 21312 15438
rect 22020 14482 22048 17002
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22112 16726 22140 16934
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 22204 16590 22232 16934
rect 22296 16590 22324 17206
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22480 16590 22508 17138
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22284 16584 22336 16590
rect 22468 16584 22520 16590
rect 22284 16526 22336 16532
rect 22388 16544 22468 16572
rect 22204 16182 22232 16526
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22296 15910 22324 16526
rect 22388 16182 22416 16544
rect 22468 16526 22520 16532
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22112 15026 22140 15370
rect 22296 15162 22324 15846
rect 22388 15706 22416 16118
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22572 15502 22600 19654
rect 22848 18766 22876 20742
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19854 23060 20198
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22940 19514 22968 19790
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22664 18290 22692 18702
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22756 17882 22784 18566
rect 22940 18426 22968 18566
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 23032 18358 23060 19450
rect 23124 19378 23152 19654
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23020 18352 23072 18358
rect 23020 18294 23072 18300
rect 23112 18148 23164 18154
rect 23112 18090 23164 18096
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 16454 22692 17682
rect 22756 17678 22784 17818
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 16182 22692 16390
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 15502 22784 15846
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22572 15026 22600 15438
rect 23124 15026 23152 18090
rect 23216 17678 23244 21422
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23308 19378 23336 20742
rect 23400 20330 23428 20878
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23400 18902 23428 19722
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23308 15094 23336 17274
rect 23400 16182 23428 18022
rect 23584 17338 23612 26930
rect 24216 26920 24268 26926
rect 24216 26862 24268 26868
rect 24412 26874 24440 41210
rect 24676 41064 24728 41070
rect 24676 41006 24728 41012
rect 24688 40050 24716 41006
rect 24964 40934 24992 42094
rect 27264 41818 27292 42162
rect 27528 42016 27580 42022
rect 27528 41958 27580 41964
rect 27252 41812 27304 41818
rect 27252 41754 27304 41760
rect 26976 41540 27028 41546
rect 26976 41482 27028 41488
rect 26238 41304 26294 41313
rect 26238 41239 26294 41248
rect 25228 41132 25280 41138
rect 25228 41074 25280 41080
rect 25964 41132 26016 41138
rect 25964 41074 26016 41080
rect 24952 40928 25004 40934
rect 24952 40870 25004 40876
rect 24860 40656 24912 40662
rect 24860 40598 24912 40604
rect 24872 40526 24900 40598
rect 24860 40520 24912 40526
rect 24860 40462 24912 40468
rect 24768 40452 24820 40458
rect 24768 40394 24820 40400
rect 24780 40050 24808 40394
rect 24964 40186 24992 40870
rect 25240 40730 25268 41074
rect 25228 40724 25280 40730
rect 25228 40666 25280 40672
rect 25976 40526 26004 41074
rect 26252 41070 26280 41239
rect 26240 41064 26292 41070
rect 26240 41006 26292 41012
rect 26252 40594 26280 41006
rect 26240 40588 26292 40594
rect 26240 40530 26292 40536
rect 26516 40588 26568 40594
rect 26516 40530 26568 40536
rect 25964 40520 26016 40526
rect 25964 40462 26016 40468
rect 25976 40390 26004 40462
rect 26148 40452 26200 40458
rect 26148 40394 26200 40400
rect 25964 40384 26016 40390
rect 25964 40326 26016 40332
rect 24952 40180 25004 40186
rect 24952 40122 25004 40128
rect 26160 40050 26188 40394
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 24676 40044 24728 40050
rect 24676 39986 24728 39992
rect 24768 40044 24820 40050
rect 24768 39986 24820 39992
rect 26148 40044 26200 40050
rect 26148 39986 26200 39992
rect 25044 39976 25096 39982
rect 25044 39918 25096 39924
rect 24584 39908 24636 39914
rect 24584 39850 24636 39856
rect 24492 38956 24544 38962
rect 24492 38898 24544 38904
rect 24504 37874 24532 38898
rect 24596 38758 24624 39850
rect 24952 39364 25004 39370
rect 24952 39306 25004 39312
rect 24964 38962 24992 39306
rect 24952 38956 25004 38962
rect 24952 38898 25004 38904
rect 25056 38826 25084 39918
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 25044 38820 25096 38826
rect 25044 38762 25096 38768
rect 24584 38752 24636 38758
rect 24584 38694 24636 38700
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 24492 37664 24544 37670
rect 24492 37606 24544 37612
rect 24504 36242 24532 37606
rect 24596 36922 24624 38694
rect 24860 38548 24912 38554
rect 24860 38490 24912 38496
rect 24872 38010 24900 38490
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 24768 37800 24820 37806
rect 24768 37742 24820 37748
rect 24780 37398 24808 37742
rect 24768 37392 24820 37398
rect 24768 37334 24820 37340
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 24872 36786 24900 37946
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 25056 37210 25084 38762
rect 25136 38208 25188 38214
rect 25136 38150 25188 38156
rect 25228 38208 25280 38214
rect 25228 38150 25280 38156
rect 25148 37874 25176 38150
rect 25240 37942 25268 38150
rect 25228 37936 25280 37942
rect 25228 37878 25280 37884
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25228 37664 25280 37670
rect 25228 37606 25280 37612
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24860 36644 24912 36650
rect 24860 36586 24912 36592
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 24584 35828 24636 35834
rect 24584 35770 24636 35776
rect 24596 34746 24624 35770
rect 24768 35488 24820 35494
rect 24768 35430 24820 35436
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 24780 34474 24808 35430
rect 24872 35018 24900 36586
rect 24964 36310 24992 37198
rect 25056 37182 25176 37210
rect 25240 37194 25268 37606
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 25056 36786 25084 37062
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 24952 36304 25004 36310
rect 24952 36246 25004 36252
rect 24860 35012 24912 35018
rect 24860 34954 24912 34960
rect 24860 34672 24912 34678
rect 24860 34614 24912 34620
rect 24768 34468 24820 34474
rect 24768 34410 24820 34416
rect 24780 32978 24808 34410
rect 24872 33998 24900 34614
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 33318 24900 33458
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 24780 32858 24808 32914
rect 24688 32830 24808 32858
rect 24688 31822 24716 32830
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24780 32502 24808 32710
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24872 31822 24900 33254
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24964 31686 24992 36246
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 25056 35766 25084 36110
rect 25148 36038 25176 37182
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25148 35766 25176 35974
rect 25044 35760 25096 35766
rect 25136 35760 25188 35766
rect 25044 35702 25096 35708
rect 25134 35728 25136 35737
rect 25188 35728 25190 35737
rect 25134 35663 25190 35672
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25148 35290 25176 35566
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 25044 35012 25096 35018
rect 25044 34954 25096 34960
rect 25056 34542 25084 34954
rect 25044 34536 25096 34542
rect 25044 34478 25096 34484
rect 25240 33114 25268 37130
rect 25332 34610 25360 39782
rect 26252 39273 26280 40122
rect 26238 39264 26294 39273
rect 26238 39199 26294 39208
rect 26528 39098 26556 40530
rect 26988 40526 27016 41482
rect 27264 41138 27292 41754
rect 27540 41682 27568 41958
rect 27344 41676 27396 41682
rect 27344 41618 27396 41624
rect 27528 41676 27580 41682
rect 27528 41618 27580 41624
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 27068 40928 27120 40934
rect 27068 40870 27120 40876
rect 27080 40526 27108 40870
rect 26976 40520 27028 40526
rect 26976 40462 27028 40468
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26792 40384 26844 40390
rect 26792 40326 26844 40332
rect 26608 39840 26660 39846
rect 26608 39782 26660 39788
rect 26516 39092 26568 39098
rect 26516 39034 26568 39040
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 26068 38826 26096 38898
rect 26424 38888 26476 38894
rect 26620 38842 26648 39782
rect 26476 38836 26648 38842
rect 26424 38830 26648 38836
rect 26056 38820 26108 38826
rect 26436 38814 26648 38830
rect 26056 38762 26108 38768
rect 25872 38480 25924 38486
rect 25872 38422 25924 38428
rect 25412 38004 25464 38010
rect 25412 37946 25464 37952
rect 25424 36825 25452 37946
rect 25884 37874 25912 38422
rect 25964 38344 26016 38350
rect 25964 38286 26016 38292
rect 25872 37868 25924 37874
rect 25872 37810 25924 37816
rect 25780 37800 25832 37806
rect 25780 37742 25832 37748
rect 25688 37664 25740 37670
rect 25688 37606 25740 37612
rect 25596 37392 25648 37398
rect 25596 37334 25648 37340
rect 25504 37256 25556 37262
rect 25504 37198 25556 37204
rect 25410 36816 25466 36825
rect 25410 36751 25466 36760
rect 25412 36032 25464 36038
rect 25412 35974 25464 35980
rect 25424 35562 25452 35974
rect 25412 35556 25464 35562
rect 25412 35498 25464 35504
rect 25412 34944 25464 34950
rect 25412 34886 25464 34892
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25424 34490 25452 34886
rect 25332 34462 25452 34490
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25332 32722 25360 34462
rect 25412 34400 25464 34406
rect 25412 34342 25464 34348
rect 25424 33522 25452 34342
rect 25516 34066 25544 37198
rect 25608 36582 25636 37334
rect 25700 37330 25728 37606
rect 25688 37324 25740 37330
rect 25688 37266 25740 37272
rect 25792 37262 25820 37742
rect 25884 37738 25912 37810
rect 25872 37732 25924 37738
rect 25872 37674 25924 37680
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25872 36848 25924 36854
rect 25872 36790 25924 36796
rect 25596 36576 25648 36582
rect 25596 36518 25648 36524
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25516 33590 25544 34002
rect 25504 33584 25556 33590
rect 25504 33526 25556 33532
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25332 32694 25636 32722
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 24952 31680 25004 31686
rect 24952 31622 25004 31628
rect 24860 31272 24912 31278
rect 24860 31214 24912 31220
rect 24492 31204 24544 31210
rect 24492 31146 24544 31152
rect 24504 30190 24532 31146
rect 24872 30598 24900 31214
rect 25148 30938 25176 31894
rect 25240 31822 25268 32370
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25332 31754 25360 32506
rect 25332 31726 25452 31754
rect 25320 31680 25372 31686
rect 25320 31622 25372 31628
rect 25332 31346 25360 31622
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24492 30184 24544 30190
rect 24492 30126 24544 30132
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 24596 28082 24624 28562
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24596 27470 24624 28018
rect 24688 27606 24716 28086
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24872 27538 24900 30534
rect 24964 28082 24992 30874
rect 25240 30870 25268 31078
rect 25424 30938 25452 31726
rect 25412 30932 25464 30938
rect 25412 30874 25464 30880
rect 25228 30864 25280 30870
rect 25228 30806 25280 30812
rect 25044 30796 25096 30802
rect 25044 30738 25096 30744
rect 25056 30258 25084 30738
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25332 29646 25360 30194
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25424 29102 25452 30670
rect 25608 30258 25636 32694
rect 25700 31754 25728 35634
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25792 34678 25820 35022
rect 25884 35018 25912 36790
rect 25976 36582 26004 38286
rect 26068 37466 26096 38762
rect 26148 38752 26200 38758
rect 26148 38694 26200 38700
rect 26160 37670 26188 38694
rect 26700 37868 26752 37874
rect 26700 37810 26752 37816
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 26148 37664 26200 37670
rect 26148 37606 26200 37612
rect 26056 37460 26108 37466
rect 26056 37402 26108 37408
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 26160 35494 26188 37606
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 26252 35170 26280 37742
rect 26516 37324 26568 37330
rect 26516 37266 26568 37272
rect 26528 36174 26556 37266
rect 26712 37126 26740 37810
rect 26700 37120 26752 37126
rect 26700 37062 26752 37068
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26160 35142 26280 35170
rect 26160 35086 26188 35142
rect 26148 35080 26200 35086
rect 26148 35022 26200 35028
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25780 34672 25832 34678
rect 25780 34614 25832 34620
rect 25792 32502 25820 34614
rect 25872 34536 25924 34542
rect 26252 34490 26280 35022
rect 26344 34610 26372 35566
rect 26332 34604 26384 34610
rect 26332 34546 26384 34552
rect 25872 34478 25924 34484
rect 25884 34134 25912 34478
rect 26068 34462 26280 34490
rect 25872 34128 25924 34134
rect 25872 34070 25924 34076
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 25884 31822 25912 34070
rect 25962 33960 26018 33969
rect 26068 33930 26096 34462
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 25962 33895 25964 33904
rect 26016 33895 26018 33904
rect 26056 33924 26108 33930
rect 25964 33866 26016 33872
rect 26056 33866 26108 33872
rect 25964 33652 26016 33658
rect 25964 33594 26016 33600
rect 25976 32570 26004 33594
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 26068 32434 26096 33866
rect 26148 32836 26200 32842
rect 26148 32778 26200 32784
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26068 31822 26096 32370
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26160 31804 26188 32778
rect 26252 31958 26280 33934
rect 26240 31952 26292 31958
rect 26240 31894 26292 31900
rect 26240 31816 26292 31822
rect 26160 31776 26240 31804
rect 25688 31748 25740 31754
rect 25688 31690 25740 31696
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25700 29782 25728 31690
rect 26068 30954 26096 31758
rect 25884 30926 26096 30954
rect 25884 30734 25912 30926
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25780 30388 25832 30394
rect 25780 30330 25832 30336
rect 25688 29776 25740 29782
rect 25688 29718 25740 29724
rect 25412 29096 25464 29102
rect 25412 29038 25464 29044
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24872 26994 24900 27474
rect 25056 27470 25084 27950
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 25240 26926 25268 27270
rect 25228 26920 25280 26926
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 23952 25702 23980 25910
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23768 24274 23796 24754
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23860 22642 23888 24550
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23860 22234 23888 22578
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23768 18766 23796 19858
rect 23952 19854 23980 20402
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23952 19514 23980 19790
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23860 19394 23888 19450
rect 24044 19394 24072 20266
rect 23860 19378 24072 19394
rect 23860 19372 24084 19378
rect 23860 19366 24032 19372
rect 24032 19314 24084 19320
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 24136 17814 24164 23530
rect 24228 22094 24256 26862
rect 24412 26846 24716 26874
rect 25424 26897 25452 28018
rect 25792 27674 25820 30330
rect 25884 30326 25912 30670
rect 25872 30320 25924 30326
rect 25872 30262 25924 30268
rect 26056 30116 26108 30122
rect 26056 30058 26108 30064
rect 26068 29034 26096 30058
rect 26160 29306 26188 31776
rect 26344 31793 26372 34546
rect 26422 33688 26478 33697
rect 26422 33623 26424 33632
rect 26476 33623 26478 33632
rect 26424 33594 26476 33600
rect 26528 32722 26556 36110
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26620 33522 26648 35430
rect 26608 33516 26660 33522
rect 26608 33458 26660 33464
rect 26712 32978 26740 37062
rect 26804 34202 26832 40326
rect 26988 38962 27016 40462
rect 27080 40186 27108 40462
rect 27160 40452 27212 40458
rect 27160 40394 27212 40400
rect 27252 40452 27304 40458
rect 27252 40394 27304 40400
rect 27068 40180 27120 40186
rect 27068 40122 27120 40128
rect 27172 40050 27200 40394
rect 27264 40118 27292 40394
rect 27252 40112 27304 40118
rect 27252 40054 27304 40060
rect 27160 40044 27212 40050
rect 27160 39986 27212 39992
rect 27068 39976 27120 39982
rect 27068 39918 27120 39924
rect 26976 38956 27028 38962
rect 26976 38898 27028 38904
rect 27080 38654 27108 39918
rect 27252 39908 27304 39914
rect 27252 39850 27304 39856
rect 27160 39500 27212 39506
rect 27160 39442 27212 39448
rect 27172 39098 27200 39442
rect 27264 39273 27292 39850
rect 27356 39506 27384 41618
rect 27896 41472 27948 41478
rect 27896 41414 27948 41420
rect 27620 40724 27672 40730
rect 27620 40666 27672 40672
rect 27632 40225 27660 40666
rect 27908 40526 27936 41414
rect 28080 41064 28132 41070
rect 28080 41006 28132 41012
rect 28092 40526 28120 41006
rect 27896 40520 27948 40526
rect 27896 40462 27948 40468
rect 28080 40520 28132 40526
rect 28080 40462 28132 40468
rect 27618 40216 27674 40225
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 27540 40174 27618 40202
rect 27344 39500 27396 39506
rect 27344 39442 27396 39448
rect 27250 39264 27306 39273
rect 27250 39199 27306 39208
rect 27160 39092 27212 39098
rect 27160 39034 27212 39040
rect 26988 38626 27108 38654
rect 26988 37262 27016 38626
rect 27068 38344 27120 38350
rect 27068 38286 27120 38292
rect 27160 38344 27212 38350
rect 27160 38286 27212 38292
rect 27080 37874 27108 38286
rect 27068 37868 27120 37874
rect 27068 37810 27120 37816
rect 27172 37262 27200 38286
rect 27448 37346 27476 40122
rect 27540 38282 27568 40174
rect 27618 40151 27674 40160
rect 27620 40044 27672 40050
rect 27620 39986 27672 39992
rect 27632 39642 27660 39986
rect 27620 39636 27672 39642
rect 27620 39578 27672 39584
rect 27632 38944 27660 39578
rect 27908 39438 27936 40462
rect 28092 40186 28120 40462
rect 28080 40180 28132 40186
rect 28080 40122 28132 40128
rect 28368 40089 28396 42230
rect 30564 42220 30616 42226
rect 30564 42162 30616 42168
rect 34152 42220 34204 42226
rect 34152 42162 34204 42168
rect 30012 42084 30064 42090
rect 30012 42026 30064 42032
rect 28540 41608 28592 41614
rect 28540 41550 28592 41556
rect 28908 41608 28960 41614
rect 28908 41550 28960 41556
rect 28446 41168 28502 41177
rect 28446 41103 28502 41112
rect 28460 41070 28488 41103
rect 28448 41064 28500 41070
rect 28448 41006 28500 41012
rect 28552 41002 28580 41550
rect 28920 41414 28948 41550
rect 29920 41540 29972 41546
rect 29920 41482 29972 41488
rect 28920 41386 29132 41414
rect 28906 41304 28962 41313
rect 28632 41268 28684 41274
rect 28816 41268 28868 41274
rect 28632 41210 28684 41216
rect 28736 41228 28816 41256
rect 28644 41041 28672 41210
rect 28736 41177 28764 41228
rect 29104 41274 29132 41386
rect 28906 41239 28962 41248
rect 29000 41268 29052 41274
rect 28816 41210 28868 41216
rect 28920 41206 28948 41239
rect 29000 41210 29052 41216
rect 29092 41268 29144 41274
rect 29092 41210 29144 41216
rect 28908 41200 28960 41206
rect 28722 41168 28778 41177
rect 28908 41142 28960 41148
rect 28722 41103 28778 41112
rect 28816 41064 28868 41070
rect 28630 41032 28686 41041
rect 28540 40996 28592 41002
rect 28814 41032 28816 41041
rect 28868 41032 28870 41041
rect 28630 40967 28686 40976
rect 28724 40996 28776 41002
rect 28540 40938 28592 40944
rect 28448 40928 28500 40934
rect 28448 40870 28500 40876
rect 28460 40769 28488 40870
rect 28446 40760 28502 40769
rect 28446 40695 28502 40704
rect 28540 40384 28592 40390
rect 28540 40326 28592 40332
rect 28354 40080 28410 40089
rect 28354 40015 28410 40024
rect 28172 39976 28224 39982
rect 28172 39918 28224 39924
rect 27896 39432 27948 39438
rect 27896 39374 27948 39380
rect 27804 38956 27856 38962
rect 27632 38916 27804 38944
rect 27528 38276 27580 38282
rect 27528 38218 27580 38224
rect 27528 37868 27580 37874
rect 27528 37810 27580 37816
rect 27264 37318 27476 37346
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 26882 36272 26938 36281
rect 26882 36207 26884 36216
rect 26936 36207 26938 36216
rect 26884 36178 26936 36184
rect 26792 34196 26844 34202
rect 26792 34138 26844 34144
rect 26804 33590 26832 34138
rect 26896 33998 26924 36178
rect 26988 34474 27016 37198
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 27172 36242 27200 36654
rect 27160 36236 27212 36242
rect 27160 36178 27212 36184
rect 27068 35692 27120 35698
rect 27068 35634 27120 35640
rect 27080 35290 27108 35634
rect 27264 35578 27292 37318
rect 27436 37188 27488 37194
rect 27436 37130 27488 37136
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27172 35550 27292 35578
rect 27068 35284 27120 35290
rect 27068 35226 27120 35232
rect 27068 35148 27120 35154
rect 27172 35136 27200 35550
rect 27120 35108 27200 35136
rect 27068 35090 27120 35096
rect 27068 35012 27120 35018
rect 27068 34954 27120 34960
rect 26976 34468 27028 34474
rect 26976 34410 27028 34416
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26884 33856 26936 33862
rect 26884 33798 26936 33804
rect 26896 33590 26924 33798
rect 26792 33584 26844 33590
rect 26792 33526 26844 33532
rect 26884 33584 26936 33590
rect 26884 33526 26936 33532
rect 26976 33040 27028 33046
rect 26976 32982 27028 32988
rect 26700 32972 26752 32978
rect 26700 32914 26752 32920
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 26528 32694 26740 32722
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 26240 31758 26292 31764
rect 26330 31784 26386 31793
rect 26330 31719 26386 31728
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26252 30734 26280 31622
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26344 30258 26372 31719
rect 26528 31278 26556 32370
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 26436 31142 26464 31214
rect 26424 31136 26476 31142
rect 26424 31078 26476 31084
rect 26436 30802 26464 31078
rect 26424 30796 26476 30802
rect 26424 30738 26476 30744
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26528 29578 26556 31214
rect 26712 30870 26740 32694
rect 26792 32292 26844 32298
rect 26792 32234 26844 32240
rect 26700 30864 26752 30870
rect 26700 30806 26752 30812
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26056 29028 26108 29034
rect 26056 28970 26108 28976
rect 26436 28422 26464 29106
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 25686 27432 25742 27441
rect 25686 27367 25688 27376
rect 25740 27367 25742 27376
rect 25688 27338 25740 27344
rect 25976 26994 26004 27610
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25228 26862 25280 26868
rect 25410 26888 25466 26897
rect 24688 26790 24716 26846
rect 25410 26823 25466 26832
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24504 24177 24532 25434
rect 24584 24200 24636 24206
rect 24490 24168 24546 24177
rect 24584 24142 24636 24148
rect 24490 24103 24492 24112
rect 24544 24103 24546 24112
rect 24492 24074 24544 24080
rect 24596 23866 24624 24142
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24584 23860 24636 23866
rect 24584 23802 24636 23808
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 23322 24348 23666
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24412 22778 24440 23802
rect 24688 23798 24716 24006
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 24780 23322 24808 25638
rect 24964 24886 24992 25842
rect 24952 24880 25004 24886
rect 24952 24822 25004 24828
rect 25424 24818 25452 26823
rect 26252 26790 26280 27066
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 25596 26512 25648 26518
rect 25596 26454 25648 26460
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24228 22066 24348 22094
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24228 19854 24256 20470
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23584 16794 23612 17138
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23952 16794 23980 17070
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23584 16250 23612 16526
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23400 15502 23428 16118
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 22020 12850 22048 14418
rect 23124 13190 23152 14962
rect 23400 14890 23428 15438
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23676 14278 23704 15030
rect 23860 14414 23888 15982
rect 24136 15638 24164 15982
rect 24124 15632 24176 15638
rect 24124 15574 24176 15580
rect 24320 15434 24348 22066
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24688 21690 24716 21830
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24780 21298 24808 23054
rect 24872 22982 24900 24686
rect 25320 24336 25372 24342
rect 25320 24278 25372 24284
rect 25332 23594 25360 24278
rect 25424 23594 25452 24754
rect 25608 23798 25636 26454
rect 26436 25906 26464 28358
rect 26528 27470 26556 29514
rect 26700 29096 26752 29102
rect 26700 29038 26752 29044
rect 26608 27600 26660 27606
rect 26608 27542 26660 27548
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26528 25906 26556 27270
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25700 24954 25728 25230
rect 25884 24954 25912 25230
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25320 23588 25372 23594
rect 25320 23530 25372 23536
rect 25412 23588 25464 23594
rect 25412 23530 25464 23536
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25056 23186 25084 23462
rect 25148 23186 25176 23462
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 25332 22710 25360 23530
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25332 22522 25360 22646
rect 24952 22432 25004 22438
rect 25240 22420 25268 22510
rect 25332 22494 25452 22522
rect 25240 22392 25360 22420
rect 24952 22374 25004 22380
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24872 21554 24900 21966
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24964 21486 24992 22374
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24860 21344 24912 21350
rect 24688 21292 24860 21298
rect 24688 21286 24912 21292
rect 24688 21270 24900 21286
rect 24688 19990 24716 21270
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24780 20806 24808 21082
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24872 20466 24900 20878
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24964 20346 24992 21082
rect 24872 20318 24992 20346
rect 24872 20058 24900 20318
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24676 19984 24728 19990
rect 24676 19926 24728 19932
rect 24768 19984 24820 19990
rect 24768 19926 24820 19932
rect 24780 19378 24808 19926
rect 24964 19854 24992 20198
rect 25056 19922 25084 21422
rect 25148 21146 25176 21966
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25240 20942 25268 22170
rect 25332 20942 25360 22392
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24872 19242 24900 19790
rect 25056 19378 25084 19858
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 25240 18970 25268 19722
rect 25332 19378 25360 20334
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25424 18902 25452 22494
rect 25516 19854 25544 22918
rect 25608 22574 25636 23734
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 22438 25636 22510
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25792 22234 25820 22986
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25884 22094 25912 24890
rect 26620 23254 26648 27542
rect 26712 23798 26740 29038
rect 26804 28558 26832 32234
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26896 28150 26924 32846
rect 26988 32774 27016 32982
rect 26976 32768 27028 32774
rect 26976 32710 27028 32716
rect 26988 31822 27016 32710
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26988 31346 27016 31758
rect 27080 31754 27108 34954
rect 27172 34678 27200 35108
rect 27160 34672 27212 34678
rect 27160 34614 27212 34620
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 27172 33318 27200 33934
rect 27252 33516 27304 33522
rect 27252 33458 27304 33464
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 31890 27200 33254
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 27068 31748 27120 31754
rect 27068 31690 27120 31696
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 27068 31136 27120 31142
rect 27068 31078 27120 31084
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 26988 29646 27016 30670
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 27080 29594 27108 31078
rect 27264 29714 27292 33458
rect 27356 32570 27384 36722
rect 27448 36038 27476 37130
rect 27540 36854 27568 37810
rect 27632 37466 27660 38916
rect 27804 38898 27856 38904
rect 27712 38820 27764 38826
rect 27712 38762 27764 38768
rect 27724 37670 27752 38762
rect 27712 37664 27764 37670
rect 27712 37606 27764 37612
rect 27620 37460 27672 37466
rect 27620 37402 27672 37408
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27632 37194 27660 37266
rect 27908 37262 27936 39374
rect 27988 39024 28040 39030
rect 27988 38966 28040 38972
rect 27896 37256 27948 37262
rect 27896 37198 27948 37204
rect 27620 37188 27672 37194
rect 27620 37130 27672 37136
rect 27528 36848 27580 36854
rect 27528 36790 27580 36796
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27710 36680 27766 36689
rect 27540 36378 27568 36654
rect 27710 36615 27766 36624
rect 27724 36582 27752 36615
rect 28000 36582 28028 38966
rect 28080 38820 28132 38826
rect 28080 38762 28132 38768
rect 28092 37874 28120 38762
rect 28184 38350 28212 39918
rect 28552 39574 28580 40326
rect 28540 39568 28592 39574
rect 28540 39510 28592 39516
rect 28264 39364 28316 39370
rect 28264 39306 28316 39312
rect 28172 38344 28224 38350
rect 28172 38286 28224 38292
rect 28276 38214 28304 39306
rect 28540 38956 28592 38962
rect 28540 38898 28592 38904
rect 28354 38448 28410 38457
rect 28552 38418 28580 38898
rect 28354 38383 28410 38392
rect 28540 38412 28592 38418
rect 28264 38208 28316 38214
rect 28264 38150 28316 38156
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 27988 36576 28040 36582
rect 27988 36518 28040 36524
rect 28080 36576 28132 36582
rect 28080 36518 28132 36524
rect 28092 36394 28120 36518
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 27908 36366 28120 36394
rect 27908 36242 27936 36366
rect 27896 36236 27948 36242
rect 27896 36178 27948 36184
rect 28080 36236 28132 36242
rect 28080 36178 28132 36184
rect 27712 36168 27764 36174
rect 27712 36110 27764 36116
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27448 30802 27476 35974
rect 27632 35834 27660 36042
rect 27724 35834 27752 36110
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 27620 35828 27672 35834
rect 27620 35770 27672 35776
rect 27712 35828 27764 35834
rect 27908 35816 27936 36042
rect 27712 35770 27764 35776
rect 27816 35788 27936 35816
rect 27712 35692 27764 35698
rect 27712 35634 27764 35640
rect 27724 35136 27752 35634
rect 27816 35290 27844 35788
rect 27986 35728 28042 35737
rect 27896 35692 27948 35698
rect 27986 35663 28042 35672
rect 27896 35634 27948 35640
rect 27908 35290 27936 35634
rect 28000 35562 28028 35663
rect 27988 35556 28040 35562
rect 27988 35498 28040 35504
rect 27804 35284 27856 35290
rect 27804 35226 27856 35232
rect 27896 35284 27948 35290
rect 27896 35226 27948 35232
rect 27988 35216 28040 35222
rect 27908 35164 27988 35170
rect 27908 35158 28040 35164
rect 27908 35142 28028 35158
rect 27724 35108 27844 35136
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27620 35080 27672 35086
rect 27816 35068 27844 35108
rect 27908 35068 27936 35142
rect 27672 35040 27752 35068
rect 27620 35022 27672 35028
rect 27540 33998 27568 35022
rect 27620 34944 27672 34950
rect 27620 34886 27672 34892
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27540 33862 27568 33934
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27632 33538 27660 34886
rect 27724 34542 27752 35040
rect 27816 35040 27936 35068
rect 27816 34542 27844 35040
rect 28092 34678 28120 36178
rect 28170 34776 28226 34785
rect 28170 34711 28172 34720
rect 28224 34711 28226 34720
rect 28172 34682 28224 34688
rect 28080 34672 28132 34678
rect 28080 34614 28132 34620
rect 27712 34536 27764 34542
rect 27712 34478 27764 34484
rect 27804 34536 27856 34542
rect 27804 34478 27856 34484
rect 27540 33510 27660 33538
rect 27540 33454 27568 33510
rect 27528 33448 27580 33454
rect 27528 33390 27580 33396
rect 27620 33448 27672 33454
rect 27620 33390 27672 33396
rect 27632 33114 27660 33390
rect 27620 33108 27672 33114
rect 27620 33050 27672 33056
rect 27724 32570 27752 34478
rect 27988 34128 28040 34134
rect 27988 34070 28040 34076
rect 27896 33856 27948 33862
rect 27896 33798 27948 33804
rect 27804 33312 27856 33318
rect 27802 33280 27804 33289
rect 27856 33280 27858 33289
rect 27802 33215 27858 33224
rect 27528 32564 27580 32570
rect 27528 32506 27580 32512
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27540 32434 27568 32506
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27712 32292 27764 32298
rect 27712 32234 27764 32240
rect 27724 32026 27752 32234
rect 27712 32020 27764 32026
rect 27712 31962 27764 31968
rect 27908 31822 27936 33798
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 27436 30796 27488 30802
rect 27436 30738 27488 30744
rect 28000 30682 28028 34070
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 28092 33318 28120 33934
rect 28080 33312 28132 33318
rect 28080 33254 28132 33260
rect 28092 32230 28120 33254
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 28092 31346 28120 32166
rect 28184 31822 28212 34682
rect 28276 34490 28304 38150
rect 28368 35766 28396 38383
rect 28540 38354 28592 38360
rect 28448 38344 28500 38350
rect 28448 38286 28500 38292
rect 28460 37330 28488 38286
rect 28552 37913 28580 38354
rect 28538 37904 28594 37913
rect 28644 37874 28672 40967
rect 28814 40967 28870 40976
rect 28724 40938 28776 40944
rect 28736 40662 28764 40938
rect 28816 40928 28868 40934
rect 28816 40870 28868 40876
rect 28724 40656 28776 40662
rect 28724 40598 28776 40604
rect 28828 40526 28856 40870
rect 28906 40760 28962 40769
rect 28906 40695 28908 40704
rect 28960 40695 28962 40704
rect 28908 40666 28960 40672
rect 28908 40588 28960 40594
rect 28908 40530 28960 40536
rect 28724 40520 28776 40526
rect 28724 40462 28776 40468
rect 28816 40520 28868 40526
rect 28816 40462 28868 40468
rect 28736 38826 28764 40462
rect 28816 39976 28868 39982
rect 28814 39944 28816 39953
rect 28868 39944 28870 39953
rect 28814 39879 28870 39888
rect 28920 39828 28948 40530
rect 29012 40118 29040 41210
rect 29932 41002 29960 41482
rect 29920 40996 29972 41002
rect 29920 40938 29972 40944
rect 29932 40526 29960 40938
rect 29920 40520 29972 40526
rect 29920 40462 29972 40468
rect 29092 40452 29144 40458
rect 29092 40394 29144 40400
rect 29184 40452 29236 40458
rect 29184 40394 29236 40400
rect 29000 40112 29052 40118
rect 29000 40054 29052 40060
rect 28828 39800 28948 39828
rect 28828 39030 28856 39800
rect 29104 39506 29132 40394
rect 29196 40050 29224 40394
rect 29828 40384 29880 40390
rect 29828 40326 29880 40332
rect 29840 40118 29868 40326
rect 29828 40112 29880 40118
rect 29828 40054 29880 40060
rect 29184 40044 29236 40050
rect 29184 39986 29236 39992
rect 29092 39500 29144 39506
rect 29092 39442 29144 39448
rect 28816 39024 28868 39030
rect 28816 38966 28868 38972
rect 28906 38992 28962 39001
rect 28906 38927 28962 38936
rect 28724 38820 28776 38826
rect 28724 38762 28776 38768
rect 28920 38418 28948 38927
rect 29000 38752 29052 38758
rect 29000 38694 29052 38700
rect 29012 38486 29040 38694
rect 29000 38480 29052 38486
rect 29000 38422 29052 38428
rect 28908 38412 28960 38418
rect 28908 38354 28960 38360
rect 28538 37839 28594 37848
rect 28632 37868 28684 37874
rect 28632 37810 28684 37816
rect 28644 37754 28672 37810
rect 28552 37726 28672 37754
rect 28448 37324 28500 37330
rect 28448 37266 28500 37272
rect 28460 36174 28488 37266
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28356 35760 28408 35766
rect 28356 35702 28408 35708
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 28368 34610 28396 35566
rect 28460 35086 28488 36110
rect 28552 35154 28580 37726
rect 28632 37664 28684 37670
rect 28632 37606 28684 37612
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 28644 36378 28672 37606
rect 28736 37126 28764 37606
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28816 37120 28868 37126
rect 28816 37062 28868 37068
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 28540 35148 28592 35154
rect 28540 35090 28592 35096
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28460 34746 28488 35022
rect 28448 34740 28500 34746
rect 28448 34682 28500 34688
rect 28632 34672 28684 34678
rect 28632 34614 28684 34620
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28538 34504 28594 34513
rect 28276 34462 28396 34490
rect 28264 34196 28316 34202
rect 28264 34138 28316 34144
rect 28276 33114 28304 34138
rect 28264 33108 28316 33114
rect 28264 33050 28316 33056
rect 28276 32502 28304 33050
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28276 31346 28304 32302
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 27908 30654 28028 30682
rect 27252 29708 27304 29714
rect 27252 29650 27304 29656
rect 26884 28144 26936 28150
rect 26884 28086 26936 28092
rect 26988 27538 27016 29582
rect 27080 29566 27292 29594
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 27172 28490 27200 28698
rect 27160 28484 27212 28490
rect 27160 28426 27212 28432
rect 27172 28082 27200 28426
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 26976 27532 27028 27538
rect 26976 27474 27028 27480
rect 26792 26920 26844 26926
rect 26792 26862 26844 26868
rect 26804 26382 26832 26862
rect 26884 26852 26936 26858
rect 26884 26794 26936 26800
rect 26896 26450 26924 26794
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26988 26382 27016 27474
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26884 25764 26936 25770
rect 26884 25706 26936 25712
rect 26896 25226 26924 25706
rect 27080 25294 27108 27406
rect 27264 27316 27292 29566
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27448 27470 27476 28970
rect 27540 27470 27568 29514
rect 27908 29238 27936 30654
rect 27988 30592 28040 30598
rect 27988 30534 28040 30540
rect 28000 29646 28028 30534
rect 28078 30288 28134 30297
rect 28368 30258 28396 34462
rect 28538 34439 28594 34448
rect 28448 34400 28500 34406
rect 28448 34342 28500 34348
rect 28460 34202 28488 34342
rect 28448 34196 28500 34202
rect 28448 34138 28500 34144
rect 28446 33688 28502 33697
rect 28446 33623 28448 33632
rect 28500 33623 28502 33632
rect 28448 33594 28500 33600
rect 28552 33522 28580 34439
rect 28540 33516 28592 33522
rect 28540 33458 28592 33464
rect 28448 33380 28500 33386
rect 28448 33322 28500 33328
rect 28460 33289 28488 33322
rect 28644 33318 28672 34614
rect 28632 33312 28684 33318
rect 28446 33280 28502 33289
rect 28632 33254 28684 33260
rect 28446 33215 28502 33224
rect 28630 33144 28686 33153
rect 28630 33079 28686 33088
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28460 31822 28488 32370
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28540 31816 28592 31822
rect 28540 31758 28592 31764
rect 28552 30818 28580 31758
rect 28460 30790 28580 30818
rect 28460 30666 28488 30790
rect 28644 30682 28672 33079
rect 28736 32842 28764 37062
rect 28828 36718 28856 37062
rect 28816 36712 28868 36718
rect 28816 36654 28868 36660
rect 28920 36258 28948 38354
rect 29104 37262 29132 39442
rect 29644 38888 29696 38894
rect 29644 38830 29696 38836
rect 29656 38457 29684 38830
rect 29642 38448 29698 38457
rect 30024 38418 30052 42026
rect 30472 41676 30524 41682
rect 30472 41618 30524 41624
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 30196 41132 30248 41138
rect 30196 41074 30248 41080
rect 30116 40934 30144 41074
rect 30104 40928 30156 40934
rect 30104 40870 30156 40876
rect 30116 39438 30144 40870
rect 30208 40225 30236 41074
rect 30288 40588 30340 40594
rect 30288 40530 30340 40536
rect 30194 40216 30250 40225
rect 30194 40151 30250 40160
rect 30208 40050 30236 40151
rect 30300 40118 30328 40530
rect 30288 40112 30340 40118
rect 30288 40054 30340 40060
rect 30196 40044 30248 40050
rect 30196 39986 30248 39992
rect 30104 39432 30156 39438
rect 30104 39374 30156 39380
rect 30116 38826 30144 39374
rect 30484 39080 30512 41618
rect 30576 40662 30604 42162
rect 31576 42084 31628 42090
rect 31576 42026 31628 42032
rect 32588 42084 32640 42090
rect 32588 42026 32640 42032
rect 30840 41472 30892 41478
rect 30840 41414 30892 41420
rect 31116 41472 31168 41478
rect 31116 41414 31168 41420
rect 31588 41414 31616 42026
rect 31668 42016 31720 42022
rect 31668 41958 31720 41964
rect 31680 41546 31708 41958
rect 31668 41540 31720 41546
rect 31668 41482 31720 41488
rect 32496 41540 32548 41546
rect 32496 41482 32548 41488
rect 30852 41274 30880 41414
rect 31036 41386 31156 41414
rect 31588 41386 31708 41414
rect 30840 41268 30892 41274
rect 30840 41210 30892 41216
rect 31036 41138 31064 41386
rect 31680 41138 31708 41386
rect 32508 41138 32536 41482
rect 32600 41449 32628 42026
rect 33968 41608 34020 41614
rect 33968 41550 34020 41556
rect 33876 41472 33928 41478
rect 32586 41440 32642 41449
rect 33876 41414 33928 41420
rect 32586 41375 32642 41384
rect 31024 41132 31076 41138
rect 31024 41074 31076 41080
rect 31116 41132 31168 41138
rect 31116 41074 31168 41080
rect 31668 41132 31720 41138
rect 31668 41074 31720 41080
rect 32496 41132 32548 41138
rect 32496 41074 32548 41080
rect 33692 41132 33744 41138
rect 33692 41074 33744 41080
rect 30564 40656 30616 40662
rect 30564 40598 30616 40604
rect 30656 40520 30708 40526
rect 30656 40462 30708 40468
rect 30668 40390 30696 40462
rect 30656 40384 30708 40390
rect 30656 40326 30708 40332
rect 31036 40050 31064 41074
rect 31128 40594 31156 41074
rect 31680 40594 31708 41074
rect 32036 41064 32088 41070
rect 32036 41006 32088 41012
rect 31852 40928 31904 40934
rect 31852 40870 31904 40876
rect 31116 40588 31168 40594
rect 31116 40530 31168 40536
rect 31668 40588 31720 40594
rect 31668 40530 31720 40536
rect 31484 40384 31536 40390
rect 31484 40326 31536 40332
rect 31496 40050 31524 40326
rect 31024 40044 31076 40050
rect 31024 39986 31076 39992
rect 31484 40044 31536 40050
rect 31484 39986 31536 39992
rect 31300 39500 31352 39506
rect 31300 39442 31352 39448
rect 30564 39296 30616 39302
rect 30564 39238 30616 39244
rect 30392 39052 30512 39080
rect 30104 38820 30156 38826
rect 30104 38762 30156 38768
rect 29642 38383 29698 38392
rect 30012 38412 30064 38418
rect 30012 38354 30064 38360
rect 30116 38350 30144 38762
rect 30104 38344 30156 38350
rect 30104 38286 30156 38292
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 30012 37800 30064 37806
rect 30012 37742 30064 37748
rect 29092 37256 29144 37262
rect 29472 37233 29500 37742
rect 29552 37664 29604 37670
rect 29552 37606 29604 37612
rect 29092 37198 29144 37204
rect 29458 37224 29514 37233
rect 29104 37097 29132 37198
rect 29458 37159 29514 37168
rect 29090 37088 29146 37097
rect 29090 37023 29146 37032
rect 29368 36304 29420 36310
rect 28828 36230 29316 36258
rect 29368 36246 29420 36252
rect 28828 36174 28856 36230
rect 28816 36168 28868 36174
rect 28816 36110 28868 36116
rect 28908 36168 28960 36174
rect 28960 36128 29040 36156
rect 28908 36110 28960 36116
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 28816 35080 28868 35086
rect 28816 35022 28868 35028
rect 28828 33454 28856 35022
rect 28920 34950 28948 35702
rect 29012 35494 29040 36128
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 28908 34944 28960 34950
rect 28908 34886 28960 34892
rect 28920 34678 28948 34886
rect 29196 34678 29224 35974
rect 28908 34672 28960 34678
rect 28908 34614 28960 34620
rect 29184 34672 29236 34678
rect 29184 34614 29236 34620
rect 29092 34468 29144 34474
rect 29092 34410 29144 34416
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 29012 34066 29040 34342
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 28816 33448 28868 33454
rect 28816 33390 28868 33396
rect 28920 33114 28948 33458
rect 28908 33108 28960 33114
rect 28908 33050 28960 33056
rect 28724 32836 28776 32842
rect 28724 32778 28776 32784
rect 28816 32836 28868 32842
rect 28816 32778 28868 32784
rect 28828 32502 28856 32778
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 28828 32337 28856 32438
rect 29104 32434 29132 34410
rect 29288 34066 29316 36230
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28814 32328 28870 32337
rect 28814 32263 28870 32272
rect 29380 31754 29408 36246
rect 29564 35290 29592 37606
rect 29920 36712 29972 36718
rect 29920 36654 29972 36660
rect 29932 36310 29960 36654
rect 30024 36378 30052 37742
rect 30012 36372 30064 36378
rect 30012 36314 30064 36320
rect 29920 36304 29972 36310
rect 29920 36246 29972 36252
rect 30116 35698 30144 38286
rect 30392 38010 30420 39052
rect 30472 38956 30524 38962
rect 30472 38898 30524 38904
rect 30484 38350 30512 38898
rect 30472 38344 30524 38350
rect 30472 38286 30524 38292
rect 30380 38004 30432 38010
rect 30380 37946 30432 37952
rect 30196 37868 30248 37874
rect 30196 37810 30248 37816
rect 30380 37868 30432 37874
rect 30380 37810 30432 37816
rect 30208 37262 30236 37810
rect 30288 37664 30340 37670
rect 30288 37606 30340 37612
rect 30196 37256 30248 37262
rect 30196 37198 30248 37204
rect 30300 36378 30328 37606
rect 30392 36854 30420 37810
rect 30380 36848 30432 36854
rect 30380 36790 30432 36796
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 30300 36174 30328 36314
rect 30576 36174 30604 39238
rect 31312 39030 31340 39442
rect 31300 39024 31352 39030
rect 31300 38966 31352 38972
rect 31312 38758 31340 38966
rect 31300 38752 31352 38758
rect 31300 38694 31352 38700
rect 31024 38480 31076 38486
rect 31024 38422 31076 38428
rect 31036 36786 31064 38422
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 30748 36712 30800 36718
rect 30748 36654 30800 36660
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 30380 36168 30432 36174
rect 30380 36110 30432 36116
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30392 36020 30420 36110
rect 30760 36106 30788 36654
rect 31024 36236 31076 36242
rect 31024 36178 31076 36184
rect 30748 36100 30800 36106
rect 30748 36042 30800 36048
rect 30300 35992 30420 36020
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 29460 35080 29512 35086
rect 29460 35022 29512 35028
rect 29472 34542 29500 35022
rect 29564 35018 29592 35226
rect 29552 35012 29604 35018
rect 29552 34954 29604 34960
rect 29460 34536 29512 34542
rect 29460 34478 29512 34484
rect 29196 31726 29408 31754
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 29092 31680 29144 31686
rect 29092 31622 29144 31628
rect 29012 30734 29040 31622
rect 28448 30660 28500 30666
rect 28448 30602 28500 30608
rect 28552 30654 28672 30682
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 29104 30666 29132 31622
rect 29092 30660 29144 30666
rect 28078 30223 28080 30232
rect 28132 30223 28134 30232
rect 28356 30252 28408 30258
rect 28080 30194 28132 30200
rect 28356 30194 28408 30200
rect 28264 30116 28316 30122
rect 28264 30058 28316 30064
rect 27988 29640 28040 29646
rect 27988 29582 28040 29588
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28092 29306 28120 29582
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 27896 29232 27948 29238
rect 27896 29174 27948 29180
rect 28276 28694 28304 30058
rect 28368 29238 28396 30194
rect 28552 29322 28580 30654
rect 29092 30602 29144 30608
rect 28632 30592 28684 30598
rect 28632 30534 28684 30540
rect 28460 29294 28580 29322
rect 28644 29306 28672 30534
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28736 30122 28764 30194
rect 28724 30116 28776 30122
rect 28724 30058 28776 30064
rect 28736 29510 28764 30058
rect 28724 29504 28776 29510
rect 28724 29446 28776 29452
rect 28632 29300 28684 29306
rect 28356 29232 28408 29238
rect 28356 29174 28408 29180
rect 28460 29102 28488 29294
rect 28632 29242 28684 29248
rect 28736 29238 28764 29446
rect 28724 29232 28776 29238
rect 28724 29174 28776 29180
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28448 29096 28500 29102
rect 28448 29038 28500 29044
rect 27620 28688 27672 28694
rect 27620 28630 27672 28636
rect 28264 28688 28316 28694
rect 28264 28630 28316 28636
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27344 27328 27396 27334
rect 27264 27288 27344 27316
rect 27344 27270 27396 27276
rect 27252 27056 27304 27062
rect 27252 26998 27304 27004
rect 27264 26042 27292 26998
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27356 25922 27384 27270
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27264 25894 27384 25922
rect 27264 25838 27292 25894
rect 27252 25832 27304 25838
rect 27252 25774 27304 25780
rect 27342 25528 27398 25537
rect 27342 25463 27398 25472
rect 27356 25294 27384 25463
rect 27448 25378 27476 26318
rect 27540 25537 27568 27406
rect 27526 25528 27582 25537
rect 27526 25463 27582 25472
rect 27448 25350 27568 25378
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 26884 25220 26936 25226
rect 26884 25162 26936 25168
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26988 23866 27016 25094
rect 27080 24206 27108 25230
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26700 23792 26752 23798
rect 26700 23734 26752 23740
rect 26608 23248 26660 23254
rect 26608 23190 26660 23196
rect 26988 23186 27016 23802
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 27080 22642 27108 24142
rect 27160 23792 27212 23798
rect 27160 23734 27212 23740
rect 27172 23662 27200 23734
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27264 23526 27292 24346
rect 27356 24206 27384 25230
rect 27540 24206 27568 25350
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27264 23118 27292 23462
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 26056 22568 26108 22574
rect 26056 22510 26108 22516
rect 25792 22066 25912 22094
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25608 21690 25636 21898
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25608 21350 25636 21422
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25700 21146 25728 21490
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25516 19514 25544 19790
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25700 19446 25728 20402
rect 25688 19440 25740 19446
rect 25688 19382 25740 19388
rect 25412 18896 25464 18902
rect 25412 18838 25464 18844
rect 25700 18766 25728 19382
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25700 18290 25728 18702
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25792 17270 25820 22066
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25884 21554 25912 21830
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25884 21010 25912 21490
rect 25872 21004 25924 21010
rect 25872 20946 25924 20952
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 25884 19242 25912 20810
rect 26068 20466 26096 22510
rect 27080 22030 27108 22578
rect 27448 22438 27476 23122
rect 27436 22432 27488 22438
rect 27436 22374 27488 22380
rect 27632 22094 27660 28630
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 28000 28218 28028 28494
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 27712 28144 27764 28150
rect 27712 28086 27764 28092
rect 27724 27878 27752 28086
rect 28460 28014 28488 29038
rect 28552 28014 28580 29106
rect 28630 28520 28686 28529
rect 28630 28455 28686 28464
rect 28644 28150 28672 28455
rect 28632 28144 28684 28150
rect 28632 28086 28684 28092
rect 28644 28014 28672 28086
rect 28356 28008 28408 28014
rect 28356 27950 28408 27956
rect 28448 28008 28500 28014
rect 28448 27950 28500 27956
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 28632 28008 28684 28014
rect 28632 27950 28684 27956
rect 27712 27872 27764 27878
rect 27712 27814 27764 27820
rect 27804 27872 27856 27878
rect 27804 27814 27856 27820
rect 27724 27470 27752 27814
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27724 25498 27752 25842
rect 27712 25492 27764 25498
rect 27712 25434 27764 25440
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27724 24274 27752 24618
rect 27712 24268 27764 24274
rect 27712 24210 27764 24216
rect 27712 24132 27764 24138
rect 27712 24074 27764 24080
rect 27724 22642 27752 24074
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27540 22066 27660 22094
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26988 20942 27016 21830
rect 27080 21486 27108 21966
rect 27540 21690 27568 22066
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 27080 20466 27108 21422
rect 27436 21072 27488 21078
rect 27436 21014 27488 21020
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27264 19854 27292 20198
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26068 19378 26096 19654
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 26068 18970 26096 19314
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24688 16590 24716 16934
rect 26344 16794 26372 17614
rect 27160 17604 27212 17610
rect 27160 17546 27212 17552
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27172 17338 27200 17546
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 26344 15502 26372 16730
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 24308 15428 24360 15434
rect 24308 15370 24360 15376
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 22020 11234 22048 12786
rect 22664 12442 22692 12786
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11762 23152 12038
rect 23216 11898 23244 13194
rect 23400 12986 23428 13942
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23492 13530 23520 13874
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23676 13462 23704 14214
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23400 12238 23428 12922
rect 23676 12714 23704 13398
rect 23952 13326 23980 14758
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 14074 25176 14282
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24688 12850 24716 13670
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 24780 12374 24808 13874
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24872 12442 24900 12786
rect 25148 12646 25176 13738
rect 25332 13394 25360 15370
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25516 14074 25544 14214
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 12238 24808 12310
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 21928 11206 22048 11234
rect 21928 11150 21956 11206
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 22756 11082 22784 11494
rect 23216 11354 23244 11834
rect 25148 11694 25176 12582
rect 25332 12238 25360 13330
rect 25608 13190 25636 14418
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26160 13326 26188 14350
rect 26988 14346 27016 16730
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 14550 27108 16390
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15434 27200 15846
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27068 14544 27120 14550
rect 27068 14486 27120 14492
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26620 13870 26648 14214
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26424 13796 26476 13802
rect 26424 13738 26476 13744
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25608 12238 25636 13126
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25700 12238 25728 12650
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 24688 11150 24716 11494
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 25884 10674 25912 11494
rect 26160 11218 26188 13262
rect 26436 12374 26464 13738
rect 26988 12850 27016 14282
rect 27080 14074 27108 14350
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27264 13802 27292 17546
rect 27448 17270 27476 21014
rect 27540 20806 27568 21490
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27540 17338 27568 17478
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 27448 16250 27476 17206
rect 27632 16658 27660 21966
rect 27724 21894 27752 22578
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27724 21554 27752 21830
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27816 21162 27844 27814
rect 28262 27568 28318 27577
rect 28262 27503 28318 27512
rect 28276 27130 28304 27503
rect 28368 27130 28396 27950
rect 28736 27826 28764 29174
rect 28908 28620 28960 28626
rect 28908 28562 28960 28568
rect 28552 27798 28764 27826
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 28264 27124 28316 27130
rect 28264 27066 28316 27072
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 27896 26240 27948 26246
rect 27894 26208 27896 26217
rect 27948 26208 27950 26217
rect 27894 26143 27950 26152
rect 27908 25702 27936 26143
rect 27896 25696 27948 25702
rect 27896 25638 27948 25644
rect 27908 25294 27936 25638
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 28000 25106 28028 27066
rect 28552 26994 28580 27798
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 28080 26580 28132 26586
rect 28080 26522 28132 26528
rect 28092 26450 28120 26522
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28552 26314 28580 26930
rect 28540 26308 28592 26314
rect 28540 26250 28592 26256
rect 28632 26240 28684 26246
rect 28632 26182 28684 26188
rect 28080 25832 28132 25838
rect 28080 25774 28132 25780
rect 27908 25078 28028 25106
rect 27908 22642 27936 25078
rect 28092 24410 28120 25774
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28184 25226 28212 25298
rect 28172 25220 28224 25226
rect 28172 25162 28224 25168
rect 28540 24948 28592 24954
rect 28540 24890 28592 24896
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28092 23866 28120 24346
rect 28368 24206 28396 24754
rect 28552 24206 28580 24890
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28356 24200 28408 24206
rect 28540 24200 28592 24206
rect 28356 24142 28408 24148
rect 28538 24168 28540 24177
rect 28592 24168 28594 24177
rect 28276 23866 28304 24142
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28092 23662 28120 23802
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28184 23186 28212 23666
rect 28368 23526 28396 24142
rect 28538 24103 28594 24112
rect 28644 24070 28672 26182
rect 28828 26042 28856 26930
rect 28920 26926 28948 28562
rect 29090 27024 29146 27033
rect 29090 26959 29146 26968
rect 28908 26920 28960 26926
rect 28908 26862 28960 26868
rect 28908 26376 28960 26382
rect 28908 26318 28960 26324
rect 28920 26042 28948 26318
rect 28816 26036 28868 26042
rect 28816 25978 28868 25984
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 28920 23730 28948 24142
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 27908 22506 27936 22578
rect 27896 22500 27948 22506
rect 27896 22442 27948 22448
rect 28000 22030 28028 22714
rect 28184 22030 28212 23122
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28368 22710 28396 22986
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28632 22160 28684 22166
rect 28632 22102 28684 22108
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28276 21706 28304 21966
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 28092 21678 28304 21706
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27724 21134 27844 21162
rect 27724 17338 27752 21134
rect 27804 21072 27856 21078
rect 27804 21014 27856 21020
rect 27816 20874 27844 21014
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27908 20602 27936 21490
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 27816 19922 27844 20402
rect 27908 20398 27936 20538
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27356 13870 27384 14486
rect 27448 13938 27476 16186
rect 27540 16114 27568 16526
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27540 15706 27568 16050
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27816 14618 27844 19314
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13258 27200 13670
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26620 11762 26648 12174
rect 26804 11830 26832 12174
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26160 10742 26188 11154
rect 26620 10810 26648 11698
rect 26804 11354 26832 11766
rect 27356 11694 27384 13806
rect 27540 13530 27568 14010
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27816 12850 27844 14350
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27908 11898 27936 19654
rect 28000 14278 28028 21626
rect 28092 21622 28120 21678
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28080 20868 28132 20874
rect 28080 20810 28132 20816
rect 28092 20346 28120 20810
rect 28552 20466 28580 21422
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28092 20318 28488 20346
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28092 18154 28120 19790
rect 28184 18970 28212 19790
rect 28368 19378 28396 19994
rect 28460 19786 28488 20318
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 28460 19378 28488 19722
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28172 18964 28224 18970
rect 28172 18906 28224 18912
rect 28080 18148 28132 18154
rect 28080 18090 28132 18096
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28276 16658 28304 17750
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28368 16794 28396 17546
rect 28644 16794 28672 22102
rect 28920 22094 28948 22374
rect 28920 22066 29040 22094
rect 29012 21146 29040 22066
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 29104 20992 29132 26959
rect 29196 24274 29224 31726
rect 29368 31204 29420 31210
rect 29368 31146 29420 31152
rect 29276 30796 29328 30802
rect 29276 30738 29328 30744
rect 29288 30394 29316 30738
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 29380 30258 29408 31146
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29472 28558 29500 34478
rect 29656 34474 29684 35430
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29644 34468 29696 34474
rect 29644 34410 29696 34416
rect 29656 32774 29684 34410
rect 29932 33998 29960 35022
rect 30012 34400 30064 34406
rect 30012 34342 30064 34348
rect 29920 33992 29972 33998
rect 29920 33934 29972 33940
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29644 32768 29696 32774
rect 29644 32710 29696 32716
rect 29552 30388 29604 30394
rect 29552 30330 29604 30336
rect 29564 30258 29592 30330
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 29460 28552 29512 28558
rect 29460 28494 29512 28500
rect 29552 28416 29604 28422
rect 29552 28358 29604 28364
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29276 27396 29328 27402
rect 29276 27338 29328 27344
rect 29288 25242 29316 27338
rect 29380 26994 29408 28018
rect 29564 27606 29592 28358
rect 29656 28150 29684 32710
rect 29748 31822 29776 32914
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 29840 32570 29868 32846
rect 29828 32564 29880 32570
rect 29828 32506 29880 32512
rect 29840 31822 29868 32506
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29840 29170 29868 31758
rect 30024 31414 30052 34342
rect 30196 34128 30248 34134
rect 30196 34070 30248 34076
rect 30104 33856 30156 33862
rect 30104 33798 30156 33804
rect 30012 31408 30064 31414
rect 30012 31350 30064 31356
rect 30116 31346 30144 33798
rect 30208 33454 30236 34070
rect 30196 33448 30248 33454
rect 30196 33390 30248 33396
rect 30208 32978 30236 33390
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 30300 32910 30328 35992
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30392 35630 30420 35702
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 30380 35624 30432 35630
rect 30380 35566 30432 35572
rect 30392 34950 30420 35566
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30472 34944 30524 34950
rect 30472 34886 30524 34892
rect 30484 32910 30512 34886
rect 30576 33998 30604 35634
rect 30656 34944 30708 34950
rect 30656 34886 30708 34892
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30576 33522 30604 33798
rect 30668 33658 30696 34886
rect 30656 33652 30708 33658
rect 30656 33594 30708 33600
rect 30760 33522 30788 36042
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 30852 35222 30880 35566
rect 30932 35556 30984 35562
rect 30932 35498 30984 35504
rect 30944 35222 30972 35498
rect 30840 35216 30892 35222
rect 30840 35158 30892 35164
rect 30932 35216 30984 35222
rect 30932 35158 30984 35164
rect 30852 33998 30880 35158
rect 31036 34134 31064 36178
rect 31208 35624 31260 35630
rect 31208 35566 31260 35572
rect 31220 35290 31248 35566
rect 31208 35284 31260 35290
rect 31208 35226 31260 35232
rect 31312 34746 31340 38694
rect 31392 38344 31444 38350
rect 31392 38286 31444 38292
rect 31404 35222 31432 38286
rect 31496 37194 31524 39986
rect 31680 39642 31708 40530
rect 31864 40526 31892 40870
rect 32048 40526 32076 41006
rect 32508 40730 32536 41074
rect 32588 40996 32640 41002
rect 32588 40938 32640 40944
rect 32496 40724 32548 40730
rect 32496 40666 32548 40672
rect 31852 40520 31904 40526
rect 31852 40462 31904 40468
rect 32036 40520 32088 40526
rect 32036 40462 32088 40468
rect 31760 39840 31812 39846
rect 31760 39782 31812 39788
rect 31668 39636 31720 39642
rect 31668 39578 31720 39584
rect 31576 39432 31628 39438
rect 31576 39374 31628 39380
rect 31588 38350 31616 39374
rect 31680 38894 31708 39578
rect 31772 39370 31800 39782
rect 31760 39364 31812 39370
rect 31760 39306 31812 39312
rect 31772 38962 31800 39306
rect 31760 38956 31812 38962
rect 31760 38898 31812 38904
rect 31668 38888 31720 38894
rect 31720 38836 31800 38842
rect 31668 38830 31800 38836
rect 31680 38814 31800 38830
rect 31772 38350 31800 38814
rect 31576 38344 31628 38350
rect 31576 38286 31628 38292
rect 31760 38344 31812 38350
rect 31760 38286 31812 38292
rect 31668 38276 31720 38282
rect 31668 38218 31720 38224
rect 31680 37942 31708 38218
rect 31668 37936 31720 37942
rect 31668 37878 31720 37884
rect 31484 37188 31536 37194
rect 31484 37130 31536 37136
rect 31576 37188 31628 37194
rect 31680 37176 31708 37878
rect 31628 37148 31708 37176
rect 31576 37130 31628 37136
rect 31496 36582 31524 37130
rect 31680 36786 31708 37148
rect 31668 36780 31720 36786
rect 31668 36722 31720 36728
rect 31484 36576 31536 36582
rect 31484 36518 31536 36524
rect 31496 35698 31524 36518
rect 31680 36174 31708 36722
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 31484 35692 31536 35698
rect 31484 35634 31536 35640
rect 31772 35630 31800 38286
rect 31864 37330 31892 40462
rect 31944 39500 31996 39506
rect 31944 39442 31996 39448
rect 31956 38486 31984 39442
rect 32048 39438 32076 40462
rect 32128 40384 32180 40390
rect 32128 40326 32180 40332
rect 32036 39432 32088 39438
rect 32036 39374 32088 39380
rect 32140 39098 32168 40326
rect 32128 39092 32180 39098
rect 32128 39034 32180 39040
rect 31944 38480 31996 38486
rect 31944 38422 31996 38428
rect 32036 37664 32088 37670
rect 32036 37606 32088 37612
rect 31852 37324 31904 37330
rect 31852 37266 31904 37272
rect 31864 36224 31892 37266
rect 32048 37262 32076 37606
rect 32036 37256 32088 37262
rect 32034 37224 32036 37233
rect 32088 37224 32090 37233
rect 32140 37210 32168 39034
rect 32312 38956 32364 38962
rect 32312 38898 32364 38904
rect 32324 37874 32352 38898
rect 32404 38208 32456 38214
rect 32404 38150 32456 38156
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32416 37777 32444 38150
rect 32402 37768 32458 37777
rect 32402 37703 32458 37712
rect 32404 37664 32456 37670
rect 32404 37606 32456 37612
rect 32140 37182 32260 37210
rect 32034 37159 32090 37168
rect 31944 36236 31996 36242
rect 31864 36196 31944 36224
rect 31944 36178 31996 36184
rect 32128 36168 32180 36174
rect 32128 36110 32180 36116
rect 31944 35828 31996 35834
rect 31944 35770 31996 35776
rect 31760 35624 31812 35630
rect 31760 35566 31812 35572
rect 31392 35216 31444 35222
rect 31392 35158 31444 35164
rect 31404 35086 31432 35158
rect 31392 35080 31444 35086
rect 31392 35022 31444 35028
rect 31300 34740 31352 34746
rect 31300 34682 31352 34688
rect 31312 34610 31340 34682
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31404 34542 31432 35022
rect 31482 34776 31538 34785
rect 31482 34711 31484 34720
rect 31536 34711 31538 34720
rect 31484 34682 31536 34688
rect 31392 34536 31444 34542
rect 31392 34478 31444 34484
rect 31668 34196 31720 34202
rect 31668 34138 31720 34144
rect 31024 34128 31076 34134
rect 31024 34070 31076 34076
rect 30840 33992 30892 33998
rect 30840 33934 30892 33940
rect 31022 33960 31078 33969
rect 31022 33895 31078 33904
rect 31484 33924 31536 33930
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30748 33516 30800 33522
rect 30748 33458 30800 33464
rect 30748 33312 30800 33318
rect 30748 33254 30800 33260
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 30472 32904 30524 32910
rect 30472 32846 30524 32852
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30104 31340 30156 31346
rect 30104 31282 30156 31288
rect 30012 31204 30064 31210
rect 30012 31146 30064 31152
rect 30024 29782 30052 31146
rect 30012 29776 30064 29782
rect 30012 29718 30064 29724
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29552 27600 29604 27606
rect 29552 27542 29604 27548
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29288 25214 29408 25242
rect 29276 25152 29328 25158
rect 29276 25094 29328 25100
rect 29288 24750 29316 25094
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29184 24268 29236 24274
rect 29184 24210 29236 24216
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29196 23594 29224 23666
rect 29184 23588 29236 23594
rect 29184 23530 29236 23536
rect 29380 21418 29408 25214
rect 29472 24818 29500 26930
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29564 24698 29592 27542
rect 29748 27470 29776 28018
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 29748 26382 29776 27270
rect 29840 26994 29868 28494
rect 30024 27470 30052 29718
rect 30116 29714 30144 31282
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30300 30122 30328 30330
rect 30288 30116 30340 30122
rect 30288 30058 30340 30064
rect 30392 30054 30420 32302
rect 30656 31408 30708 31414
rect 30656 31350 30708 31356
rect 30668 30734 30696 31350
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30668 30258 30696 30670
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30380 30048 30432 30054
rect 30380 29990 30432 29996
rect 30104 29708 30156 29714
rect 30104 29650 30156 29656
rect 30380 29708 30432 29714
rect 30380 29650 30432 29656
rect 30392 28778 30420 29650
rect 30760 29617 30788 33254
rect 30840 32904 30892 32910
rect 30840 32846 30892 32852
rect 30852 32026 30880 32846
rect 30840 32020 30892 32026
rect 30840 31962 30892 31968
rect 30852 31346 30880 31962
rect 31036 31822 31064 33895
rect 31484 33866 31536 33872
rect 31392 33856 31444 33862
rect 31392 33798 31444 33804
rect 31116 33652 31168 33658
rect 31116 33594 31168 33600
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 30852 30734 30880 31282
rect 31022 31240 31078 31249
rect 31022 31175 31078 31184
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 30932 30660 30984 30666
rect 30932 30602 30984 30608
rect 30746 29608 30802 29617
rect 30746 29543 30802 29552
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30300 28750 30420 28778
rect 30300 28558 30328 28750
rect 30380 28688 30432 28694
rect 30380 28630 30432 28636
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 30012 27464 30064 27470
rect 29932 27412 30012 27418
rect 29932 27406 30064 27412
rect 29932 27390 30052 27406
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29840 26382 29868 26930
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29748 24750 29776 25230
rect 29472 24670 29592 24698
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29368 21412 29420 21418
rect 29368 21354 29420 21360
rect 29380 21078 29408 21354
rect 29472 21078 29500 24670
rect 29748 24274 29776 24686
rect 29736 24268 29788 24274
rect 29736 24210 29788 24216
rect 29552 22500 29604 22506
rect 29552 22442 29604 22448
rect 29368 21072 29420 21078
rect 29368 21014 29420 21020
rect 29460 21072 29512 21078
rect 29460 21014 29512 21020
rect 28920 20964 29132 20992
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28736 20466 28764 20538
rect 28920 20466 28948 20964
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28920 19990 28948 20402
rect 29472 20058 29500 21014
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29460 19848 29512 19854
rect 29460 19790 29512 19796
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28736 19514 28764 19654
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28736 18902 28764 19450
rect 28920 19378 28948 19450
rect 29104 19446 29132 19790
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28736 18290 28764 18838
rect 28920 18766 28948 19314
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29012 18834 29040 19246
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 29012 18426 29040 18770
rect 29104 18698 29132 19246
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 29000 18420 29052 18426
rect 29000 18362 29052 18368
rect 29104 18358 29132 18634
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29368 18216 29420 18222
rect 29368 18158 29420 18164
rect 29380 17746 29408 18158
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 28184 14006 28212 16390
rect 28552 15026 28580 16594
rect 29104 16522 29132 16934
rect 29092 16516 29144 16522
rect 29092 16458 29144 16464
rect 29472 16182 29500 19790
rect 29460 16176 29512 16182
rect 29460 16118 29512 16124
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28172 14000 28224 14006
rect 28172 13942 28224 13948
rect 28552 13734 28580 14962
rect 28736 13870 28764 15438
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28552 13326 28580 13670
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 27896 11892 27948 11898
rect 27896 11834 27948 11840
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 28092 11150 28120 11494
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 28276 10266 28304 10610
rect 28264 10260 28316 10266
rect 28264 10202 28316 10208
rect 28552 10130 28580 11766
rect 28644 10198 28672 12106
rect 28736 10742 28764 13806
rect 28828 12238 28856 14758
rect 29012 14346 29040 15506
rect 29000 14340 29052 14346
rect 29000 14282 29052 14288
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 29196 14006 29224 14214
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28828 11898 28856 12038
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 28828 11354 28856 11834
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28920 10810 28948 12106
rect 29012 11218 29040 13670
rect 29564 12850 29592 22442
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29656 20942 29684 21830
rect 29736 21140 29788 21146
rect 29736 21082 29788 21088
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29656 20058 29684 20878
rect 29644 20052 29696 20058
rect 29644 19994 29696 20000
rect 29656 19378 29684 19994
rect 29748 19922 29776 21082
rect 29932 20913 29960 27390
rect 30012 26512 30064 26518
rect 30012 26454 30064 26460
rect 30024 22098 30052 26454
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 30104 25220 30156 25226
rect 30104 25162 30156 25168
rect 30116 24818 30144 25162
rect 30104 24812 30156 24818
rect 30104 24754 30156 24760
rect 30116 24410 30144 24754
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 30116 24206 30144 24346
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30116 23526 30144 24142
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 30104 23248 30156 23254
rect 30104 23190 30156 23196
rect 30116 22642 30144 23190
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 30012 20936 30064 20942
rect 29918 20904 29974 20913
rect 30012 20878 30064 20884
rect 29918 20839 29974 20848
rect 29932 20806 29960 20839
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29748 15094 29776 15302
rect 29736 15088 29788 15094
rect 29736 15030 29788 15036
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29748 14414 29776 14894
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 13326 29776 14350
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29748 12918 29776 13262
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 29840 11898 29868 20198
rect 29932 19922 29960 20538
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29932 19514 29960 19858
rect 30024 19854 30052 20878
rect 30116 20534 30144 22374
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30116 20369 30144 20470
rect 30102 20360 30158 20369
rect 30102 20295 30158 20304
rect 30012 19848 30064 19854
rect 30012 19790 30064 19796
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 30116 19310 30144 19790
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30208 18358 30236 26386
rect 30286 26344 30342 26353
rect 30286 26279 30288 26288
rect 30340 26279 30342 26288
rect 30288 26250 30340 26256
rect 30288 25152 30340 25158
rect 30288 25094 30340 25100
rect 30300 24138 30328 25094
rect 30288 24132 30340 24138
rect 30288 24074 30340 24080
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30300 23118 30328 23258
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30300 22642 30328 23054
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30300 22030 30328 22578
rect 30392 22574 30420 28630
rect 30484 28558 30512 29446
rect 30760 29170 30788 29543
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30840 28552 30892 28558
rect 30840 28494 30892 28500
rect 30852 28082 30880 28494
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30564 27600 30616 27606
rect 30564 27542 30616 27548
rect 30576 27130 30604 27542
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30472 27056 30524 27062
rect 30472 26998 30524 27004
rect 30484 26489 30512 26998
rect 30470 26480 30526 26489
rect 30470 26415 30526 26424
rect 30576 25378 30604 27066
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30668 25906 30696 26998
rect 30852 26994 30880 27814
rect 30944 27470 30972 30602
rect 31036 27606 31064 31175
rect 31128 31142 31156 33594
rect 31404 33522 31432 33798
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31220 32026 31248 33458
rect 31312 32298 31340 33458
rect 31496 32434 31524 33866
rect 31576 33516 31628 33522
rect 31576 33458 31628 33464
rect 31588 32502 31616 33458
rect 31680 33386 31708 34138
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 33658 31800 33934
rect 31956 33862 31984 35770
rect 32036 35624 32088 35630
rect 32036 35566 32088 35572
rect 32048 35086 32076 35566
rect 32140 35494 32168 36110
rect 32128 35488 32180 35494
rect 32128 35430 32180 35436
rect 32140 35154 32168 35430
rect 32128 35148 32180 35154
rect 32128 35090 32180 35096
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 31944 33856 31996 33862
rect 31944 33798 31996 33804
rect 31760 33652 31812 33658
rect 31760 33594 31812 33600
rect 31668 33380 31720 33386
rect 31668 33322 31720 33328
rect 31576 32496 31628 32502
rect 31576 32438 31628 32444
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31300 32292 31352 32298
rect 31300 32234 31352 32240
rect 31208 32020 31260 32026
rect 31208 31962 31260 31968
rect 31116 31136 31168 31142
rect 31116 31078 31168 31084
rect 31128 30394 31156 31078
rect 31576 30932 31628 30938
rect 31576 30874 31628 30880
rect 31484 30592 31536 30598
rect 31484 30534 31536 30540
rect 31116 30388 31168 30394
rect 31116 30330 31168 30336
rect 31114 29744 31170 29753
rect 31114 29679 31170 29688
rect 31300 29708 31352 29714
rect 31128 29578 31156 29679
rect 31300 29650 31352 29656
rect 31116 29572 31168 29578
rect 31116 29514 31168 29520
rect 31208 29572 31260 29578
rect 31208 29514 31260 29520
rect 31116 29300 31168 29306
rect 31116 29242 31168 29248
rect 31128 29170 31156 29242
rect 31116 29164 31168 29170
rect 31116 29106 31168 29112
rect 31024 27600 31076 27606
rect 31024 27542 31076 27548
rect 30932 27464 30984 27470
rect 30984 27424 31064 27452
rect 30932 27406 30984 27412
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 30944 26994 30972 27270
rect 31036 27130 31064 27424
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 31128 26466 31156 29106
rect 31220 28558 31248 29514
rect 31312 29209 31340 29650
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31298 29200 31354 29209
rect 31298 29135 31354 29144
rect 31312 29102 31340 29135
rect 31300 29096 31352 29102
rect 31404 29073 31432 29582
rect 31496 29170 31524 30534
rect 31588 29714 31616 30874
rect 31680 30190 31708 33322
rect 31852 32292 31904 32298
rect 31852 32234 31904 32240
rect 31758 30560 31814 30569
rect 31758 30495 31814 30504
rect 31668 30184 31720 30190
rect 31668 30126 31720 30132
rect 31772 29753 31800 30495
rect 31758 29744 31814 29753
rect 31576 29708 31628 29714
rect 31758 29679 31814 29688
rect 31576 29650 31628 29656
rect 31588 29458 31616 29650
rect 31772 29578 31800 29679
rect 31864 29646 31892 32234
rect 32232 31754 32260 37182
rect 32416 33930 32444 37606
rect 32508 37262 32536 40666
rect 32600 40662 32628 40938
rect 33508 40928 33560 40934
rect 33508 40870 33560 40876
rect 32588 40656 32640 40662
rect 32588 40598 32640 40604
rect 33048 40520 33100 40526
rect 33048 40462 33100 40468
rect 32772 39976 32824 39982
rect 32772 39918 32824 39924
rect 32864 39976 32916 39982
rect 32864 39918 32916 39924
rect 32784 39098 32812 39918
rect 32876 39370 32904 39918
rect 33060 39642 33088 40462
rect 33520 40118 33548 40870
rect 33600 40520 33652 40526
rect 33600 40462 33652 40468
rect 33508 40112 33560 40118
rect 33508 40054 33560 40060
rect 33612 39930 33640 40462
rect 33704 40186 33732 41074
rect 33784 40452 33836 40458
rect 33784 40394 33836 40400
rect 33692 40180 33744 40186
rect 33692 40122 33744 40128
rect 33796 39953 33824 40394
rect 33520 39902 33640 39930
rect 33782 39944 33838 39953
rect 33048 39636 33100 39642
rect 33048 39578 33100 39584
rect 32864 39364 32916 39370
rect 32864 39306 32916 39312
rect 32772 39092 32824 39098
rect 32772 39034 32824 39040
rect 32680 38820 32732 38826
rect 32680 38762 32732 38768
rect 32692 38350 32720 38762
rect 32680 38344 32732 38350
rect 32680 38286 32732 38292
rect 32772 38344 32824 38350
rect 32772 38286 32824 38292
rect 32496 37256 32548 37262
rect 32680 37256 32732 37262
rect 32548 37216 32628 37244
rect 32496 37198 32548 37204
rect 32600 36786 32628 37216
rect 32680 37198 32732 37204
rect 32588 36780 32640 36786
rect 32588 36722 32640 36728
rect 32600 36174 32628 36722
rect 32692 36310 32720 37198
rect 32784 37126 32812 38286
rect 32876 38214 32904 39306
rect 33048 38752 33100 38758
rect 33048 38694 33100 38700
rect 33060 38350 33088 38694
rect 33048 38344 33100 38350
rect 33048 38286 33100 38292
rect 32864 38208 32916 38214
rect 32864 38150 32916 38156
rect 32772 37120 32824 37126
rect 32772 37062 32824 37068
rect 32680 36304 32732 36310
rect 32680 36246 32732 36252
rect 32588 36168 32640 36174
rect 32588 36110 32640 36116
rect 32772 36032 32824 36038
rect 32772 35974 32824 35980
rect 32680 35760 32732 35766
rect 32680 35702 32732 35708
rect 32588 35284 32640 35290
rect 32588 35226 32640 35232
rect 32600 34746 32628 35226
rect 32588 34740 32640 34746
rect 32588 34682 32640 34688
rect 32692 34626 32720 35702
rect 32784 35154 32812 35974
rect 32772 35148 32824 35154
rect 32772 35090 32824 35096
rect 32600 34598 32720 34626
rect 32496 34536 32548 34542
rect 32496 34478 32548 34484
rect 32404 33924 32456 33930
rect 32404 33866 32456 33872
rect 32416 32842 32444 33866
rect 32508 33590 32536 34478
rect 32496 33584 32548 33590
rect 32496 33526 32548 33532
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32494 32600 32550 32609
rect 32494 32535 32550 32544
rect 32508 32502 32536 32535
rect 32496 32496 32548 32502
rect 32496 32438 32548 32444
rect 32508 31890 32536 32438
rect 32496 31884 32548 31890
rect 32496 31826 32548 31832
rect 32232 31726 32444 31754
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32324 30666 32352 31418
rect 32416 31346 32444 31726
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32324 30190 32352 30602
rect 32416 30258 32444 31282
rect 32404 30252 32456 30258
rect 32404 30194 32456 30200
rect 32312 30184 32364 30190
rect 32312 30126 32364 30132
rect 32402 30152 32458 30161
rect 32128 29844 32180 29850
rect 32128 29786 32180 29792
rect 32140 29646 32168 29786
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 31760 29572 31812 29578
rect 31760 29514 31812 29520
rect 31588 29430 31800 29458
rect 31484 29164 31536 29170
rect 31484 29106 31536 29112
rect 31300 29038 31352 29044
rect 31390 29064 31446 29073
rect 31208 28552 31260 28558
rect 31208 28494 31260 28500
rect 31208 28416 31260 28422
rect 31208 28358 31260 28364
rect 31036 26438 31156 26466
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30748 25968 30800 25974
rect 30746 25936 30748 25945
rect 30800 25936 30802 25945
rect 30656 25900 30708 25906
rect 30746 25871 30802 25880
rect 30656 25842 30708 25848
rect 30840 25424 30892 25430
rect 30576 25350 30696 25378
rect 30840 25366 30892 25372
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30484 24750 30512 25162
rect 30576 24818 30604 25230
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 30484 24070 30512 24686
rect 30668 24682 30696 25350
rect 30852 24818 30880 25366
rect 30944 25294 30972 26182
rect 31036 25702 31064 26438
rect 31220 26382 31248 28358
rect 31312 26518 31340 29038
rect 31772 29050 31800 29430
rect 31390 28999 31446 29008
rect 31588 29022 31800 29050
rect 31300 26512 31352 26518
rect 31300 26454 31352 26460
rect 31208 26376 31260 26382
rect 31208 26318 31260 26324
rect 31116 26308 31168 26314
rect 31116 26250 31168 26256
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30656 24676 30708 24682
rect 30656 24618 30708 24624
rect 30760 24410 30788 24754
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30852 24070 30880 24550
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30484 23730 30512 24006
rect 30472 23724 30524 23730
rect 30472 23666 30524 23672
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30484 21486 30512 23666
rect 30576 23594 30604 23666
rect 30564 23588 30616 23594
rect 30564 23530 30616 23536
rect 30944 23526 30972 24074
rect 30932 23520 30984 23526
rect 30932 23462 30984 23468
rect 30840 22976 30892 22982
rect 30840 22918 30892 22924
rect 30852 22642 30880 22918
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30930 21992 30986 22001
rect 30930 21927 30932 21936
rect 30984 21927 30986 21936
rect 30932 21898 30984 21904
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30380 21140 30432 21146
rect 30380 21082 30432 21088
rect 30288 21072 30340 21078
rect 30288 21014 30340 21020
rect 30300 20806 30328 21014
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30392 20602 30420 21082
rect 30380 20596 30432 20602
rect 30380 20538 30432 20544
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30668 20058 30696 20402
rect 30656 20052 30708 20058
rect 30656 19994 30708 20000
rect 30378 19952 30434 19961
rect 30378 19887 30434 19896
rect 30392 19786 30420 19887
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 29932 16046 29960 17274
rect 30024 16250 30052 17546
rect 30668 16590 30696 18294
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 30208 16182 30236 16458
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29932 15570 29960 15982
rect 30104 15972 30156 15978
rect 30104 15914 30156 15920
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 30116 15502 30144 15914
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 30116 15162 30144 15438
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30208 14346 30236 16118
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 30196 14340 30248 14346
rect 30196 14282 30248 14288
rect 29932 13258 29960 14282
rect 30300 14006 30328 16050
rect 30472 15564 30524 15570
rect 30472 15506 30524 15512
rect 30484 14346 30512 15506
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30576 14482 30604 14962
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 29920 13252 29972 13258
rect 29920 13194 29972 13200
rect 29932 12986 29960 13194
rect 29920 12980 29972 12986
rect 29920 12922 29972 12928
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 30300 11694 30328 13942
rect 30484 12646 30512 14282
rect 30576 14074 30604 14418
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 29000 11212 29052 11218
rect 29000 11154 29052 11160
rect 30104 11212 30156 11218
rect 30104 11154 30156 11160
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 28724 10736 28776 10742
rect 28724 10678 28776 10684
rect 28632 10192 28684 10198
rect 28632 10134 28684 10140
rect 28540 10124 28592 10130
rect 28540 10066 28592 10072
rect 28920 10062 28948 10746
rect 30116 10674 30144 11154
rect 30392 11150 30420 11494
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30392 10266 30420 10610
rect 30484 10282 30512 12582
rect 30576 12442 30604 12718
rect 30668 12442 30696 12786
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30380 10260 30432 10266
rect 30484 10254 30604 10282
rect 30380 10202 30432 10208
rect 30576 10198 30604 10254
rect 30564 10192 30616 10198
rect 30564 10134 30616 10140
rect 30944 10130 30972 11834
rect 31036 10742 31064 24550
rect 31128 22642 31156 26250
rect 31312 25974 31340 26454
rect 31300 25968 31352 25974
rect 31300 25910 31352 25916
rect 31208 25900 31260 25906
rect 31208 25842 31260 25848
rect 31220 24274 31248 25842
rect 31312 25430 31340 25910
rect 31404 25906 31432 28999
rect 31588 28558 31616 29022
rect 31666 28928 31722 28937
rect 31666 28863 31722 28872
rect 31576 28552 31628 28558
rect 31576 28494 31628 28500
rect 31680 28082 31708 28863
rect 31772 28150 31800 29022
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 32048 28558 32076 28902
rect 32036 28552 32088 28558
rect 31850 28520 31906 28529
rect 32036 28494 32088 28500
rect 31850 28455 31852 28464
rect 31904 28455 31906 28464
rect 31852 28426 31904 28432
rect 31760 28144 31812 28150
rect 31760 28086 31812 28092
rect 31668 28076 31720 28082
rect 31668 28018 31720 28024
rect 31576 27600 31628 27606
rect 31576 27542 31628 27548
rect 31484 26920 31536 26926
rect 31484 26862 31536 26868
rect 31496 26382 31524 26862
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31300 25424 31352 25430
rect 31300 25366 31352 25372
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31208 24268 31260 24274
rect 31208 24210 31260 24216
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 31220 23662 31248 23802
rect 31208 23656 31260 23662
rect 31208 23598 31260 23604
rect 31312 23594 31340 25230
rect 31404 25158 31432 25434
rect 31496 25294 31524 26318
rect 31588 26314 31616 27542
rect 31668 27464 31720 27470
rect 31668 27406 31720 27412
rect 31680 27130 31708 27406
rect 31772 27402 31800 28086
rect 31864 27577 31892 28426
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 31850 27568 31906 27577
rect 32048 27538 32076 27950
rect 31850 27503 31906 27512
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31668 27124 31720 27130
rect 31668 27066 31720 27072
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31392 25152 31444 25158
rect 31392 25094 31444 25100
rect 31404 24886 31432 25094
rect 31392 24880 31444 24886
rect 31392 24822 31444 24828
rect 31300 23588 31352 23594
rect 31300 23530 31352 23536
rect 31404 22778 31432 24822
rect 31576 24676 31628 24682
rect 31576 24618 31628 24624
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31116 22636 31168 22642
rect 31116 22578 31168 22584
rect 31116 22500 31168 22506
rect 31116 22442 31168 22448
rect 31128 22234 31156 22442
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31208 22092 31260 22098
rect 31404 22094 31432 22714
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31208 22034 31260 22040
rect 31312 22066 31432 22094
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 31128 21690 31156 21830
rect 31220 21729 31248 22034
rect 31206 21720 31262 21729
rect 31116 21684 31168 21690
rect 31206 21655 31262 21664
rect 31116 21626 31168 21632
rect 31220 21622 31248 21655
rect 31312 21622 31340 22066
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31300 21616 31352 21622
rect 31300 21558 31352 21564
rect 31116 21480 31168 21486
rect 31116 21422 31168 21428
rect 31128 19922 31156 21422
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31116 17536 31168 17542
rect 31116 17478 31168 17484
rect 31128 16658 31156 17478
rect 31208 17128 31260 17134
rect 31208 17070 31260 17076
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 31128 16250 31156 16594
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31128 15162 31156 16050
rect 31116 15156 31168 15162
rect 31116 15098 31168 15104
rect 31220 14822 31248 17070
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31404 15434 31432 16050
rect 31392 15428 31444 15434
rect 31392 15370 31444 15376
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 31404 12434 31432 14214
rect 31496 12918 31524 22510
rect 31588 21078 31616 24618
rect 31576 21072 31628 21078
rect 31576 21014 31628 21020
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 31588 19417 31616 20878
rect 31574 19408 31630 19417
rect 31574 19343 31630 19352
rect 31576 17128 31628 17134
rect 31576 17070 31628 17076
rect 31588 14346 31616 17070
rect 31680 16522 31708 27066
rect 31850 27024 31906 27033
rect 31850 26959 31852 26968
rect 31904 26959 31906 26968
rect 31852 26930 31904 26936
rect 31956 26926 31984 27474
rect 32034 27432 32090 27441
rect 32034 27367 32090 27376
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 31944 25696 31996 25702
rect 31944 25638 31996 25644
rect 31760 25424 31812 25430
rect 31760 25366 31812 25372
rect 31852 25424 31904 25430
rect 31852 25366 31904 25372
rect 31772 24818 31800 25366
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 31772 20942 31800 23258
rect 31864 21010 31892 25366
rect 31956 25362 31984 25638
rect 31944 25356 31996 25362
rect 31944 25298 31996 25304
rect 32048 23662 32076 27367
rect 32036 23656 32088 23662
rect 32036 23598 32088 23604
rect 32048 22094 32076 23598
rect 32140 22642 32168 29582
rect 32324 29306 32352 30126
rect 32402 30087 32458 30096
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32416 29238 32444 30087
rect 32404 29232 32456 29238
rect 32404 29174 32456 29180
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32508 28626 32536 28698
rect 32496 28620 32548 28626
rect 32496 28562 32548 28568
rect 32600 28558 32628 34598
rect 32784 34202 32812 35090
rect 32876 34406 32904 38150
rect 33324 37392 33376 37398
rect 33324 37334 33376 37340
rect 33046 37088 33102 37097
rect 33046 37023 33102 37032
rect 33060 36854 33088 37023
rect 33140 36916 33192 36922
rect 33140 36858 33192 36864
rect 33048 36848 33100 36854
rect 33048 36790 33100 36796
rect 33152 36174 33180 36858
rect 33232 36304 33284 36310
rect 33232 36246 33284 36252
rect 32956 36168 33008 36174
rect 32956 36110 33008 36116
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 32968 35154 32996 36110
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 32956 35148 33008 35154
rect 32956 35090 33008 35096
rect 33060 35034 33088 35770
rect 33152 35630 33180 36110
rect 33140 35624 33192 35630
rect 33140 35566 33192 35572
rect 32968 35006 33088 35034
rect 32864 34400 32916 34406
rect 32864 34342 32916 34348
rect 32772 34196 32824 34202
rect 32772 34138 32824 34144
rect 32968 34082 32996 35006
rect 33048 34944 33100 34950
rect 33048 34886 33100 34892
rect 33060 34746 33088 34886
rect 33048 34740 33100 34746
rect 33048 34682 33100 34688
rect 33140 34740 33192 34746
rect 33140 34682 33192 34688
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 32692 34054 32996 34082
rect 32220 28552 32272 28558
rect 32220 28494 32272 28500
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32232 25498 32260 28494
rect 32588 28076 32640 28082
rect 32692 28064 32720 34054
rect 32956 33652 33008 33658
rect 32956 33594 33008 33600
rect 32968 33402 32996 33594
rect 33060 33590 33088 34342
rect 33048 33584 33100 33590
rect 33048 33526 33100 33532
rect 33152 33436 33180 34682
rect 33244 34610 33272 36246
rect 33336 36106 33364 37334
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 33428 36650 33456 36722
rect 33416 36644 33468 36650
rect 33416 36586 33468 36592
rect 33428 36106 33456 36586
rect 33324 36100 33376 36106
rect 33324 36042 33376 36048
rect 33416 36100 33468 36106
rect 33416 36042 33468 36048
rect 33336 35986 33364 36042
rect 33336 35958 33456 35986
rect 33428 35698 33456 35958
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33416 35692 33468 35698
rect 33416 35634 33468 35640
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 32876 33374 32996 33402
rect 33060 33408 33180 33436
rect 32876 28490 32904 33374
rect 32956 31272 33008 31278
rect 32956 31214 33008 31220
rect 32968 30870 32996 31214
rect 32956 30864 33008 30870
rect 32956 30806 33008 30812
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32968 28762 32996 29582
rect 32956 28756 33008 28762
rect 32956 28698 33008 28704
rect 32864 28484 32916 28490
rect 32864 28426 32916 28432
rect 33060 28370 33088 33408
rect 33138 33144 33194 33153
rect 33138 33079 33194 33088
rect 33152 31958 33180 33079
rect 33336 32910 33364 35634
rect 33416 35080 33468 35086
rect 33416 35022 33468 35028
rect 33428 33844 33456 35022
rect 33520 33946 33548 39902
rect 33782 39879 33838 39888
rect 33796 39574 33824 39879
rect 33784 39568 33836 39574
rect 33784 39510 33836 39516
rect 33888 38962 33916 41414
rect 33980 41138 34008 41550
rect 33968 41132 34020 41138
rect 33968 41074 34020 41080
rect 34164 39438 34192 42162
rect 35624 42016 35676 42022
rect 35624 41958 35676 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34612 41676 34664 41682
rect 34612 41618 34664 41624
rect 34244 41608 34296 41614
rect 34244 41550 34296 41556
rect 34256 41206 34284 41550
rect 34244 41200 34296 41206
rect 34244 41142 34296 41148
rect 34244 40996 34296 41002
rect 34244 40938 34296 40944
rect 34060 39432 34112 39438
rect 34060 39374 34112 39380
rect 34152 39432 34204 39438
rect 34152 39374 34204 39380
rect 34072 39284 34100 39374
rect 34072 39256 34192 39284
rect 33968 39024 34020 39030
rect 33968 38966 34020 38972
rect 33784 38956 33836 38962
rect 33784 38898 33836 38904
rect 33876 38956 33928 38962
rect 33876 38898 33928 38904
rect 33796 38282 33824 38898
rect 33600 38276 33652 38282
rect 33600 38218 33652 38224
rect 33784 38276 33836 38282
rect 33784 38218 33836 38224
rect 33612 38010 33640 38218
rect 33600 38004 33652 38010
rect 33600 37946 33652 37952
rect 33796 37874 33824 38218
rect 33980 37874 34008 38966
rect 34164 37913 34192 39256
rect 34256 38350 34284 40938
rect 34624 40118 34652 41618
rect 35532 41608 35584 41614
rect 35532 41550 35584 41556
rect 35348 41540 35400 41546
rect 35348 41482 35400 41488
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40730 35388 41482
rect 35544 41138 35572 41550
rect 35636 41206 35664 41958
rect 38016 41540 38068 41546
rect 38016 41482 38068 41488
rect 35900 41472 35952 41478
rect 35900 41414 35952 41420
rect 35624 41200 35676 41206
rect 35624 41142 35676 41148
rect 35532 41132 35584 41138
rect 35532 41074 35584 41080
rect 35440 41064 35492 41070
rect 35440 41006 35492 41012
rect 35348 40724 35400 40730
rect 35348 40666 35400 40672
rect 34796 40520 34848 40526
rect 34796 40462 34848 40468
rect 34980 40520 35032 40526
rect 34980 40462 35032 40468
rect 34704 40180 34756 40186
rect 34704 40122 34756 40128
rect 34612 40112 34664 40118
rect 34612 40054 34664 40060
rect 34520 40044 34572 40050
rect 34520 39986 34572 39992
rect 34428 39840 34480 39846
rect 34428 39782 34480 39788
rect 34440 39438 34468 39782
rect 34532 39642 34560 39986
rect 34612 39840 34664 39846
rect 34612 39782 34664 39788
rect 34520 39636 34572 39642
rect 34520 39578 34572 39584
rect 34428 39432 34480 39438
rect 34428 39374 34480 39380
rect 34244 38344 34296 38350
rect 34244 38286 34296 38292
rect 34428 38344 34480 38350
rect 34428 38286 34480 38292
rect 34336 38004 34388 38010
rect 34336 37946 34388 37952
rect 34150 37904 34206 37913
rect 33784 37868 33836 37874
rect 33784 37810 33836 37816
rect 33968 37868 34020 37874
rect 34150 37839 34206 37848
rect 33968 37810 34020 37816
rect 33600 37800 33652 37806
rect 33600 37742 33652 37748
rect 33612 36786 33640 37742
rect 33796 37346 33824 37810
rect 33796 37318 34008 37346
rect 33980 37262 34008 37318
rect 33876 37256 33928 37262
rect 33874 37224 33876 37233
rect 33968 37256 34020 37262
rect 33928 37224 33930 37233
rect 33968 37198 34020 37204
rect 33874 37159 33930 37168
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33692 36032 33744 36038
rect 33692 35974 33744 35980
rect 33600 35488 33652 35494
rect 33600 35430 33652 35436
rect 33612 34406 33640 35430
rect 33704 34610 33732 35974
rect 33980 35086 34008 37198
rect 34060 36780 34112 36786
rect 34060 36722 34112 36728
rect 34072 36174 34100 36722
rect 34060 36168 34112 36174
rect 34060 36110 34112 36116
rect 34164 35578 34192 37839
rect 34244 37256 34296 37262
rect 34244 37198 34296 37204
rect 34256 36718 34284 37198
rect 34244 36712 34296 36718
rect 34244 36654 34296 36660
rect 34256 35698 34284 36654
rect 34348 35698 34376 37946
rect 34440 37942 34468 38286
rect 34520 38276 34572 38282
rect 34520 38218 34572 38224
rect 34428 37936 34480 37942
rect 34428 37878 34480 37884
rect 34428 37732 34480 37738
rect 34428 37674 34480 37680
rect 34440 36922 34468 37674
rect 34428 36916 34480 36922
rect 34428 36858 34480 36864
rect 34532 36802 34560 38218
rect 34440 36774 34560 36802
rect 34244 35692 34296 35698
rect 34244 35634 34296 35640
rect 34336 35692 34388 35698
rect 34336 35634 34388 35640
rect 34164 35550 34376 35578
rect 33968 35080 34020 35086
rect 33968 35022 34020 35028
rect 34244 34944 34296 34950
rect 34244 34886 34296 34892
rect 33692 34604 33744 34610
rect 33692 34546 33744 34552
rect 33600 34400 33652 34406
rect 33600 34342 33652 34348
rect 33704 34066 33732 34546
rect 33874 34504 33930 34513
rect 34256 34474 34284 34886
rect 33874 34439 33930 34448
rect 34152 34468 34204 34474
rect 33784 34196 33836 34202
rect 33784 34138 33836 34144
rect 33692 34060 33744 34066
rect 33692 34002 33744 34008
rect 33796 33969 33824 34138
rect 33782 33960 33838 33969
rect 33520 33918 33732 33946
rect 33600 33856 33652 33862
rect 33428 33816 33548 33844
rect 33416 33448 33468 33454
rect 33416 33390 33468 33396
rect 33428 32910 33456 33390
rect 33520 32978 33548 33816
rect 33600 33798 33652 33804
rect 33508 32972 33560 32978
rect 33508 32914 33560 32920
rect 33324 32904 33376 32910
rect 33324 32846 33376 32852
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33140 31952 33192 31958
rect 33140 31894 33192 31900
rect 33152 30734 33180 31894
rect 33232 31816 33284 31822
rect 33232 31758 33284 31764
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 33244 29850 33272 31758
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 33336 31346 33364 31690
rect 33428 31414 33456 32846
rect 33508 32428 33560 32434
rect 33508 32370 33560 32376
rect 33520 31958 33548 32370
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33416 31408 33468 31414
rect 33416 31350 33468 31356
rect 33324 31340 33376 31346
rect 33324 31282 33376 31288
rect 33508 30864 33560 30870
rect 33508 30806 33560 30812
rect 33416 30592 33468 30598
rect 33416 30534 33468 30540
rect 33428 30433 33456 30534
rect 33414 30424 33470 30433
rect 33414 30359 33470 30368
rect 33232 29844 33284 29850
rect 33232 29786 33284 29792
rect 33324 29844 33376 29850
rect 33324 29786 33376 29792
rect 33138 29744 33194 29753
rect 33138 29679 33194 29688
rect 33152 29646 33180 29679
rect 33140 29640 33192 29646
rect 33140 29582 33192 29588
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 33140 29164 33192 29170
rect 33140 29106 33192 29112
rect 33152 29073 33180 29106
rect 33138 29064 33194 29073
rect 33138 28999 33194 29008
rect 33244 28558 33272 29174
rect 33232 28552 33284 28558
rect 33232 28494 33284 28500
rect 33140 28484 33192 28490
rect 33140 28426 33192 28432
rect 32968 28342 33088 28370
rect 32968 28132 32996 28342
rect 32968 28104 33088 28132
rect 32772 28076 32824 28082
rect 32692 28036 32772 28064
rect 32588 28018 32640 28024
rect 32772 28018 32824 28024
rect 32600 27985 32628 28018
rect 32956 28008 33008 28014
rect 32586 27976 32642 27985
rect 32956 27950 33008 27956
rect 32586 27911 32642 27920
rect 32312 27872 32364 27878
rect 32312 27814 32364 27820
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32324 25294 32352 27814
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32220 24744 32272 24750
rect 32220 24686 32272 24692
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32048 22066 32168 22094
rect 32140 21049 32168 22066
rect 32232 21146 32260 24686
rect 32312 21956 32364 21962
rect 32312 21898 32364 21904
rect 32324 21486 32352 21898
rect 32312 21480 32364 21486
rect 32312 21422 32364 21428
rect 32220 21140 32272 21146
rect 32220 21082 32272 21088
rect 32126 21040 32182 21049
rect 31852 21004 31904 21010
rect 32126 20975 32182 20984
rect 31852 20946 31904 20952
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 31864 19854 31892 19926
rect 31760 19848 31812 19854
rect 31852 19848 31904 19854
rect 31760 19790 31812 19796
rect 31850 19816 31852 19825
rect 31904 19816 31906 19825
rect 31772 19514 31800 19790
rect 31850 19751 31906 19760
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 32140 19446 32168 20975
rect 32232 20262 32260 21082
rect 32416 21010 32444 27814
rect 32772 27668 32824 27674
rect 32772 27610 32824 27616
rect 32588 27532 32640 27538
rect 32588 27474 32640 27480
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32508 25294 32536 26930
rect 32600 26625 32628 27474
rect 32784 27418 32812 27610
rect 32968 27606 32996 27950
rect 32956 27600 33008 27606
rect 32956 27542 33008 27548
rect 32784 27390 32904 27418
rect 32772 27328 32824 27334
rect 32772 27270 32824 27276
rect 32586 26616 32642 26625
rect 32586 26551 32642 26560
rect 32784 26382 32812 27270
rect 32876 26382 32904 27390
rect 32956 27396 33008 27402
rect 32956 27338 33008 27344
rect 32968 26790 32996 27338
rect 32956 26784 33008 26790
rect 32956 26726 33008 26732
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32680 25968 32732 25974
rect 32680 25910 32732 25916
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32508 23322 32536 25230
rect 32692 25208 32720 25910
rect 32784 25906 32812 26318
rect 32956 26036 33008 26042
rect 32956 25978 33008 25984
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32772 25220 32824 25226
rect 32692 25180 32772 25208
rect 32692 24886 32720 25180
rect 32772 25162 32824 25168
rect 32680 24880 32732 24886
rect 32680 24822 32732 24828
rect 32862 24848 32918 24857
rect 32862 24783 32864 24792
rect 32916 24783 32918 24792
rect 32864 24754 32916 24760
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32600 23730 32628 24550
rect 32968 24138 32996 25978
rect 33060 25974 33088 28104
rect 33152 27470 33180 28426
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33140 27464 33192 27470
rect 33140 27406 33192 27412
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33152 26897 33180 26930
rect 33138 26888 33194 26897
rect 33138 26823 33194 26832
rect 33244 26466 33272 27950
rect 33152 26438 33272 26466
rect 33152 26246 33180 26438
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33140 26240 33192 26246
rect 33140 26182 33192 26188
rect 33152 25974 33180 26182
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 33140 25968 33192 25974
rect 33140 25910 33192 25916
rect 33244 25498 33272 26318
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 33336 24324 33364 29786
rect 33416 29640 33468 29646
rect 33414 29608 33416 29617
rect 33468 29608 33470 29617
rect 33414 29543 33470 29552
rect 33520 28150 33548 30806
rect 33508 28144 33560 28150
rect 33508 28086 33560 28092
rect 33520 27441 33548 28086
rect 33506 27432 33562 27441
rect 33506 27367 33562 27376
rect 33416 26784 33468 26790
rect 33416 26726 33468 26732
rect 33428 25906 33456 26726
rect 33508 26308 33560 26314
rect 33508 26250 33560 26256
rect 33416 25900 33468 25906
rect 33416 25842 33468 25848
rect 33520 24954 33548 26250
rect 33508 24948 33560 24954
rect 33508 24890 33560 24896
rect 33244 24296 33364 24324
rect 33048 24200 33100 24206
rect 33048 24142 33100 24148
rect 32956 24132 33008 24138
rect 32956 24074 33008 24080
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 33060 23526 33088 24142
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33048 23520 33100 23526
rect 33048 23462 33100 23468
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 33060 22098 33088 23258
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 33152 21434 33180 23802
rect 33244 22001 33272 24296
rect 33508 23520 33560 23526
rect 33508 23462 33560 23468
rect 33324 22976 33376 22982
rect 33324 22918 33376 22924
rect 33336 22710 33364 22918
rect 33324 22704 33376 22710
rect 33324 22646 33376 22652
rect 33230 21992 33286 22001
rect 33230 21927 33286 21936
rect 33336 21434 33364 22646
rect 33416 21956 33468 21962
rect 33416 21898 33468 21904
rect 33428 21554 33456 21898
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33152 21406 33272 21434
rect 33336 21406 33456 21434
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 32404 21004 32456 21010
rect 32404 20946 32456 20952
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32588 19780 32640 19786
rect 32588 19722 32640 19728
rect 32128 19440 32180 19446
rect 31758 19408 31814 19417
rect 32128 19382 32180 19388
rect 31758 19343 31814 19352
rect 31772 17746 31800 19343
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31760 17604 31812 17610
rect 31760 17546 31812 17552
rect 31772 17338 31800 17546
rect 31852 17536 31904 17542
rect 31852 17478 31904 17484
rect 31760 17332 31812 17338
rect 31760 17274 31812 17280
rect 31864 17202 31892 17478
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 31668 16516 31720 16522
rect 31668 16458 31720 16464
rect 31772 16250 31800 16526
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 32048 15366 32076 16526
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31680 14414 31708 14962
rect 32048 14890 32076 15302
rect 32324 14958 32352 16594
rect 32416 16590 32444 17138
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32036 14884 32088 14890
rect 32036 14826 32088 14832
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31576 14340 31628 14346
rect 31576 14282 31628 14288
rect 31484 12912 31536 12918
rect 31484 12854 31536 12860
rect 31588 12850 31616 14282
rect 31680 13938 31708 14350
rect 32048 13938 32076 14826
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 32036 13932 32088 13938
rect 32036 13874 32088 13880
rect 32324 13462 32352 14894
rect 32312 13456 32364 13462
rect 32312 13398 32364 13404
rect 32324 13190 32352 13398
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 31312 12406 31432 12434
rect 31312 12306 31340 12406
rect 31300 12300 31352 12306
rect 31300 12242 31352 12248
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31220 10810 31248 12038
rect 31312 11762 31340 12038
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 31312 11354 31340 11698
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 32416 11218 32444 12786
rect 32600 12306 32628 19722
rect 33048 16040 33100 16046
rect 33048 15982 33100 15988
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32772 14340 32824 14346
rect 32772 14282 32824 14288
rect 32784 14074 32812 14282
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32968 13326 32996 15438
rect 33060 15162 33088 15982
rect 33152 15366 33180 21286
rect 33140 15360 33192 15366
rect 33140 15302 33192 15308
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33060 14414 33088 15098
rect 33152 15026 33180 15302
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33140 14816 33192 14822
rect 33140 14758 33192 14764
rect 33152 14414 33180 14758
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 33060 12918 33088 14350
rect 33244 14074 33272 21406
rect 33428 19786 33456 21406
rect 33416 19780 33468 19786
rect 33416 19722 33468 19728
rect 33414 17912 33470 17921
rect 33414 17847 33470 17856
rect 33428 17678 33456 17847
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33520 17202 33548 23462
rect 33612 22030 33640 33798
rect 33704 31822 33732 33918
rect 33782 33895 33838 33904
rect 33782 33824 33838 33833
rect 33782 33759 33838 33768
rect 33692 31816 33744 31822
rect 33692 31758 33744 31764
rect 33704 30734 33732 31758
rect 33796 30870 33824 33759
rect 33784 30864 33836 30870
rect 33784 30806 33836 30812
rect 33692 30728 33744 30734
rect 33692 30670 33744 30676
rect 33888 27538 33916 34439
rect 34152 34410 34204 34416
rect 34244 34468 34296 34474
rect 34244 34410 34296 34416
rect 34164 33998 34192 34410
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 34152 33992 34204 33998
rect 34152 33934 34204 33940
rect 33980 32978 34008 33934
rect 34348 33538 34376 35550
rect 34440 34746 34468 36774
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34428 34740 34480 34746
rect 34428 34682 34480 34688
rect 34428 34604 34480 34610
rect 34428 34546 34480 34552
rect 34440 33930 34468 34546
rect 34532 34134 34560 35974
rect 34520 34128 34572 34134
rect 34520 34070 34572 34076
rect 34428 33924 34480 33930
rect 34428 33866 34480 33872
rect 34256 33510 34376 33538
rect 33968 32972 34020 32978
rect 33968 32914 34020 32920
rect 34150 31512 34206 31521
rect 34150 31447 34152 31456
rect 34204 31447 34206 31456
rect 34152 31418 34204 31424
rect 34256 31346 34284 33510
rect 34440 33402 34468 33866
rect 34520 33856 34572 33862
rect 34520 33798 34572 33804
rect 34348 33374 34468 33402
rect 34348 32774 34376 33374
rect 34428 33312 34480 33318
rect 34428 33254 34480 33260
rect 34440 32910 34468 33254
rect 34428 32904 34480 32910
rect 34428 32846 34480 32852
rect 34336 32768 34388 32774
rect 34532 32722 34560 33798
rect 34336 32710 34388 32716
rect 34348 32570 34376 32710
rect 34440 32694 34560 32722
rect 34336 32564 34388 32570
rect 34336 32506 34388 32512
rect 34440 32434 34468 32694
rect 34520 32496 34572 32502
rect 34624 32484 34652 39782
rect 34716 39302 34744 40122
rect 34704 39296 34756 39302
rect 34704 39238 34756 39244
rect 34716 38826 34744 39238
rect 34808 38962 34836 40462
rect 34992 39846 35020 40462
rect 34980 39840 35032 39846
rect 34980 39782 35032 39788
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34888 39636 34940 39642
rect 34888 39578 34940 39584
rect 34900 39438 34928 39578
rect 34888 39432 34940 39438
rect 34888 39374 34940 39380
rect 34796 38956 34848 38962
rect 34796 38898 34848 38904
rect 34704 38820 34756 38826
rect 34704 38762 34756 38768
rect 34572 32456 34652 32484
rect 34520 32438 34572 32444
rect 34428 32428 34480 32434
rect 34428 32370 34480 32376
rect 34612 32224 34664 32230
rect 34612 32166 34664 32172
rect 34336 31476 34388 31482
rect 34336 31418 34388 31424
rect 34244 31340 34296 31346
rect 34244 31282 34296 31288
rect 34348 31142 34376 31418
rect 34428 31408 34480 31414
rect 34428 31350 34480 31356
rect 34336 31136 34388 31142
rect 34336 31078 34388 31084
rect 34244 30728 34296 30734
rect 34244 30670 34296 30676
rect 33968 30660 34020 30666
rect 33968 30602 34020 30608
rect 33980 29850 34008 30602
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 33968 29844 34020 29850
rect 33968 29786 34020 29792
rect 34072 29560 34100 30194
rect 34152 29572 34204 29578
rect 34072 29532 34152 29560
rect 34152 29514 34204 29520
rect 33968 29096 34020 29102
rect 33968 29038 34020 29044
rect 33980 27606 34008 29038
rect 34164 28626 34192 29514
rect 34152 28620 34204 28626
rect 34152 28562 34204 28568
rect 33968 27600 34020 27606
rect 33968 27542 34020 27548
rect 33876 27532 33928 27538
rect 33876 27474 33928 27480
rect 33784 26852 33836 26858
rect 33784 26794 33836 26800
rect 33796 26382 33824 26794
rect 33980 26382 34008 27542
rect 34164 27112 34192 28562
rect 34256 28490 34284 30670
rect 34336 30048 34388 30054
rect 34336 29990 34388 29996
rect 34348 28558 34376 29990
rect 34440 29170 34468 31350
rect 34520 31136 34572 31142
rect 34520 31078 34572 31084
rect 34532 30433 34560 31078
rect 34518 30424 34574 30433
rect 34518 30359 34574 30368
rect 34520 30184 34572 30190
rect 34520 30126 34572 30132
rect 34532 29850 34560 30126
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34532 29646 34560 29786
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34532 29306 34560 29582
rect 34520 29300 34572 29306
rect 34520 29242 34572 29248
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34624 29050 34652 32166
rect 34716 31346 34744 38762
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35072 38344 35124 38350
rect 35072 38286 35124 38292
rect 34796 38208 34848 38214
rect 34796 38150 34848 38156
rect 34808 36854 34836 38150
rect 35084 37874 35112 38286
rect 35072 37868 35124 37874
rect 35072 37810 35124 37816
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37330 35480 41006
rect 35636 40458 35664 41142
rect 35912 40526 35940 41414
rect 38028 41274 38056 41482
rect 38016 41268 38068 41274
rect 38016 41210 38068 41216
rect 38384 41200 38436 41206
rect 38384 41142 38436 41148
rect 37556 41064 37608 41070
rect 37556 41006 37608 41012
rect 36912 40928 36964 40934
rect 36912 40870 36964 40876
rect 36924 40730 36952 40870
rect 36912 40724 36964 40730
rect 36912 40666 36964 40672
rect 35900 40520 35952 40526
rect 35900 40462 35952 40468
rect 35624 40452 35676 40458
rect 35624 40394 35676 40400
rect 36452 39908 36504 39914
rect 36452 39850 36504 39856
rect 36084 39364 36136 39370
rect 36084 39306 36136 39312
rect 36096 38894 36124 39306
rect 36464 38962 36492 39850
rect 36636 39500 36688 39506
rect 36636 39442 36688 39448
rect 37004 39500 37056 39506
rect 37004 39442 37056 39448
rect 36544 39024 36596 39030
rect 36648 39012 36676 39442
rect 36910 39400 36966 39409
rect 36910 39335 36966 39344
rect 36728 39092 36780 39098
rect 36728 39034 36780 39040
rect 36596 38984 36676 39012
rect 36544 38966 36596 38972
rect 36268 38956 36320 38962
rect 36268 38898 36320 38904
rect 36452 38956 36504 38962
rect 36452 38898 36504 38904
rect 36084 38888 36136 38894
rect 36084 38830 36136 38836
rect 35532 38752 35584 38758
rect 35530 38720 35532 38729
rect 35584 38720 35586 38729
rect 35530 38655 35586 38664
rect 36096 38350 36124 38830
rect 36176 38412 36228 38418
rect 36176 38354 36228 38360
rect 36084 38344 36136 38350
rect 36084 38286 36136 38292
rect 35992 38208 36044 38214
rect 35992 38150 36044 38156
rect 35900 37868 35952 37874
rect 35900 37810 35952 37816
rect 35808 37392 35860 37398
rect 35912 37369 35940 37810
rect 36004 37806 36032 38150
rect 36096 38010 36124 38286
rect 36188 38010 36216 38354
rect 36280 38010 36308 38898
rect 36464 38842 36492 38898
rect 36464 38814 36584 38842
rect 36740 38826 36768 39034
rect 36924 38894 36952 39335
rect 36912 38888 36964 38894
rect 36912 38830 36964 38836
rect 36360 38344 36412 38350
rect 36360 38286 36412 38292
rect 36084 38004 36136 38010
rect 36084 37946 36136 37952
rect 36176 38004 36228 38010
rect 36176 37946 36228 37952
rect 36268 38004 36320 38010
rect 36268 37946 36320 37952
rect 35992 37800 36044 37806
rect 35992 37742 36044 37748
rect 35808 37334 35860 37340
rect 35898 37360 35954 37369
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35532 37188 35584 37194
rect 35532 37130 35584 37136
rect 34796 36848 34848 36854
rect 34796 36790 34848 36796
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 34808 36242 34836 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35070 36272 35126 36281
rect 34796 36236 34848 36242
rect 35070 36207 35126 36216
rect 34796 36178 34848 36184
rect 35084 36174 35112 36207
rect 35072 36168 35124 36174
rect 35072 36110 35124 36116
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34888 35284 34940 35290
rect 34888 35226 34940 35232
rect 34900 34542 34928 35226
rect 35348 34944 35400 34950
rect 35348 34886 35400 34892
rect 34888 34536 34940 34542
rect 34888 34478 34940 34484
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35256 33924 35308 33930
rect 35360 33912 35388 34886
rect 35440 34060 35492 34066
rect 35440 34002 35492 34008
rect 35308 33884 35388 33912
rect 35256 33866 35308 33872
rect 34796 33584 34848 33590
rect 34796 33526 34848 33532
rect 34808 32230 34836 33526
rect 35348 33312 35400 33318
rect 35348 33254 35400 33260
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 32978 35388 33254
rect 35256 32972 35308 32978
rect 35256 32914 35308 32920
rect 35348 32972 35400 32978
rect 35348 32914 35400 32920
rect 35268 32858 35296 32914
rect 34980 32836 35032 32842
rect 35268 32830 35388 32858
rect 34980 32778 35032 32784
rect 34992 32434 35020 32778
rect 34980 32428 35032 32434
rect 34980 32370 35032 32376
rect 35256 32428 35308 32434
rect 35256 32370 35308 32376
rect 35268 32337 35296 32370
rect 35254 32328 35310 32337
rect 35254 32263 35310 32272
rect 34796 32224 34848 32230
rect 34796 32166 34848 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35256 32020 35308 32026
rect 35256 31962 35308 31968
rect 34796 31952 34848 31958
rect 35268 31929 35296 31962
rect 34796 31894 34848 31900
rect 35254 31920 35310 31929
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34808 30240 34836 31894
rect 35254 31855 35310 31864
rect 35164 31816 35216 31822
rect 35162 31784 35164 31793
rect 35216 31784 35218 31793
rect 35162 31719 35218 31728
rect 35268 31090 35296 31855
rect 35360 31210 35388 32830
rect 35452 31958 35480 34002
rect 35544 33590 35572 37130
rect 35728 36310 35756 37198
rect 35716 36304 35768 36310
rect 35716 36246 35768 36252
rect 35624 35624 35676 35630
rect 35624 35566 35676 35572
rect 35532 33584 35584 33590
rect 35532 33526 35584 33532
rect 35532 33040 35584 33046
rect 35532 32982 35584 32988
rect 35440 31952 35492 31958
rect 35440 31894 35492 31900
rect 35440 31272 35492 31278
rect 35438 31240 35440 31249
rect 35492 31240 35494 31249
rect 35348 31204 35400 31210
rect 35438 31175 35494 31184
rect 35348 31146 35400 31152
rect 35268 31062 35388 31090
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34980 30728 35032 30734
rect 34980 30670 35032 30676
rect 35164 30728 35216 30734
rect 35164 30670 35216 30676
rect 34716 30212 34836 30240
rect 34888 30252 34940 30258
rect 34716 29209 34744 30212
rect 34888 30194 34940 30200
rect 34900 30161 34928 30194
rect 34886 30152 34942 30161
rect 34796 30116 34848 30122
rect 34992 30122 35020 30670
rect 35176 30326 35204 30670
rect 35164 30320 35216 30326
rect 35164 30262 35216 30268
rect 34886 30087 34942 30096
rect 34980 30116 35032 30122
rect 34796 30058 34848 30064
rect 34980 30058 35032 30064
rect 34808 29628 34836 30058
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34980 29640 35032 29646
rect 34808 29600 34980 29628
rect 34980 29582 35032 29588
rect 34702 29200 34758 29209
rect 34796 29164 34848 29170
rect 34758 29144 34796 29152
rect 34702 29135 34796 29144
rect 34716 29124 34796 29135
rect 34796 29106 34848 29112
rect 34532 29022 34652 29050
rect 34796 29028 34848 29034
rect 34336 28552 34388 28558
rect 34336 28494 34388 28500
rect 34244 28484 34296 28490
rect 34244 28426 34296 28432
rect 34348 28082 34376 28494
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 34440 28014 34468 28426
rect 34428 28008 34480 28014
rect 34428 27950 34480 27956
rect 34164 27084 34284 27112
rect 34256 26994 34284 27084
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33980 23730 34008 26318
rect 34060 26308 34112 26314
rect 34060 26250 34112 26256
rect 34072 25702 34100 26250
rect 34164 25945 34192 26930
rect 34244 26512 34296 26518
rect 34244 26454 34296 26460
rect 34256 26382 34284 26454
rect 34440 26382 34468 27950
rect 34532 27674 34560 29022
rect 34796 28970 34848 28976
rect 34612 28416 34664 28422
rect 34612 28358 34664 28364
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34624 26586 34652 28358
rect 34808 27538 34836 28970
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35072 28552 35124 28558
rect 35072 28494 35124 28500
rect 35084 28082 35112 28494
rect 35256 28484 35308 28490
rect 35256 28426 35308 28432
rect 35268 28218 35296 28426
rect 35256 28212 35308 28218
rect 35256 28154 35308 28160
rect 35072 28076 35124 28082
rect 35072 28018 35124 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 34980 27464 35032 27470
rect 34980 27406 35032 27412
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34612 26580 34664 26586
rect 34612 26522 34664 26528
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 34518 26344 34574 26353
rect 34150 25936 34206 25945
rect 34150 25871 34206 25880
rect 34060 25696 34112 25702
rect 34060 25638 34112 25644
rect 34256 25362 34284 26318
rect 34518 26279 34574 26288
rect 34426 25936 34482 25945
rect 34426 25871 34428 25880
rect 34480 25871 34482 25880
rect 34428 25842 34480 25848
rect 34244 25356 34296 25362
rect 34244 25298 34296 25304
rect 34058 23760 34114 23769
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33968 23724 34020 23730
rect 34058 23695 34060 23704
rect 33968 23666 34020 23672
rect 34112 23695 34114 23704
rect 34060 23666 34112 23672
rect 33704 23118 33732 23666
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 33692 23112 33744 23118
rect 33744 23060 33824 23066
rect 33692 23054 33824 23060
rect 33704 23038 33824 23054
rect 33692 22704 33744 22710
rect 33692 22646 33744 22652
rect 33600 22024 33652 22030
rect 33600 21966 33652 21972
rect 33612 21486 33640 21966
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33600 21004 33652 21010
rect 33600 20946 33652 20952
rect 33612 17202 33640 20946
rect 33704 20942 33732 22646
rect 33796 22642 33824 23038
rect 33784 22636 33836 22642
rect 33784 22578 33836 22584
rect 34072 22094 34100 23462
rect 34256 23118 34284 25298
rect 34428 24268 34480 24274
rect 34428 24210 34480 24216
rect 34244 23112 34296 23118
rect 34244 23054 34296 23060
rect 34152 23044 34204 23050
rect 34152 22986 34204 22992
rect 34164 22506 34192 22986
rect 34256 22642 34284 23054
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34152 22500 34204 22506
rect 34152 22442 34204 22448
rect 34244 22500 34296 22506
rect 34244 22442 34296 22448
rect 34072 22066 34192 22094
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 33784 21888 33836 21894
rect 33784 21830 33836 21836
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33704 20398 33732 20878
rect 33692 20392 33744 20398
rect 33692 20334 33744 20340
rect 33704 20058 33732 20334
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 33692 19712 33744 19718
rect 33692 19654 33744 19660
rect 33704 18766 33732 19654
rect 33796 18970 33824 21830
rect 33968 21616 34020 21622
rect 34072 21604 34100 21898
rect 34020 21576 34100 21604
rect 33968 21558 34020 21564
rect 33876 20868 33928 20874
rect 33876 20810 33928 20816
rect 33888 19854 33916 20810
rect 34072 20602 34100 21576
rect 34164 21554 34192 22066
rect 34256 21962 34284 22442
rect 34244 21956 34296 21962
rect 34244 21898 34296 21904
rect 34336 21956 34388 21962
rect 34336 21898 34388 21904
rect 34152 21548 34204 21554
rect 34152 21490 34204 21496
rect 34164 20942 34192 21490
rect 34348 21418 34376 21898
rect 34440 21894 34468 24210
rect 34532 22642 34560 26279
rect 34612 24132 34664 24138
rect 34612 24074 34664 24080
rect 34624 23730 34652 24074
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34624 23526 34652 23666
rect 34612 23520 34664 23526
rect 34612 23462 34664 23468
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 34428 21888 34480 21894
rect 34428 21830 34480 21836
rect 34244 21412 34296 21418
rect 34244 21354 34296 21360
rect 34336 21412 34388 21418
rect 34336 21354 34388 21360
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34072 19854 34100 20538
rect 34256 20466 34284 21354
rect 34440 21010 34468 21830
rect 34532 21486 34560 22578
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 34334 20632 34390 20641
rect 34334 20567 34390 20576
rect 34244 20460 34296 20466
rect 34244 20402 34296 20408
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 34060 19848 34112 19854
rect 34060 19790 34112 19796
rect 34256 19378 34284 20402
rect 34348 19854 34376 20567
rect 34532 20466 34560 21286
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34336 19848 34388 19854
rect 34336 19790 34388 19796
rect 34428 19780 34480 19786
rect 34428 19722 34480 19728
rect 34440 19514 34468 19722
rect 34428 19508 34480 19514
rect 34428 19450 34480 19456
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 33784 18964 33836 18970
rect 33784 18906 33836 18912
rect 33692 18760 33744 18766
rect 33692 18702 33744 18708
rect 33704 18154 33732 18702
rect 33796 18290 33824 18906
rect 33784 18284 33836 18290
rect 33784 18226 33836 18232
rect 33692 18148 33744 18154
rect 33692 18090 33744 18096
rect 33876 17808 33928 17814
rect 33876 17750 33928 17756
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33692 16992 33744 16998
rect 33692 16934 33744 16940
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33336 14890 33364 16050
rect 33324 14884 33376 14890
rect 33324 14826 33376 14832
rect 33416 14884 33468 14890
rect 33416 14826 33468 14832
rect 33428 14770 33456 14826
rect 33336 14742 33456 14770
rect 33336 14618 33364 14742
rect 33324 14612 33376 14618
rect 33324 14554 33376 14560
rect 33232 14068 33284 14074
rect 33232 14010 33284 14016
rect 33336 13870 33364 14554
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 33048 12912 33100 12918
rect 33048 12854 33100 12860
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 32784 12442 32812 12786
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 33336 12374 33364 13806
rect 33324 12368 33376 12374
rect 33324 12310 33376 12316
rect 32588 12300 32640 12306
rect 32588 12242 32640 12248
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32864 11076 32916 11082
rect 32864 11018 32916 11024
rect 32876 10810 32904 11018
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 32864 10804 32916 10810
rect 32864 10746 32916 10752
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 31220 10062 31248 10746
rect 33336 10606 33364 12310
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 33704 6798 33732 16934
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33796 14006 33824 14554
rect 33784 14000 33836 14006
rect 33784 13942 33836 13948
rect 33888 13818 33916 17750
rect 34520 16584 34572 16590
rect 34520 16526 34572 16532
rect 34428 15904 34480 15910
rect 34428 15846 34480 15852
rect 34440 15502 34468 15846
rect 34532 15706 34560 16526
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 34428 15496 34480 15502
rect 34428 15438 34480 15444
rect 33968 15428 34020 15434
rect 33968 15370 34020 15376
rect 33980 13938 34008 15370
rect 34440 15094 34468 15438
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34428 14340 34480 14346
rect 34428 14282 34480 14288
rect 34440 14074 34468 14282
rect 34532 14074 34560 14962
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 33796 13790 33916 13818
rect 33796 8498 33824 13790
rect 33980 13394 34008 13874
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33980 12850 34008 13330
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33888 12238 33916 12582
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 34164 11914 34192 12786
rect 34072 11886 34192 11914
rect 34072 11830 34100 11886
rect 34060 11824 34112 11830
rect 34060 11766 34112 11772
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 33980 11354 34008 11698
rect 33968 11348 34020 11354
rect 33968 11290 34020 11296
rect 33980 10810 34008 11290
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 34624 6914 34652 22918
rect 34716 21690 34744 27270
rect 34992 27130 35020 27406
rect 34980 27124 35032 27130
rect 34980 27066 35032 27072
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 34808 25906 34836 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35164 26376 35216 26382
rect 35164 26318 35216 26324
rect 35176 26246 35204 26318
rect 35164 26240 35216 26246
rect 35164 26182 35216 26188
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24206 35388 31062
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 35452 28558 35480 30194
rect 35544 30122 35572 32982
rect 35532 30116 35584 30122
rect 35532 30058 35584 30064
rect 35532 29844 35584 29850
rect 35532 29786 35584 29792
rect 35544 28994 35572 29786
rect 35636 29238 35664 35566
rect 35820 35290 35848 37334
rect 35898 37295 35954 37304
rect 36096 36174 36124 37946
rect 36188 37890 36216 37946
rect 36188 37862 36308 37890
rect 36176 36236 36228 36242
rect 36176 36178 36228 36184
rect 36084 36168 36136 36174
rect 36084 36110 36136 36116
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35808 35284 35860 35290
rect 35808 35226 35860 35232
rect 35808 35080 35860 35086
rect 35900 35080 35952 35086
rect 35808 35022 35860 35028
rect 35898 35048 35900 35057
rect 35952 35048 35954 35057
rect 35716 35012 35768 35018
rect 35716 34954 35768 34960
rect 35728 33998 35756 34954
rect 35820 34746 35848 35022
rect 35898 34983 35954 34992
rect 35808 34740 35860 34746
rect 35808 34682 35860 34688
rect 35912 34678 35940 34983
rect 35900 34672 35952 34678
rect 35900 34614 35952 34620
rect 36004 34610 36032 35974
rect 36188 35766 36216 36178
rect 36176 35760 36228 35766
rect 36176 35702 36228 35708
rect 36084 35216 36136 35222
rect 36084 35158 36136 35164
rect 36096 35018 36124 35158
rect 36084 35012 36136 35018
rect 36084 34954 36136 34960
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 35808 34400 35860 34406
rect 35808 34342 35860 34348
rect 35716 33992 35768 33998
rect 35716 33934 35768 33940
rect 35820 33862 35848 34342
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 35716 33856 35768 33862
rect 35716 33798 35768 33804
rect 35808 33856 35860 33862
rect 35808 33798 35860 33804
rect 35728 32910 35756 33798
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35728 32230 35756 32846
rect 35716 32224 35768 32230
rect 35716 32166 35768 32172
rect 35716 31952 35768 31958
rect 35714 31920 35716 31929
rect 35768 31920 35770 31929
rect 35714 31855 35770 31864
rect 35820 31804 35848 33798
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 35912 32026 35940 32846
rect 36004 32434 36032 34138
rect 36096 32774 36124 34954
rect 36188 34649 36216 34954
rect 36174 34640 36230 34649
rect 36174 34575 36230 34584
rect 36176 34468 36228 34474
rect 36176 34410 36228 34416
rect 36188 33833 36216 34410
rect 36174 33824 36230 33833
rect 36174 33759 36230 33768
rect 36188 33590 36216 33759
rect 36176 33584 36228 33590
rect 36176 33526 36228 33532
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 36084 32768 36136 32774
rect 36084 32710 36136 32716
rect 35992 32428 36044 32434
rect 35992 32370 36044 32376
rect 35900 32020 35952 32026
rect 35900 31962 35952 31968
rect 36004 31822 36032 32370
rect 36084 32020 36136 32026
rect 36084 31962 36136 31968
rect 35728 31776 35848 31804
rect 35992 31816 36044 31822
rect 35990 31784 35992 31793
rect 36044 31784 36046 31793
rect 35728 30394 35756 31776
rect 35990 31719 36046 31728
rect 35900 31680 35952 31686
rect 35900 31622 35952 31628
rect 35992 31680 36044 31686
rect 35992 31622 36044 31628
rect 35912 31210 35940 31622
rect 36004 31346 36032 31622
rect 36096 31414 36124 31962
rect 36084 31408 36136 31414
rect 36084 31350 36136 31356
rect 35992 31340 36044 31346
rect 35992 31282 36044 31288
rect 35808 31204 35860 31210
rect 35808 31146 35860 31152
rect 35900 31204 35952 31210
rect 35900 31146 35952 31152
rect 35820 30410 35848 31146
rect 36084 31136 36136 31142
rect 36084 31078 36136 31084
rect 36096 30734 36124 31078
rect 36188 30818 36216 32846
rect 36280 30938 36308 37862
rect 36372 37738 36400 38286
rect 36452 37868 36504 37874
rect 36452 37810 36504 37816
rect 36360 37732 36412 37738
rect 36360 37674 36412 37680
rect 36464 37466 36492 37810
rect 36452 37460 36504 37466
rect 36452 37402 36504 37408
rect 36360 36100 36412 36106
rect 36360 36042 36412 36048
rect 36372 34610 36400 36042
rect 36464 36038 36492 37402
rect 36452 36032 36504 36038
rect 36452 35974 36504 35980
rect 36452 35080 36504 35086
rect 36450 35048 36452 35057
rect 36504 35048 36506 35057
rect 36450 34983 36506 34992
rect 36360 34604 36412 34610
rect 36360 34546 36412 34552
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 36372 32570 36400 34546
rect 36464 33658 36492 34546
rect 36452 33652 36504 33658
rect 36452 33594 36504 33600
rect 36464 33318 36492 33594
rect 36452 33312 36504 33318
rect 36452 33254 36504 33260
rect 36452 32836 36504 32842
rect 36452 32778 36504 32784
rect 36360 32564 36412 32570
rect 36360 32506 36412 32512
rect 36372 31890 36400 32506
rect 36360 31884 36412 31890
rect 36360 31826 36412 31832
rect 36464 31346 36492 32778
rect 36556 32026 36584 38814
rect 36728 38820 36780 38826
rect 36728 38762 36780 38768
rect 36728 38344 36780 38350
rect 36728 38286 36780 38292
rect 36740 37874 36768 38286
rect 37016 38282 37044 39442
rect 37096 39432 37148 39438
rect 37096 39374 37148 39380
rect 37188 39432 37240 39438
rect 37188 39374 37240 39380
rect 37108 38554 37136 39374
rect 37200 39273 37228 39374
rect 37280 39296 37332 39302
rect 37186 39264 37242 39273
rect 37280 39238 37332 39244
rect 37186 39199 37242 39208
rect 37200 38758 37228 39199
rect 37188 38752 37240 38758
rect 37188 38694 37240 38700
rect 37096 38548 37148 38554
rect 37096 38490 37148 38496
rect 36820 38276 36872 38282
rect 36820 38218 36872 38224
rect 37004 38276 37056 38282
rect 37004 38218 37056 38224
rect 36728 37868 36780 37874
rect 36728 37810 36780 37816
rect 36832 37176 36860 38218
rect 36912 38208 36964 38214
rect 36912 38150 36964 38156
rect 36924 37369 36952 38150
rect 37292 37874 37320 39238
rect 37568 39098 37596 41006
rect 38396 40526 38424 41142
rect 38568 41132 38620 41138
rect 38568 41074 38620 41080
rect 38476 41064 38528 41070
rect 38476 41006 38528 41012
rect 38488 40730 38516 41006
rect 38476 40724 38528 40730
rect 38476 40666 38528 40672
rect 38580 40526 38608 41074
rect 38384 40520 38436 40526
rect 38384 40462 38436 40468
rect 38568 40520 38620 40526
rect 38568 40462 38620 40468
rect 38844 40520 38896 40526
rect 38844 40462 38896 40468
rect 38396 39642 38424 40462
rect 38580 39846 38608 40462
rect 38856 40118 38884 40462
rect 38660 40112 38712 40118
rect 38660 40054 38712 40060
rect 38844 40112 38896 40118
rect 38844 40054 38896 40060
rect 38568 39840 38620 39846
rect 38568 39782 38620 39788
rect 38384 39636 38436 39642
rect 38384 39578 38436 39584
rect 37740 39500 37792 39506
rect 37660 39460 37740 39488
rect 37556 39092 37608 39098
rect 37556 39034 37608 39040
rect 37660 38962 37688 39460
rect 37740 39442 37792 39448
rect 37924 39432 37976 39438
rect 37924 39374 37976 39380
rect 37936 39098 37964 39374
rect 37924 39092 37976 39098
rect 37924 39034 37976 39040
rect 37740 39024 37792 39030
rect 37792 38984 37872 39012
rect 37740 38966 37792 38972
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 37648 38956 37700 38962
rect 37648 38898 37700 38904
rect 37280 37868 37332 37874
rect 37280 37810 37332 37816
rect 37188 37460 37240 37466
rect 37188 37402 37240 37408
rect 36910 37360 36966 37369
rect 36910 37295 36966 37304
rect 37200 37262 37228 37402
rect 37188 37256 37240 37262
rect 37188 37198 37240 37204
rect 36912 37188 36964 37194
rect 36832 37148 36912 37176
rect 37280 37188 37332 37194
rect 36964 37148 37044 37176
rect 36912 37130 36964 37136
rect 36636 37120 36688 37126
rect 36636 37062 36688 37068
rect 36648 36922 36676 37062
rect 36636 36916 36688 36922
rect 36636 36858 36688 36864
rect 36820 36712 36872 36718
rect 36820 36654 36872 36660
rect 36636 36168 36688 36174
rect 36636 36110 36688 36116
rect 36648 34610 36676 36110
rect 36728 35148 36780 35154
rect 36728 35090 36780 35096
rect 36740 34746 36768 35090
rect 36728 34740 36780 34746
rect 36728 34682 36780 34688
rect 36636 34604 36688 34610
rect 36636 34546 36688 34552
rect 36648 34202 36676 34546
rect 36636 34196 36688 34202
rect 36636 34138 36688 34144
rect 36728 33448 36780 33454
rect 36728 33390 36780 33396
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 36544 32020 36596 32026
rect 36544 31962 36596 31968
rect 36648 31958 36676 32302
rect 36636 31952 36688 31958
rect 36636 31894 36688 31900
rect 36648 31754 36676 31894
rect 36636 31748 36688 31754
rect 36636 31690 36688 31696
rect 36452 31340 36504 31346
rect 36452 31282 36504 31288
rect 36544 31340 36596 31346
rect 36544 31282 36596 31288
rect 36268 30932 36320 30938
rect 36268 30874 36320 30880
rect 36556 30870 36584 31282
rect 36636 31204 36688 31210
rect 36636 31146 36688 31152
rect 36544 30864 36596 30870
rect 36188 30790 36400 30818
rect 36544 30806 36596 30812
rect 36372 30734 36400 30790
rect 36084 30728 36136 30734
rect 36084 30670 36136 30676
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 36360 30728 36412 30734
rect 36360 30670 36412 30676
rect 35716 30388 35768 30394
rect 35820 30382 36032 30410
rect 36188 30394 36216 30670
rect 35716 30330 35768 30336
rect 35714 30288 35770 30297
rect 35714 30223 35716 30232
rect 35768 30223 35770 30232
rect 35808 30252 35860 30258
rect 35716 30194 35768 30200
rect 35808 30194 35860 30200
rect 35624 29232 35676 29238
rect 35624 29174 35676 29180
rect 35544 28966 35664 28994
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 35636 28082 35664 28966
rect 35624 28076 35676 28082
rect 35624 28018 35676 28024
rect 35636 27606 35664 28018
rect 35624 27600 35676 27606
rect 35624 27542 35676 27548
rect 35440 27396 35492 27402
rect 35440 27338 35492 27344
rect 35452 25294 35480 27338
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 35544 26246 35572 26522
rect 35532 26240 35584 26246
rect 35636 26228 35664 27542
rect 35728 26353 35756 30194
rect 35820 29714 35848 30194
rect 35900 30184 35952 30190
rect 35900 30126 35952 30132
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 35912 27062 35940 30126
rect 36004 29646 36032 30382
rect 36176 30388 36228 30394
rect 36176 30330 36228 30336
rect 36176 29844 36228 29850
rect 36176 29786 36228 29792
rect 35992 29640 36044 29646
rect 35992 29582 36044 29588
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 36004 28082 36032 29106
rect 36084 28144 36136 28150
rect 36084 28086 36136 28092
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 36004 27674 36032 28018
rect 35992 27668 36044 27674
rect 35992 27610 36044 27616
rect 35900 27056 35952 27062
rect 35900 26998 35952 27004
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35714 26344 35770 26353
rect 35714 26279 35770 26288
rect 35636 26200 35756 26228
rect 35532 26182 35584 26188
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 35268 23594 35296 24006
rect 35360 23730 35388 24142
rect 35544 24138 35572 26182
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 35636 25294 35664 25774
rect 35624 25288 35676 25294
rect 35624 25230 35676 25236
rect 35728 25226 35756 26200
rect 35820 25906 35848 26454
rect 35808 25900 35860 25906
rect 35808 25842 35860 25848
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 35808 25220 35860 25226
rect 35808 25162 35860 25168
rect 35728 24886 35756 25162
rect 35820 24954 35848 25162
rect 35808 24948 35860 24954
rect 35808 24890 35860 24896
rect 35716 24880 35768 24886
rect 35716 24822 35768 24828
rect 35820 24342 35848 24890
rect 35912 24614 35940 26998
rect 36004 26450 36032 27610
rect 36096 27470 36124 28086
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36084 27328 36136 27334
rect 36084 27270 36136 27276
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 35992 25968 36044 25974
rect 35992 25910 36044 25916
rect 36004 24818 36032 25910
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 35900 24608 35952 24614
rect 35900 24550 35952 24556
rect 35808 24336 35860 24342
rect 35808 24278 35860 24284
rect 35532 24132 35584 24138
rect 35532 24074 35584 24080
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35256 23588 35308 23594
rect 35256 23530 35308 23536
rect 35348 23588 35400 23594
rect 35348 23530 35400 23536
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 23338 35388 23530
rect 35268 23310 35388 23338
rect 35268 22710 35296 23310
rect 35544 23186 35572 23666
rect 35912 23662 35940 24550
rect 36004 23798 36032 24754
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 36004 23202 36032 23734
rect 35532 23180 35584 23186
rect 35532 23122 35584 23128
rect 35636 23174 36032 23202
rect 36096 23186 36124 27270
rect 36188 26926 36216 29786
rect 36372 27470 36400 30670
rect 36648 30258 36676 31146
rect 36636 30252 36688 30258
rect 36636 30194 36688 30200
rect 36450 30152 36506 30161
rect 36450 30087 36506 30096
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 36464 26382 36492 30087
rect 36648 29850 36676 30194
rect 36740 30054 36768 33390
rect 36728 30048 36780 30054
rect 36728 29990 36780 29996
rect 36636 29844 36688 29850
rect 36636 29786 36688 29792
rect 36728 29572 36780 29578
rect 36728 29514 36780 29520
rect 36740 29306 36768 29514
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 36634 27568 36690 27577
rect 36634 27503 36690 27512
rect 36542 26888 36598 26897
rect 36542 26823 36598 26832
rect 36452 26376 36504 26382
rect 36452 26318 36504 26324
rect 36176 26308 36228 26314
rect 36176 26250 36228 26256
rect 36188 25498 36216 26250
rect 36556 26246 36584 26823
rect 36648 26382 36676 27503
rect 36728 27396 36780 27402
rect 36728 27338 36780 27344
rect 36740 27062 36768 27338
rect 36728 27056 36780 27062
rect 36728 26998 36780 27004
rect 36740 26382 36768 26998
rect 36832 26858 36860 36654
rect 36912 36168 36964 36174
rect 36912 36110 36964 36116
rect 36924 35834 36952 36110
rect 37016 36106 37044 37148
rect 37280 37130 37332 37136
rect 37292 37074 37320 37130
rect 37200 37046 37320 37074
rect 37004 36100 37056 36106
rect 37004 36042 37056 36048
rect 36912 35828 36964 35834
rect 36912 35770 36964 35776
rect 36924 35562 36952 35770
rect 36912 35556 36964 35562
rect 36912 35498 36964 35504
rect 36912 35080 36964 35086
rect 36912 35022 36964 35028
rect 36924 32570 36952 35022
rect 37094 34504 37150 34513
rect 37094 34439 37150 34448
rect 37108 33658 37136 34439
rect 37096 33652 37148 33658
rect 37096 33594 37148 33600
rect 36912 32564 36964 32570
rect 36912 32506 36964 32512
rect 37096 31884 37148 31890
rect 37096 31826 37148 31832
rect 36912 31816 36964 31822
rect 36912 31758 36964 31764
rect 36924 31142 36952 31758
rect 37108 31754 37136 31826
rect 37096 31748 37148 31754
rect 37096 31690 37148 31696
rect 36912 31136 36964 31142
rect 36912 31078 36964 31084
rect 36924 28966 36952 31078
rect 37004 30932 37056 30938
rect 37004 30874 37056 30880
rect 36912 28960 36964 28966
rect 36912 28902 36964 28908
rect 36912 28756 36964 28762
rect 36912 28698 36964 28704
rect 36924 28558 36952 28698
rect 36912 28552 36964 28558
rect 36912 28494 36964 28500
rect 36924 28422 36952 28494
rect 36912 28416 36964 28422
rect 36912 28358 36964 28364
rect 36912 27940 36964 27946
rect 36912 27882 36964 27888
rect 36924 27033 36952 27882
rect 36910 27024 36966 27033
rect 36910 26959 36966 26968
rect 36924 26926 36952 26959
rect 36912 26920 36964 26926
rect 36912 26862 36964 26868
rect 37016 26858 37044 30874
rect 37096 30048 37148 30054
rect 37096 29990 37148 29996
rect 37108 29646 37136 29990
rect 37096 29640 37148 29646
rect 37096 29582 37148 29588
rect 37108 28150 37136 29582
rect 37096 28144 37148 28150
rect 37096 28086 37148 28092
rect 37096 27668 37148 27674
rect 37096 27610 37148 27616
rect 37108 27470 37136 27610
rect 37096 27464 37148 27470
rect 37096 27406 37148 27412
rect 37108 27062 37136 27406
rect 37096 27056 37148 27062
rect 37096 26998 37148 27004
rect 36820 26852 36872 26858
rect 36820 26794 36872 26800
rect 37004 26852 37056 26858
rect 37004 26794 37056 26800
rect 36636 26376 36688 26382
rect 36636 26318 36688 26324
rect 36728 26376 36780 26382
rect 36728 26318 36780 26324
rect 36268 26240 36320 26246
rect 36268 26182 36320 26188
rect 36452 26240 36504 26246
rect 36452 26182 36504 26188
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36280 25770 36308 26182
rect 36464 26042 36492 26182
rect 36556 26042 36584 26182
rect 36452 26036 36504 26042
rect 36452 25978 36504 25984
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 36268 25764 36320 25770
rect 36268 25706 36320 25712
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 36556 25378 36584 25978
rect 36832 25786 36860 26794
rect 37200 26586 37228 37046
rect 37384 36378 37412 38898
rect 37844 38654 37872 38984
rect 37936 38962 37964 39034
rect 38580 38962 38608 39782
rect 38672 39370 38700 40054
rect 38856 39370 38884 40054
rect 38936 39840 38988 39846
rect 38936 39782 38988 39788
rect 38948 39438 38976 39782
rect 38936 39432 38988 39438
rect 38936 39374 38988 39380
rect 38660 39364 38712 39370
rect 38660 39306 38712 39312
rect 38844 39364 38896 39370
rect 38844 39306 38896 39312
rect 37924 38956 37976 38962
rect 37924 38898 37976 38904
rect 38568 38956 38620 38962
rect 38568 38898 38620 38904
rect 37752 38626 37872 38654
rect 37464 38344 37516 38350
rect 37464 38286 37516 38292
rect 37648 38344 37700 38350
rect 37648 38286 37700 38292
rect 37476 37466 37504 38286
rect 37464 37460 37516 37466
rect 37464 37402 37516 37408
rect 37660 37398 37688 38286
rect 37752 38282 37780 38626
rect 37936 38350 37964 38898
rect 38672 38554 38700 39306
rect 38660 38548 38712 38554
rect 38660 38490 38712 38496
rect 37924 38344 37976 38350
rect 37844 38304 37924 38332
rect 37740 38276 37792 38282
rect 37740 38218 37792 38224
rect 37648 37392 37700 37398
rect 37648 37334 37700 37340
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 37372 35080 37424 35086
rect 37370 35048 37372 35057
rect 37424 35048 37426 35057
rect 37280 35012 37332 35018
rect 37370 34983 37426 34992
rect 37280 34954 37332 34960
rect 37292 31346 37320 34954
rect 37384 33046 37412 34983
rect 37556 33924 37608 33930
rect 37556 33866 37608 33872
rect 37372 33040 37424 33046
rect 37372 32982 37424 32988
rect 37384 32910 37412 32982
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 37464 32904 37516 32910
rect 37464 32846 37516 32852
rect 37476 32026 37504 32846
rect 37464 32020 37516 32026
rect 37464 31962 37516 31968
rect 37568 31822 37596 33866
rect 37556 31816 37608 31822
rect 37556 31758 37608 31764
rect 37464 31748 37516 31754
rect 37464 31690 37516 31696
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 37292 30569 37320 31282
rect 37476 30841 37504 31690
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37462 30832 37518 30841
rect 37462 30767 37464 30776
rect 37516 30767 37518 30776
rect 37464 30738 37516 30744
rect 37568 30734 37596 30874
rect 37556 30728 37608 30734
rect 37556 30670 37608 30676
rect 37278 30560 37334 30569
rect 37278 30495 37334 30504
rect 37280 30184 37332 30190
rect 37280 30126 37332 30132
rect 37292 29170 37320 30126
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37556 30048 37608 30054
rect 37556 29990 37608 29996
rect 37476 29578 37504 29990
rect 37568 29753 37596 29990
rect 37554 29744 37610 29753
rect 37554 29679 37610 29688
rect 37464 29572 37516 29578
rect 37464 29514 37516 29520
rect 37372 29300 37424 29306
rect 37660 29288 37688 37334
rect 37752 35154 37780 38218
rect 37844 36582 37872 38304
rect 37924 38286 37976 38292
rect 38660 38276 38712 38282
rect 38660 38218 38712 38224
rect 38292 37800 38344 37806
rect 38292 37742 38344 37748
rect 38304 37330 38332 37742
rect 38672 37330 38700 38218
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 38660 37324 38712 37330
rect 38660 37266 38712 37272
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 37740 35148 37792 35154
rect 37740 35090 37792 35096
rect 37844 35086 37872 36518
rect 38016 36168 38068 36174
rect 38068 36128 38148 36156
rect 38016 36110 38068 36116
rect 37924 36032 37976 36038
rect 37924 35974 37976 35980
rect 38016 36032 38068 36038
rect 38016 35974 38068 35980
rect 37936 35766 37964 35974
rect 38028 35766 38056 35974
rect 37924 35760 37976 35766
rect 37924 35702 37976 35708
rect 38016 35760 38068 35766
rect 38016 35702 38068 35708
rect 38028 35290 38056 35702
rect 38120 35494 38148 36128
rect 38108 35488 38160 35494
rect 38108 35430 38160 35436
rect 38016 35284 38068 35290
rect 38016 35226 38068 35232
rect 38120 35222 38148 35430
rect 38108 35216 38160 35222
rect 38108 35158 38160 35164
rect 37832 35080 37884 35086
rect 37832 35022 37884 35028
rect 38200 34536 38252 34542
rect 38200 34478 38252 34484
rect 37740 33516 37792 33522
rect 37740 33458 37792 33464
rect 37752 32366 37780 33458
rect 38028 32978 38148 32994
rect 38016 32972 38148 32978
rect 38068 32966 38148 32972
rect 38016 32914 38068 32920
rect 38016 32836 38068 32842
rect 38016 32778 38068 32784
rect 37832 32768 37884 32774
rect 37832 32710 37884 32716
rect 37844 32366 37872 32710
rect 37924 32496 37976 32502
rect 37924 32438 37976 32444
rect 37740 32360 37792 32366
rect 37740 32302 37792 32308
rect 37832 32360 37884 32366
rect 37832 32302 37884 32308
rect 37740 32224 37792 32230
rect 37740 32166 37792 32172
rect 37372 29242 37424 29248
rect 37476 29260 37688 29288
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37384 28966 37412 29242
rect 37372 28960 37424 28966
rect 37372 28902 37424 28908
rect 37384 28558 37412 28902
rect 37372 28552 37424 28558
rect 37372 28494 37424 28500
rect 37372 28416 37424 28422
rect 37372 28358 37424 28364
rect 37188 26580 37240 26586
rect 37188 26522 37240 26528
rect 37004 26376 37056 26382
rect 37004 26318 37056 26324
rect 37016 25906 37044 26318
rect 37004 25900 37056 25906
rect 37004 25842 37056 25848
rect 36832 25758 36952 25786
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 36372 25350 36584 25378
rect 36268 24676 36320 24682
rect 36268 24618 36320 24624
rect 35636 23118 35664 23174
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 35808 23112 35860 23118
rect 35808 23054 35860 23060
rect 35820 22778 35848 23054
rect 35808 22772 35860 22778
rect 35808 22714 35860 22720
rect 35256 22704 35308 22710
rect 35256 22646 35308 22652
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 35532 22636 35584 22642
rect 35532 22578 35584 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34808 21486 34836 22170
rect 34980 22092 35032 22098
rect 34980 22034 35032 22040
rect 34992 22001 35020 22034
rect 34978 21992 35034 22001
rect 34978 21927 35034 21936
rect 35360 21894 35388 22578
rect 35072 21888 35124 21894
rect 35072 21830 35124 21836
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 35084 21622 35112 21830
rect 35072 21616 35124 21622
rect 35072 21558 35124 21564
rect 35544 21486 35572 22578
rect 36004 22574 36032 23174
rect 36084 23180 36136 23186
rect 36084 23122 36136 23128
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 36188 22778 36216 23054
rect 36176 22772 36228 22778
rect 36176 22714 36228 22720
rect 35992 22568 36044 22574
rect 35992 22510 36044 22516
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 35624 21684 35676 21690
rect 35624 21626 35676 21632
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 35532 21480 35584 21486
rect 35532 21422 35584 21428
rect 34716 20874 34744 21422
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35440 20936 35492 20942
rect 35438 20904 35440 20913
rect 35492 20904 35494 20913
rect 34704 20868 34756 20874
rect 35438 20839 35494 20848
rect 34704 20810 34756 20816
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 34888 20800 34940 20806
rect 34888 20742 34940 20748
rect 34808 20466 34836 20742
rect 34900 20534 34928 20742
rect 34888 20528 34940 20534
rect 35348 20528 35400 20534
rect 34888 20470 34940 20476
rect 35254 20496 35310 20505
rect 34796 20460 34848 20466
rect 35348 20470 35400 20476
rect 35254 20431 35256 20440
rect 34796 20402 34848 20408
rect 35308 20431 35310 20440
rect 35256 20402 35308 20408
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 19310 34744 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34716 18902 34744 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34704 18896 34756 18902
rect 34704 18838 34756 18844
rect 35360 18834 35388 20470
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34808 17270 34836 18702
rect 35360 18222 35388 18770
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 35452 17066 35480 18906
rect 35532 17604 35584 17610
rect 35532 17546 35584 17552
rect 35440 17060 35492 17066
rect 35440 17002 35492 17008
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35256 16108 35308 16114
rect 35256 16050 35308 16056
rect 35268 15858 35296 16050
rect 35268 15830 35388 15858
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15706 35388 15830
rect 35348 15700 35400 15706
rect 35348 15642 35400 15648
rect 35348 15564 35400 15570
rect 35348 15506 35400 15512
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34704 13320 34756 13326
rect 34704 13262 34756 13268
rect 34716 12986 34744 13262
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34704 12844 34756 12850
rect 34704 12786 34756 12792
rect 34716 11898 34744 12786
rect 34704 11892 34756 11898
rect 34704 11834 34756 11840
rect 34808 11762 34836 13874
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 12918 35388 15506
rect 35544 15502 35572 17546
rect 35532 15496 35584 15502
rect 35532 15438 35584 15444
rect 35544 15162 35572 15438
rect 35532 15156 35584 15162
rect 35532 15098 35584 15104
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35452 13938 35480 14214
rect 35544 14006 35572 15098
rect 35532 14000 35584 14006
rect 35532 13942 35584 13948
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35636 12986 35664 21626
rect 35716 19440 35768 19446
rect 35716 19382 35768 19388
rect 35728 18290 35756 19382
rect 35808 18352 35860 18358
rect 35808 18294 35860 18300
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 35728 17746 35756 18226
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35728 16182 35756 17682
rect 35820 17678 35848 18294
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 36004 17610 36032 22170
rect 36280 21554 36308 24618
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 36096 19854 36124 21422
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 36004 17134 36032 17546
rect 36280 17338 36308 18702
rect 36372 17354 36400 25350
rect 36728 25288 36780 25294
rect 36648 25248 36728 25276
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36464 22094 36492 23666
rect 36544 23180 36596 23186
rect 36544 23122 36596 23128
rect 36556 22574 36584 23122
rect 36648 23118 36676 25248
rect 36728 25230 36780 25236
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36740 23118 36768 24550
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36544 22568 36596 22574
rect 36544 22510 36596 22516
rect 36556 22438 36584 22510
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36648 22234 36676 23054
rect 36636 22228 36688 22234
rect 36636 22170 36688 22176
rect 36464 22066 36584 22094
rect 36556 21010 36584 22066
rect 36728 21344 36780 21350
rect 36728 21286 36780 21292
rect 36740 21078 36768 21286
rect 36728 21072 36780 21078
rect 36728 21014 36780 21020
rect 36544 21004 36596 21010
rect 36544 20946 36596 20952
rect 36740 20874 36768 21014
rect 36728 20868 36780 20874
rect 36728 20810 36780 20816
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36464 18290 36492 18702
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 36544 18080 36596 18086
rect 36544 18022 36596 18028
rect 36556 17678 36584 18022
rect 36544 17672 36596 17678
rect 36544 17614 36596 17620
rect 36268 17332 36320 17338
rect 36372 17326 36492 17354
rect 36268 17274 36320 17280
rect 35992 17128 36044 17134
rect 35992 17070 36044 17076
rect 35808 16584 35860 16590
rect 35808 16526 35860 16532
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 35716 16176 35768 16182
rect 35716 16118 35768 16124
rect 35716 15564 35768 15570
rect 35716 15506 35768 15512
rect 35728 14482 35756 15506
rect 35820 15026 35848 16526
rect 35912 15026 35940 16526
rect 36372 15910 36400 16526
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36372 15434 36400 15846
rect 36360 15428 36412 15434
rect 36360 15370 36412 15376
rect 35808 15020 35860 15026
rect 35808 14962 35860 14968
rect 35900 15020 35952 15026
rect 35952 14980 36032 15008
rect 35900 14962 35952 14968
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35348 12912 35400 12918
rect 35348 12854 35400 12860
rect 35624 12844 35676 12850
rect 35624 12786 35676 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35544 11830 35572 12038
rect 35532 11824 35584 11830
rect 35532 11766 35584 11772
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34808 11218 34836 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35636 11354 35664 12786
rect 35728 12306 35756 14418
rect 35820 13326 35848 14962
rect 35900 14884 35952 14890
rect 35900 14826 35952 14832
rect 35912 14278 35940 14826
rect 36004 14414 36032 14980
rect 35992 14408 36044 14414
rect 35992 14350 36044 14356
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 35912 14074 35940 14214
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 36004 13954 36032 14350
rect 35912 13926 36032 13954
rect 35912 13326 35940 13926
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35900 13320 35952 13326
rect 35900 13262 35952 13268
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 35820 12782 35848 13262
rect 35808 12776 35860 12782
rect 35808 12718 35860 12724
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 35164 11076 35216 11082
rect 35164 11018 35216 11024
rect 35176 10810 35204 11018
rect 35636 10810 35664 11290
rect 35164 10804 35216 10810
rect 35164 10746 35216 10752
rect 35624 10804 35676 10810
rect 35624 10746 35676 10752
rect 35728 10690 35756 12242
rect 36096 12102 36124 13262
rect 36464 12986 36492 17326
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 36556 11898 36584 12038
rect 36832 11898 36860 25638
rect 36924 25294 36952 25758
rect 37384 25684 37412 28358
rect 37476 25838 37504 29260
rect 37556 29164 37608 29170
rect 37556 29106 37608 29112
rect 37648 29164 37700 29170
rect 37648 29106 37700 29112
rect 37568 28558 37596 29106
rect 37660 28626 37688 29106
rect 37648 28620 37700 28626
rect 37648 28562 37700 28568
rect 37556 28552 37608 28558
rect 37556 28494 37608 28500
rect 37660 28150 37688 28562
rect 37648 28144 37700 28150
rect 37648 28086 37700 28092
rect 37556 26376 37608 26382
rect 37660 26364 37688 28086
rect 37752 27062 37780 32166
rect 37936 31385 37964 32438
rect 38028 31754 38056 32778
rect 38120 31890 38148 32966
rect 38108 31884 38160 31890
rect 38108 31826 38160 31832
rect 38016 31748 38068 31754
rect 38016 31690 38068 31696
rect 38016 31476 38068 31482
rect 38016 31418 38068 31424
rect 37922 31376 37978 31385
rect 38028 31346 38056 31418
rect 37922 31311 37924 31320
rect 37976 31311 37978 31320
rect 38016 31340 38068 31346
rect 37924 31282 37976 31288
rect 38016 31282 38068 31288
rect 38028 31226 38056 31282
rect 37844 31198 38056 31226
rect 37844 30394 37872 31198
rect 38120 30784 38148 31826
rect 38028 30756 38148 30784
rect 37924 30592 37976 30598
rect 37924 30534 37976 30540
rect 37832 30388 37884 30394
rect 37832 30330 37884 30336
rect 37936 30190 37964 30534
rect 37924 30184 37976 30190
rect 37924 30126 37976 30132
rect 37936 29578 37964 30126
rect 37924 29572 37976 29578
rect 37924 29514 37976 29520
rect 37832 28076 37884 28082
rect 37832 28018 37884 28024
rect 37740 27056 37792 27062
rect 37740 26998 37792 27004
rect 37740 26852 37792 26858
rect 37740 26794 37792 26800
rect 37752 26382 37780 26794
rect 37844 26382 37872 28018
rect 37924 28008 37976 28014
rect 37924 27950 37976 27956
rect 37936 26994 37964 27950
rect 37924 26988 37976 26994
rect 37924 26930 37976 26936
rect 37608 26336 37688 26364
rect 37740 26376 37792 26382
rect 37556 26318 37608 26324
rect 37740 26318 37792 26324
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 37464 25832 37516 25838
rect 37464 25774 37516 25780
rect 37384 25656 37504 25684
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 36912 25152 36964 25158
rect 36912 25094 36964 25100
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36820 11892 36872 11898
rect 36820 11834 36872 11840
rect 35636 10662 35756 10690
rect 35636 10606 35664 10662
rect 35624 10600 35676 10606
rect 35624 10542 35676 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35636 10198 35664 10542
rect 36924 10198 36952 25094
rect 37188 23724 37240 23730
rect 37188 23666 37240 23672
rect 37200 23186 37228 23666
rect 37188 23180 37240 23186
rect 37188 23122 37240 23128
rect 37004 22976 37056 22982
rect 37004 22918 37056 22924
rect 35624 10192 35676 10198
rect 35624 10134 35676 10140
rect 36912 10192 36964 10198
rect 36912 10134 36964 10140
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34624 6886 34744 6914
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34716 2446 34744 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 37016 4146 37044 22918
rect 37280 22568 37332 22574
rect 37280 22510 37332 22516
rect 37292 21622 37320 22510
rect 37372 22500 37424 22506
rect 37372 22442 37424 22448
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37188 21480 37240 21486
rect 37188 21422 37240 21428
rect 37200 20942 37228 21422
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37188 20800 37240 20806
rect 37240 20748 37320 20754
rect 37188 20742 37320 20748
rect 37200 20726 37320 20742
rect 37292 19990 37320 20726
rect 37384 20398 37412 22442
rect 37476 21690 37504 25656
rect 37568 24274 37596 26318
rect 37648 25288 37700 25294
rect 37648 25230 37700 25236
rect 37660 24274 37688 25230
rect 37556 24268 37608 24274
rect 37556 24210 37608 24216
rect 37648 24268 37700 24274
rect 37648 24210 37700 24216
rect 37568 22574 37596 24210
rect 37844 24206 37872 26318
rect 38028 24750 38056 30756
rect 38108 30660 38160 30666
rect 38108 30602 38160 30608
rect 38120 30190 38148 30602
rect 38108 30184 38160 30190
rect 38108 30126 38160 30132
rect 38212 29102 38240 34478
rect 38304 31657 38332 37266
rect 38752 36168 38804 36174
rect 38856 36156 38884 39306
rect 38948 39098 38976 39374
rect 38936 39092 38988 39098
rect 38936 39034 38988 39040
rect 38804 36128 38884 36156
rect 38752 36110 38804 36116
rect 38764 35834 38792 36110
rect 38752 35828 38804 35834
rect 38752 35770 38804 35776
rect 38384 35692 38436 35698
rect 38384 35634 38436 35640
rect 38396 35086 38424 35634
rect 38384 35080 38436 35086
rect 38384 35022 38436 35028
rect 38396 32910 38424 35022
rect 38476 34740 38528 34746
rect 38476 34682 38528 34688
rect 38384 32904 38436 32910
rect 38384 32846 38436 32852
rect 38488 32722 38516 34682
rect 38660 33448 38712 33454
rect 38660 33390 38712 33396
rect 38396 32694 38516 32722
rect 38290 31648 38346 31657
rect 38290 31583 38346 31592
rect 38290 31240 38346 31249
rect 38290 31175 38346 31184
rect 38304 30580 38332 31175
rect 38396 30734 38424 32694
rect 38672 31906 38700 33390
rect 38844 32836 38896 32842
rect 38844 32778 38896 32784
rect 38856 32434 38884 32778
rect 38936 32768 38988 32774
rect 38936 32710 38988 32716
rect 38948 32502 38976 32710
rect 38936 32496 38988 32502
rect 38936 32438 38988 32444
rect 38844 32428 38896 32434
rect 38844 32370 38896 32376
rect 38580 31878 38700 31906
rect 38476 31816 38528 31822
rect 38476 31758 38528 31764
rect 38488 31521 38516 31758
rect 38580 31754 38608 31878
rect 38660 31816 38712 31822
rect 38660 31758 38712 31764
rect 38568 31748 38620 31754
rect 38568 31690 38620 31696
rect 38566 31648 38622 31657
rect 38566 31583 38622 31592
rect 38474 31512 38530 31521
rect 38474 31447 38530 31456
rect 38384 30728 38436 30734
rect 38384 30670 38436 30676
rect 38304 30552 38424 30580
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38108 29096 38160 29102
rect 38108 29038 38160 29044
rect 38200 29096 38252 29102
rect 38304 29073 38332 29106
rect 38200 29038 38252 29044
rect 38290 29064 38346 29073
rect 38120 28762 38148 29038
rect 38290 28999 38346 29008
rect 38108 28756 38160 28762
rect 38108 28698 38160 28704
rect 38396 27606 38424 30552
rect 38488 29306 38516 31447
rect 38476 29300 38528 29306
rect 38476 29242 38528 29248
rect 38580 29152 38608 31583
rect 38672 31482 38700 31758
rect 38752 31748 38804 31754
rect 38752 31690 38804 31696
rect 38660 31476 38712 31482
rect 38660 31418 38712 31424
rect 38764 31414 38792 31690
rect 38752 31408 38804 31414
rect 38752 31350 38804 31356
rect 38844 31272 38896 31278
rect 38844 31214 38896 31220
rect 38752 31136 38804 31142
rect 38752 31078 38804 31084
rect 38764 30734 38792 31078
rect 38752 30728 38804 30734
rect 38752 30670 38804 30676
rect 38856 30546 38884 31214
rect 38936 30932 38988 30938
rect 38936 30874 38988 30880
rect 38764 30518 38884 30546
rect 38660 29164 38712 29170
rect 38580 29124 38660 29152
rect 38660 29106 38712 29112
rect 38384 27600 38436 27606
rect 38384 27542 38436 27548
rect 38200 26920 38252 26926
rect 38200 26862 38252 26868
rect 38212 26518 38240 26862
rect 38200 26512 38252 26518
rect 38200 26454 38252 26460
rect 38016 24744 38068 24750
rect 38016 24686 38068 24692
rect 38016 24268 38068 24274
rect 38016 24210 38068 24216
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37648 23520 37700 23526
rect 37648 23462 37700 23468
rect 37660 23118 37688 23462
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37844 22642 37872 24142
rect 37832 22636 37884 22642
rect 37752 22596 37832 22624
rect 37556 22568 37608 22574
rect 37556 22510 37608 22516
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37568 21554 37596 22510
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37568 20874 37596 21490
rect 37752 21486 37780 22596
rect 37832 22578 37884 22584
rect 37924 22160 37976 22166
rect 37924 22102 37976 22108
rect 37740 21480 37792 21486
rect 37740 21422 37792 21428
rect 37832 21412 37884 21418
rect 37832 21354 37884 21360
rect 37844 21049 37872 21354
rect 37830 21040 37886 21049
rect 37830 20975 37832 20984
rect 37884 20975 37886 20984
rect 37832 20946 37884 20952
rect 37556 20868 37608 20874
rect 37556 20810 37608 20816
rect 37648 20800 37700 20806
rect 37648 20742 37700 20748
rect 37372 20392 37424 20398
rect 37372 20334 37424 20340
rect 37464 20324 37516 20330
rect 37464 20266 37516 20272
rect 37372 20052 37424 20058
rect 37372 19994 37424 20000
rect 37280 19984 37332 19990
rect 37186 19952 37242 19961
rect 37280 19926 37332 19932
rect 37186 19887 37242 19896
rect 37200 19854 37228 19887
rect 37292 19854 37320 19926
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37384 19378 37412 19994
rect 37476 19854 37504 20266
rect 37556 20256 37608 20262
rect 37556 20198 37608 20204
rect 37568 19854 37596 20198
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37556 19848 37608 19854
rect 37556 19790 37608 19796
rect 37660 19378 37688 20742
rect 37740 20392 37792 20398
rect 37740 20334 37792 20340
rect 37372 19372 37424 19378
rect 37648 19372 37700 19378
rect 37424 19320 37504 19334
rect 37372 19314 37504 19320
rect 37648 19314 37700 19320
rect 37384 19306 37504 19314
rect 37476 17882 37504 19306
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37568 18290 37596 18566
rect 37556 18284 37608 18290
rect 37556 18226 37608 18232
rect 37752 18170 37780 20334
rect 37936 19990 37964 22102
rect 37924 19984 37976 19990
rect 37924 19926 37976 19932
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 37844 19378 37872 19654
rect 37832 19372 37884 19378
rect 37832 19314 37884 19320
rect 37568 18142 37780 18170
rect 37464 17876 37516 17882
rect 37464 17818 37516 17824
rect 37568 17542 37596 18142
rect 37556 17536 37608 17542
rect 37556 17478 37608 17484
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37292 13394 37320 17138
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37476 16114 37504 16390
rect 37568 16250 37596 17478
rect 37740 16448 37792 16454
rect 37740 16390 37792 16396
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37752 15502 37780 16390
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 38028 15026 38056 24210
rect 38212 23322 38240 26454
rect 38200 23316 38252 23322
rect 38200 23258 38252 23264
rect 38396 21350 38424 27542
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38488 23254 38516 27270
rect 38672 26994 38700 29106
rect 38764 29102 38792 30518
rect 38948 30190 38976 30874
rect 38936 30184 38988 30190
rect 38936 30126 38988 30132
rect 38752 29096 38804 29102
rect 38752 29038 38804 29044
rect 38764 27946 38792 29038
rect 38844 28552 38896 28558
rect 38948 28540 38976 30126
rect 39040 28694 39068 44200
rect 42720 42226 42748 44200
rect 43994 42664 44050 42673
rect 43994 42599 44050 42608
rect 44008 42294 44036 42599
rect 43996 42288 44048 42294
rect 43996 42230 44048 42236
rect 41604 42220 41656 42226
rect 41604 42162 41656 42168
rect 42708 42220 42760 42226
rect 42708 42162 42760 42168
rect 41616 41682 41644 42162
rect 41604 41676 41656 41682
rect 41604 41618 41656 41624
rect 40132 41540 40184 41546
rect 40132 41482 40184 41488
rect 39304 41472 39356 41478
rect 39304 41414 39356 41420
rect 39316 39914 39344 41414
rect 40144 41274 40172 41482
rect 41420 41472 41472 41478
rect 41420 41414 41472 41420
rect 40132 41268 40184 41274
rect 40132 41210 40184 41216
rect 40684 41132 40736 41138
rect 40684 41074 40736 41080
rect 40040 41064 40092 41070
rect 40040 41006 40092 41012
rect 39304 39908 39356 39914
rect 39304 39850 39356 39856
rect 39212 39636 39264 39642
rect 39212 39578 39264 39584
rect 39120 39364 39172 39370
rect 39120 39306 39172 39312
rect 39132 39098 39160 39306
rect 39120 39092 39172 39098
rect 39120 39034 39172 39040
rect 39224 38962 39252 39578
rect 39672 39568 39724 39574
rect 39672 39510 39724 39516
rect 39212 38956 39264 38962
rect 39212 38898 39264 38904
rect 39212 38820 39264 38826
rect 39212 38762 39264 38768
rect 39224 38350 39252 38762
rect 39212 38344 39264 38350
rect 39212 38286 39264 38292
rect 39304 38344 39356 38350
rect 39304 38286 39356 38292
rect 39120 38276 39172 38282
rect 39120 38218 39172 38224
rect 39132 37738 39160 38218
rect 39212 38208 39264 38214
rect 39212 38150 39264 38156
rect 39120 37732 39172 37738
rect 39120 37674 39172 37680
rect 39132 37194 39160 37674
rect 39224 37670 39252 38150
rect 39316 37874 39344 38286
rect 39304 37868 39356 37874
rect 39304 37810 39356 37816
rect 39212 37664 39264 37670
rect 39212 37606 39264 37612
rect 39120 37188 39172 37194
rect 39120 37130 39172 37136
rect 39132 36922 39160 37130
rect 39120 36916 39172 36922
rect 39120 36858 39172 36864
rect 39120 36032 39172 36038
rect 39120 35974 39172 35980
rect 39132 35698 39160 35974
rect 39120 35692 39172 35698
rect 39120 35634 39172 35640
rect 39120 31340 39172 31346
rect 39120 31282 39172 31288
rect 39132 30734 39160 31282
rect 39224 31278 39252 37606
rect 39316 37466 39344 37810
rect 39684 37670 39712 39510
rect 39764 38888 39816 38894
rect 39764 38830 39816 38836
rect 39672 37664 39724 37670
rect 39672 37606 39724 37612
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 39488 37460 39540 37466
rect 39488 37402 39540 37408
rect 39316 37244 39344 37402
rect 39500 37262 39528 37402
rect 39396 37256 39448 37262
rect 39316 37216 39396 37244
rect 39396 37198 39448 37204
rect 39488 37256 39540 37262
rect 39488 37198 39540 37204
rect 39408 36106 39436 37198
rect 39396 36100 39448 36106
rect 39396 36042 39448 36048
rect 39304 36032 39356 36038
rect 39304 35974 39356 35980
rect 39316 33590 39344 35974
rect 39304 33584 39356 33590
rect 39304 33526 39356 33532
rect 39408 33454 39436 36042
rect 39396 33448 39448 33454
rect 39396 33390 39448 33396
rect 39304 31680 39356 31686
rect 39304 31622 39356 31628
rect 39212 31272 39264 31278
rect 39212 31214 39264 31220
rect 39212 31136 39264 31142
rect 39212 31078 39264 31084
rect 39224 30938 39252 31078
rect 39212 30932 39264 30938
rect 39212 30874 39264 30880
rect 39120 30728 39172 30734
rect 39120 30670 39172 30676
rect 39212 30592 39264 30598
rect 39212 30534 39264 30540
rect 39224 30326 39252 30534
rect 39212 30320 39264 30326
rect 39212 30262 39264 30268
rect 39316 30258 39344 31622
rect 39408 31346 39436 33390
rect 39580 32836 39632 32842
rect 39580 32778 39632 32784
rect 39488 32768 39540 32774
rect 39488 32710 39540 32716
rect 39500 32434 39528 32710
rect 39592 32570 39620 32778
rect 39580 32564 39632 32570
rect 39580 32506 39632 32512
rect 39488 32428 39540 32434
rect 39488 32370 39540 32376
rect 39580 31748 39632 31754
rect 39580 31690 39632 31696
rect 39396 31340 39448 31346
rect 39396 31282 39448 31288
rect 39488 31340 39540 31346
rect 39488 31282 39540 31288
rect 39304 30252 39356 30258
rect 39304 30194 39356 30200
rect 39396 29504 39448 29510
rect 39396 29446 39448 29452
rect 39212 29300 39264 29306
rect 39212 29242 39264 29248
rect 39224 29170 39252 29242
rect 39408 29170 39436 29446
rect 39120 29164 39172 29170
rect 39120 29106 39172 29112
rect 39212 29164 39264 29170
rect 39212 29106 39264 29112
rect 39396 29164 39448 29170
rect 39396 29106 39448 29112
rect 39132 28762 39160 29106
rect 39120 28756 39172 28762
rect 39120 28698 39172 28704
rect 39028 28688 39080 28694
rect 39028 28630 39080 28636
rect 38896 28512 38976 28540
rect 38844 28494 38896 28500
rect 38856 28150 38884 28494
rect 39028 28484 39080 28490
rect 38948 28444 39028 28472
rect 38844 28144 38896 28150
rect 38844 28086 38896 28092
rect 38752 27940 38804 27946
rect 38752 27882 38804 27888
rect 38660 26988 38712 26994
rect 38660 26930 38712 26936
rect 38672 26897 38700 26930
rect 38658 26888 38714 26897
rect 38658 26823 38714 26832
rect 38856 26738 38884 28086
rect 38672 26710 38884 26738
rect 38672 26382 38700 26710
rect 38660 26376 38712 26382
rect 38712 26336 38792 26364
rect 38660 26318 38712 26324
rect 38660 25900 38712 25906
rect 38580 25860 38660 25888
rect 38580 25770 38608 25860
rect 38660 25842 38712 25848
rect 38568 25764 38620 25770
rect 38568 25706 38620 25712
rect 38764 24834 38792 26336
rect 38948 26314 38976 28444
rect 39028 28426 39080 28432
rect 39028 27600 39080 27606
rect 39028 27542 39080 27548
rect 39040 27470 39068 27542
rect 39028 27464 39080 27470
rect 39028 27406 39080 27412
rect 39028 26988 39080 26994
rect 39028 26930 39080 26936
rect 39120 26988 39172 26994
rect 39224 26976 39252 29106
rect 39304 28960 39356 28966
rect 39304 28902 39356 28908
rect 39316 28558 39344 28902
rect 39304 28552 39356 28558
rect 39304 28494 39356 28500
rect 39172 26948 39252 26976
rect 39120 26930 39172 26936
rect 39040 26314 39068 26930
rect 38936 26308 38988 26314
rect 38936 26250 38988 26256
rect 39028 26308 39080 26314
rect 39028 26250 39080 26256
rect 38844 26240 38896 26246
rect 38844 26182 38896 26188
rect 38856 25906 38884 26182
rect 38844 25900 38896 25906
rect 38844 25842 38896 25848
rect 38948 25786 38976 26250
rect 39120 26240 39172 26246
rect 39120 26182 39172 26188
rect 39132 25906 39160 26182
rect 39120 25900 39172 25906
rect 39120 25842 39172 25848
rect 38580 24818 38792 24834
rect 38856 25758 38976 25786
rect 38856 24818 38884 25758
rect 39028 25696 39080 25702
rect 39028 25638 39080 25644
rect 39040 25362 39068 25638
rect 39224 25378 39252 26948
rect 39316 26382 39344 28494
rect 39408 26908 39436 29106
rect 39500 28422 39528 31282
rect 39592 30802 39620 31690
rect 39580 30796 39632 30802
rect 39580 30738 39632 30744
rect 39488 28416 39540 28422
rect 39488 28358 39540 28364
rect 39500 28082 39528 28358
rect 39488 28076 39540 28082
rect 39488 28018 39540 28024
rect 39408 26880 39620 26908
rect 39488 26784 39540 26790
rect 39488 26726 39540 26732
rect 39304 26376 39356 26382
rect 39356 26336 39436 26364
rect 39304 26318 39356 26324
rect 39028 25356 39080 25362
rect 39028 25298 39080 25304
rect 39132 25350 39252 25378
rect 38936 25288 38988 25294
rect 38936 25230 38988 25236
rect 38948 24954 38976 25230
rect 38936 24948 38988 24954
rect 38936 24890 38988 24896
rect 38568 24812 38792 24818
rect 38620 24806 38792 24812
rect 38568 24754 38620 24760
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38672 24070 38700 24550
rect 38660 24064 38712 24070
rect 38660 24006 38712 24012
rect 38476 23248 38528 23254
rect 38476 23190 38528 23196
rect 38764 23118 38792 24806
rect 38844 24812 38896 24818
rect 38844 24754 38896 24760
rect 38936 24812 38988 24818
rect 39132 24800 39160 25350
rect 39212 25288 39264 25294
rect 39212 25230 39264 25236
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 38936 24754 38988 24760
rect 39040 24772 39160 24800
rect 38948 24342 38976 24754
rect 38936 24336 38988 24342
rect 38842 24304 38898 24313
rect 38936 24278 38988 24284
rect 38842 24239 38898 24248
rect 38856 24206 38884 24239
rect 39040 24206 39068 24772
rect 39120 24676 39172 24682
rect 39120 24618 39172 24624
rect 38844 24200 38896 24206
rect 38844 24142 38896 24148
rect 39028 24200 39080 24206
rect 39028 24142 39080 24148
rect 38752 23112 38804 23118
rect 38752 23054 38804 23060
rect 38660 22636 38712 22642
rect 38660 22578 38712 22584
rect 38672 21554 38700 22578
rect 38764 22094 38792 23054
rect 38856 22642 38884 24142
rect 38936 24064 38988 24070
rect 38934 24032 38936 24041
rect 38988 24032 38990 24041
rect 38934 23967 38990 23976
rect 39040 23662 39068 24142
rect 39028 23656 39080 23662
rect 39028 23598 39080 23604
rect 39026 23488 39082 23497
rect 39026 23423 39082 23432
rect 39040 23118 39068 23423
rect 39028 23112 39080 23118
rect 39028 23054 39080 23060
rect 39132 23050 39160 24618
rect 39224 24410 39252 25230
rect 39316 24954 39344 25230
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 39408 24818 39436 26336
rect 39500 25974 39528 26726
rect 39488 25968 39540 25974
rect 39488 25910 39540 25916
rect 39396 24812 39448 24818
rect 39396 24754 39448 24760
rect 39488 24812 39540 24818
rect 39488 24754 39540 24760
rect 39212 24404 39264 24410
rect 39212 24346 39264 24352
rect 39212 24132 39264 24138
rect 39212 24074 39264 24080
rect 39224 24041 39252 24074
rect 39210 24032 39266 24041
rect 39210 23967 39266 23976
rect 39212 23656 39264 23662
rect 39212 23598 39264 23604
rect 39120 23044 39172 23050
rect 39120 22986 39172 22992
rect 39028 22976 39080 22982
rect 39028 22918 39080 22924
rect 39040 22642 39068 22918
rect 38844 22636 38896 22642
rect 38844 22578 38896 22584
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 39132 22166 39160 22986
rect 39224 22642 39252 23598
rect 39408 23118 39436 24754
rect 39500 24410 39528 24754
rect 39488 24404 39540 24410
rect 39488 24346 39540 24352
rect 39592 24206 39620 26880
rect 39684 26450 39712 37606
rect 39776 36242 39804 38830
rect 39856 37188 39908 37194
rect 39856 37130 39908 37136
rect 39764 36236 39816 36242
rect 39764 36178 39816 36184
rect 39776 36009 39804 36178
rect 39762 36000 39818 36009
rect 39762 35935 39818 35944
rect 39868 31754 39896 37130
rect 39948 36916 40000 36922
rect 39948 36858 40000 36864
rect 39960 36038 39988 36858
rect 39948 36032 40000 36038
rect 39948 35974 40000 35980
rect 40052 35154 40080 41006
rect 40696 40730 40724 41074
rect 40684 40724 40736 40730
rect 40684 40666 40736 40672
rect 40132 40588 40184 40594
rect 40132 40530 40184 40536
rect 40144 39846 40172 40530
rect 40408 39908 40460 39914
rect 40408 39850 40460 39856
rect 40132 39840 40184 39846
rect 40132 39782 40184 39788
rect 40420 38350 40448 39850
rect 41432 39642 41460 41414
rect 41512 40928 41564 40934
rect 41512 40870 41564 40876
rect 40960 39636 41012 39642
rect 40960 39578 41012 39584
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 40972 38758 41000 39578
rect 41524 39386 41552 40870
rect 41340 39358 41552 39386
rect 41340 39302 41368 39358
rect 41328 39296 41380 39302
rect 41328 39238 41380 39244
rect 41420 39296 41472 39302
rect 41420 39238 41472 39244
rect 40960 38752 41012 38758
rect 40960 38694 41012 38700
rect 40408 38344 40460 38350
rect 40408 38286 40460 38292
rect 40408 38208 40460 38214
rect 40408 38150 40460 38156
rect 40420 37806 40448 38150
rect 40972 37942 41000 38694
rect 41144 38344 41196 38350
rect 41144 38286 41196 38292
rect 40960 37936 41012 37942
rect 40960 37878 41012 37884
rect 41156 37874 41184 38286
rect 41144 37868 41196 37874
rect 41144 37810 41196 37816
rect 40408 37800 40460 37806
rect 40408 37742 40460 37748
rect 40420 37194 40448 37742
rect 40500 37392 40552 37398
rect 40500 37334 40552 37340
rect 40512 37262 40540 37334
rect 41156 37262 41184 37810
rect 40500 37256 40552 37262
rect 40500 37198 40552 37204
rect 41144 37256 41196 37262
rect 41144 37198 41196 37204
rect 40408 37188 40460 37194
rect 40408 37130 40460 37136
rect 40316 35488 40368 35494
rect 40316 35430 40368 35436
rect 40040 35148 40092 35154
rect 40040 35090 40092 35096
rect 40328 34678 40356 35430
rect 40420 35000 40448 37130
rect 40960 36032 41012 36038
rect 40960 35974 41012 35980
rect 40972 35698 41000 35974
rect 40960 35692 41012 35698
rect 40960 35634 41012 35640
rect 41156 35562 41184 37198
rect 41340 35698 41368 39238
rect 41432 37398 41460 39238
rect 41420 37392 41472 37398
rect 41420 37334 41472 37340
rect 41616 36786 41644 41618
rect 41880 41608 41932 41614
rect 41880 41550 41932 41556
rect 41892 40526 41920 41550
rect 43996 41540 44048 41546
rect 43996 41482 44048 41488
rect 44008 41177 44036 41482
rect 43994 41168 44050 41177
rect 43076 41132 43128 41138
rect 43994 41103 44050 41112
rect 43076 41074 43128 41080
rect 41880 40520 41932 40526
rect 41880 40462 41932 40468
rect 41788 39432 41840 39438
rect 41788 39374 41840 39380
rect 41800 38418 41828 39374
rect 41788 38412 41840 38418
rect 41788 38354 41840 38360
rect 41800 37262 41828 38354
rect 41788 37256 41840 37262
rect 41708 37216 41788 37244
rect 41604 36780 41656 36786
rect 41604 36722 41656 36728
rect 41236 35692 41288 35698
rect 41236 35634 41288 35640
rect 41328 35692 41380 35698
rect 41328 35634 41380 35640
rect 41144 35556 41196 35562
rect 41144 35498 41196 35504
rect 40592 35012 40644 35018
rect 40420 34972 40592 35000
rect 40592 34954 40644 34960
rect 40316 34672 40368 34678
rect 40316 34614 40368 34620
rect 40328 33590 40356 34614
rect 40316 33584 40368 33590
rect 40316 33526 40368 33532
rect 40604 33522 40632 34954
rect 40776 34944 40828 34950
rect 40776 34886 40828 34892
rect 40592 33516 40644 33522
rect 40592 33458 40644 33464
rect 40040 32768 40092 32774
rect 40040 32710 40092 32716
rect 39948 32496 40000 32502
rect 39948 32438 40000 32444
rect 39776 31726 39896 31754
rect 39672 26444 39724 26450
rect 39672 26386 39724 26392
rect 39776 24614 39804 31726
rect 39960 30258 39988 32438
rect 40052 31890 40080 32710
rect 40408 32224 40460 32230
rect 40408 32166 40460 32172
rect 40040 31884 40092 31890
rect 40040 31826 40092 31832
rect 40052 30802 40080 31826
rect 40420 31822 40448 32166
rect 40408 31816 40460 31822
rect 40408 31758 40460 31764
rect 40604 31754 40632 33458
rect 40592 31748 40644 31754
rect 40592 31690 40644 31696
rect 40788 31686 40816 34886
rect 41156 33522 41184 35498
rect 41248 35018 41276 35634
rect 41236 35012 41288 35018
rect 41236 34954 41288 34960
rect 41144 33516 41196 33522
rect 41144 33458 41196 33464
rect 40960 32360 41012 32366
rect 40960 32302 41012 32308
rect 40972 32026 41000 32302
rect 40960 32020 41012 32026
rect 40960 31962 41012 31968
rect 41156 31754 41184 33458
rect 41052 31748 41184 31754
rect 41104 31726 41184 31748
rect 41052 31690 41104 31696
rect 40776 31680 40828 31686
rect 40776 31622 40828 31628
rect 40040 30796 40092 30802
rect 40040 30738 40092 30744
rect 40408 30796 40460 30802
rect 40408 30738 40460 30744
rect 40224 30728 40276 30734
rect 40224 30670 40276 30676
rect 40236 30326 40264 30670
rect 40224 30320 40276 30326
rect 40224 30262 40276 30268
rect 39948 30252 40000 30258
rect 39948 30194 40000 30200
rect 40316 30252 40368 30258
rect 40316 30194 40368 30200
rect 39960 29238 39988 30194
rect 40132 30184 40184 30190
rect 40132 30126 40184 30132
rect 40040 29504 40092 29510
rect 40040 29446 40092 29452
rect 39948 29232 40000 29238
rect 39948 29174 40000 29180
rect 40052 29034 40080 29446
rect 40144 29170 40172 30126
rect 40328 29170 40356 30194
rect 40132 29164 40184 29170
rect 40132 29106 40184 29112
rect 40316 29164 40368 29170
rect 40316 29106 40368 29112
rect 40040 29028 40092 29034
rect 40040 28970 40092 28976
rect 40052 28558 40080 28970
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 40144 27606 40172 29106
rect 40224 29096 40276 29102
rect 40420 29050 40448 30738
rect 40276 29044 40448 29050
rect 40224 29038 40448 29044
rect 40236 29022 40448 29038
rect 40236 28626 40264 29022
rect 40224 28620 40276 28626
rect 40224 28562 40276 28568
rect 40132 27600 40184 27606
rect 40132 27542 40184 27548
rect 40040 26784 40092 26790
rect 40040 26726 40092 26732
rect 40052 26042 40080 26726
rect 40040 26036 40092 26042
rect 40040 25978 40092 25984
rect 40132 25900 40184 25906
rect 40132 25842 40184 25848
rect 40144 24818 40172 25842
rect 40236 25362 40264 28562
rect 40316 28552 40368 28558
rect 40316 28494 40368 28500
rect 40328 28218 40356 28494
rect 40316 28212 40368 28218
rect 40316 28154 40368 28160
rect 40684 27464 40736 27470
rect 40684 27406 40736 27412
rect 40316 27396 40368 27402
rect 40316 27338 40368 27344
rect 40328 26450 40356 27338
rect 40316 26444 40368 26450
rect 40316 26386 40368 26392
rect 40328 25770 40356 26386
rect 40696 26382 40724 27406
rect 40788 27334 40816 31622
rect 41064 31482 41092 31690
rect 41052 31476 41104 31482
rect 41052 31418 41104 31424
rect 41340 30682 41368 35634
rect 41420 35080 41472 35086
rect 41420 35022 41472 35028
rect 41432 32910 41460 35022
rect 41420 32904 41472 32910
rect 41420 32846 41472 32852
rect 41708 30802 41736 37216
rect 41788 37198 41840 37204
rect 41892 37074 41920 40462
rect 42616 40452 42668 40458
rect 42616 40394 42668 40400
rect 42628 40186 42656 40394
rect 42892 40384 42944 40390
rect 42892 40326 42944 40332
rect 42616 40180 42668 40186
rect 42616 40122 42668 40128
rect 42904 40118 42932 40326
rect 42892 40112 42944 40118
rect 42892 40054 42944 40060
rect 42708 39432 42760 39438
rect 42708 39374 42760 39380
rect 42720 38894 42748 39374
rect 42708 38888 42760 38894
rect 42708 38830 42760 38836
rect 42616 38752 42668 38758
rect 42616 38694 42668 38700
rect 42628 38350 42656 38694
rect 42616 38344 42668 38350
rect 42616 38286 42668 38292
rect 42720 38010 42748 38830
rect 42904 38282 42932 40054
rect 43088 39982 43116 41074
rect 43996 41064 44048 41070
rect 43996 41006 44048 41012
rect 43076 39976 43128 39982
rect 43076 39918 43128 39924
rect 43168 39976 43220 39982
rect 43168 39918 43220 39924
rect 42984 38956 43036 38962
rect 42984 38898 43036 38904
rect 42996 38332 43024 38898
rect 43088 38554 43116 39918
rect 43180 38894 43208 39918
rect 44008 39681 44036 41006
rect 43994 39672 44050 39681
rect 43994 39607 44050 39616
rect 43996 39364 44048 39370
rect 43996 39306 44048 39312
rect 43168 38888 43220 38894
rect 43168 38830 43220 38836
rect 43076 38548 43128 38554
rect 43076 38490 43128 38496
rect 42996 38304 43116 38332
rect 42892 38276 42944 38282
rect 42892 38218 42944 38224
rect 43088 38214 43116 38304
rect 43076 38208 43128 38214
rect 43076 38150 43128 38156
rect 42708 38004 42760 38010
rect 42708 37946 42760 37952
rect 43088 37942 43116 38150
rect 43076 37936 43128 37942
rect 43076 37878 43128 37884
rect 42984 37868 43036 37874
rect 42984 37810 43036 37816
rect 42616 37188 42668 37194
rect 42616 37130 42668 37136
rect 41800 37046 41920 37074
rect 41800 35766 41828 37046
rect 42628 36922 42656 37130
rect 42996 37126 43024 37810
rect 42984 37120 43036 37126
rect 42984 37062 43036 37068
rect 43076 37120 43128 37126
rect 43076 37062 43128 37068
rect 42996 36922 43024 37062
rect 42616 36916 42668 36922
rect 42616 36858 42668 36864
rect 42984 36916 43036 36922
rect 42984 36858 43036 36864
rect 43088 36786 43116 37062
rect 43076 36780 43128 36786
rect 43076 36722 43128 36728
rect 43180 36718 43208 38830
rect 44008 38185 44036 39306
rect 43994 38176 44050 38185
rect 43994 38111 44050 38120
rect 43996 37800 44048 37806
rect 43996 37742 44048 37748
rect 43168 36712 43220 36718
rect 44008 36689 44036 37742
rect 43168 36654 43220 36660
rect 43994 36680 44050 36689
rect 41880 36168 41932 36174
rect 41880 36110 41932 36116
rect 41788 35760 41840 35766
rect 41788 35702 41840 35708
rect 41800 34066 41828 35702
rect 41892 35086 41920 36110
rect 42616 36100 42668 36106
rect 42616 36042 42668 36048
rect 42628 35834 42656 36042
rect 42616 35828 42668 35834
rect 42616 35770 42668 35776
rect 41972 35624 42024 35630
rect 43180 35612 43208 36654
rect 43994 36615 44050 36624
rect 43260 36032 43312 36038
rect 43260 35974 43312 35980
rect 43272 35766 43300 35974
rect 43260 35760 43312 35766
rect 43260 35702 43312 35708
rect 43260 35624 43312 35630
rect 43180 35584 43260 35612
rect 41972 35566 42024 35572
rect 43260 35566 43312 35572
rect 41984 35086 42012 35566
rect 41880 35080 41932 35086
rect 41880 35022 41932 35028
rect 41972 35080 42024 35086
rect 41972 35022 42024 35028
rect 42892 35080 42944 35086
rect 42892 35022 42944 35028
rect 41788 34060 41840 34066
rect 41788 34002 41840 34008
rect 41800 32026 41828 34002
rect 42616 33924 42668 33930
rect 42616 33866 42668 33872
rect 42628 33658 42656 33866
rect 42616 33652 42668 33658
rect 42616 33594 42668 33600
rect 42904 33386 42932 35022
rect 43272 34406 43300 35566
rect 43994 35184 44050 35193
rect 43994 35119 43996 35128
rect 44048 35119 44050 35128
rect 43996 35090 44048 35096
rect 43996 35012 44048 35018
rect 43996 34954 44048 34960
rect 43260 34400 43312 34406
rect 43260 34342 43312 34348
rect 42984 33856 43036 33862
rect 42984 33798 43036 33804
rect 42996 33590 43024 33798
rect 42984 33584 43036 33590
rect 42984 33526 43036 33532
rect 43272 33454 43300 34342
rect 44008 33697 44036 34954
rect 43994 33688 44050 33697
rect 43994 33623 44050 33632
rect 43260 33448 43312 33454
rect 43260 33390 43312 33396
rect 42892 33380 42944 33386
rect 42892 33322 42944 33328
rect 41880 32904 41932 32910
rect 41880 32846 41932 32852
rect 42892 32904 42944 32910
rect 42892 32846 42944 32852
rect 41788 32020 41840 32026
rect 41788 31962 41840 31968
rect 41696 30796 41748 30802
rect 41696 30738 41748 30744
rect 41064 30654 41368 30682
rect 41064 30054 41092 30654
rect 41052 30048 41104 30054
rect 41052 29990 41104 29996
rect 41144 30048 41196 30054
rect 41144 29990 41196 29996
rect 41156 29646 41184 29990
rect 41708 29850 41736 30738
rect 41696 29844 41748 29850
rect 41696 29786 41748 29792
rect 41144 29640 41196 29646
rect 41144 29582 41196 29588
rect 41052 29504 41104 29510
rect 41052 29446 41104 29452
rect 41064 29306 41092 29446
rect 41052 29300 41104 29306
rect 41052 29242 41104 29248
rect 41144 29164 41196 29170
rect 41144 29106 41196 29112
rect 40776 27328 40828 27334
rect 40776 27270 40828 27276
rect 40776 26988 40828 26994
rect 40776 26930 40828 26936
rect 40788 26586 40816 26930
rect 40776 26580 40828 26586
rect 40776 26522 40828 26528
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 40316 25764 40368 25770
rect 40316 25706 40368 25712
rect 40696 25498 40724 26318
rect 41156 25906 41184 29106
rect 41892 28558 41920 32846
rect 42904 32366 42932 32846
rect 43168 32836 43220 32842
rect 43168 32778 43220 32784
rect 42984 32428 43036 32434
rect 42984 32370 43036 32376
rect 42892 32360 42944 32366
rect 42892 32302 42944 32308
rect 42616 32224 42668 32230
rect 42616 32166 42668 32172
rect 42628 31822 42656 32166
rect 42996 31958 43024 32370
rect 43180 32201 43208 32778
rect 43272 32366 43300 33390
rect 43260 32360 43312 32366
rect 43260 32302 43312 32308
rect 43166 32192 43222 32201
rect 43166 32127 43222 32136
rect 42984 31952 43036 31958
rect 42984 31894 43036 31900
rect 42616 31816 42668 31822
rect 42616 31758 42668 31764
rect 43076 31340 43128 31346
rect 43076 31282 43128 31288
rect 42984 30932 43036 30938
rect 42984 30874 43036 30880
rect 42616 30660 42668 30666
rect 42616 30602 42668 30608
rect 42628 30394 42656 30602
rect 42996 30394 43024 30874
rect 43088 30598 43116 31282
rect 43168 31272 43220 31278
rect 43168 31214 43220 31220
rect 43180 30705 43208 31214
rect 43166 30696 43222 30705
rect 43166 30631 43222 30640
rect 43076 30592 43128 30598
rect 43076 30534 43128 30540
rect 43088 30394 43116 30534
rect 42616 30388 42668 30394
rect 42616 30330 42668 30336
rect 42984 30388 43036 30394
rect 42984 30330 43036 30336
rect 43076 30388 43128 30394
rect 43076 30330 43128 30336
rect 43260 30116 43312 30122
rect 43260 30058 43312 30064
rect 43168 29572 43220 29578
rect 43168 29514 43220 29520
rect 43180 29209 43208 29514
rect 43166 29200 43222 29209
rect 43166 29135 43222 29144
rect 42984 28756 43036 28762
rect 42984 28698 43036 28704
rect 41880 28552 41932 28558
rect 41880 28494 41932 28500
rect 41892 27470 41920 28494
rect 42616 28484 42668 28490
rect 42616 28426 42668 28432
rect 42628 28218 42656 28426
rect 42996 28218 43024 28698
rect 43076 28416 43128 28422
rect 43076 28358 43128 28364
rect 43088 28218 43116 28358
rect 42616 28212 42668 28218
rect 42616 28154 42668 28160
rect 42984 28212 43036 28218
rect 42984 28154 43036 28160
rect 43076 28212 43128 28218
rect 43076 28154 43128 28160
rect 43088 27470 43116 28154
rect 43272 28014 43300 30058
rect 43260 28008 43312 28014
rect 43260 27950 43312 27956
rect 41880 27464 41932 27470
rect 41880 27406 41932 27412
rect 43076 27464 43128 27470
rect 43076 27406 43128 27412
rect 41972 26988 42024 26994
rect 41972 26930 42024 26936
rect 42984 26988 43036 26994
rect 42984 26930 43036 26936
rect 41984 26450 42012 26930
rect 42616 26784 42668 26790
rect 42616 26726 42668 26732
rect 41972 26444 42024 26450
rect 41972 26386 42024 26392
rect 41144 25900 41196 25906
rect 41144 25842 41196 25848
rect 40684 25492 40736 25498
rect 40684 25434 40736 25440
rect 40224 25356 40276 25362
rect 40224 25298 40276 25304
rect 39948 24812 40000 24818
rect 39948 24754 40000 24760
rect 40132 24812 40184 24818
rect 40132 24754 40184 24760
rect 39764 24608 39816 24614
rect 39764 24550 39816 24556
rect 39580 24200 39632 24206
rect 39580 24142 39632 24148
rect 39592 23594 39620 24142
rect 39960 23866 39988 24754
rect 39948 23860 40000 23866
rect 39948 23802 40000 23808
rect 39580 23588 39632 23594
rect 39580 23530 39632 23536
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 39224 22438 39252 22578
rect 39304 22568 39356 22574
rect 39304 22510 39356 22516
rect 39212 22432 39264 22438
rect 39212 22374 39264 22380
rect 39120 22160 39172 22166
rect 39120 22102 39172 22108
rect 38764 22066 38976 22094
rect 38660 21548 38712 21554
rect 38660 21490 38712 21496
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38384 21344 38436 21350
rect 38384 21286 38436 21292
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 38212 17202 38240 20878
rect 38764 20398 38792 21490
rect 38948 20754 38976 22066
rect 39224 21690 39252 22374
rect 39316 22094 39344 22510
rect 39408 22250 39436 23054
rect 39592 22642 39620 23530
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39580 22432 39632 22438
rect 39580 22374 39632 22380
rect 39408 22222 39528 22250
rect 39316 22066 39436 22094
rect 39304 21888 39356 21894
rect 39304 21830 39356 21836
rect 39316 21690 39344 21830
rect 39212 21684 39264 21690
rect 39212 21626 39264 21632
rect 39304 21684 39356 21690
rect 39304 21626 39356 21632
rect 39316 21010 39344 21626
rect 39408 21554 39436 22066
rect 39396 21548 39448 21554
rect 39396 21490 39448 21496
rect 39396 21344 39448 21350
rect 39396 21286 39448 21292
rect 39408 21010 39436 21286
rect 39304 21004 39356 21010
rect 39304 20946 39356 20952
rect 39396 21004 39448 21010
rect 39396 20946 39448 20952
rect 38856 20726 38976 20754
rect 39304 20800 39356 20806
rect 39304 20742 39356 20748
rect 38856 20466 38884 20726
rect 39028 20596 39080 20602
rect 39028 20538 39080 20544
rect 38844 20460 38896 20466
rect 38844 20402 38896 20408
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38856 19854 38884 20402
rect 38934 20360 38990 20369
rect 38934 20295 38990 20304
rect 38948 19854 38976 20295
rect 39040 19990 39068 20538
rect 39120 20460 39172 20466
rect 39120 20402 39172 20408
rect 39028 19984 39080 19990
rect 39028 19926 39080 19932
rect 39040 19854 39068 19926
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 38844 19848 38896 19854
rect 38844 19790 38896 19796
rect 38936 19848 38988 19854
rect 38936 19790 38988 19796
rect 39028 19848 39080 19854
rect 39132 19825 39160 20402
rect 39028 19790 39080 19796
rect 39118 19816 39174 19825
rect 38764 19718 38792 19790
rect 39118 19751 39174 19760
rect 38752 19712 38804 19718
rect 38752 19654 38804 19660
rect 38844 19508 38896 19514
rect 38844 19450 38896 19456
rect 38856 18426 38884 19450
rect 39316 19446 39344 20742
rect 39500 20466 39528 22222
rect 39592 21894 39620 22374
rect 39580 21888 39632 21894
rect 39580 21830 39632 21836
rect 39764 21888 39816 21894
rect 39764 21830 39816 21836
rect 39776 20942 39804 21830
rect 39960 21690 39988 23802
rect 40236 23186 40264 25298
rect 40316 25220 40368 25226
rect 40316 25162 40368 25168
rect 40408 25220 40460 25226
rect 40408 25162 40460 25168
rect 40328 24682 40356 25162
rect 40316 24676 40368 24682
rect 40316 24618 40368 24624
rect 40328 24274 40356 24618
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 40420 24206 40448 25162
rect 41984 24818 42012 26386
rect 42628 26382 42656 26726
rect 42996 26586 43024 26930
rect 43272 26926 43300 27950
rect 43994 27704 44050 27713
rect 43994 27639 44050 27648
rect 44008 27538 44036 27639
rect 43996 27532 44048 27538
rect 43996 27474 44048 27480
rect 43076 26920 43128 26926
rect 43076 26862 43128 26868
rect 43260 26920 43312 26926
rect 43260 26862 43312 26868
rect 42984 26580 43036 26586
rect 42984 26522 43036 26528
rect 42616 26376 42668 26382
rect 42616 26318 42668 26324
rect 43088 25906 43116 26862
rect 43166 26208 43222 26217
rect 43166 26143 43222 26152
rect 43180 25974 43208 26143
rect 43168 25968 43220 25974
rect 43168 25910 43220 25916
rect 43076 25900 43128 25906
rect 43076 25842 43128 25848
rect 43076 25288 43128 25294
rect 43076 25230 43128 25236
rect 43088 24954 43116 25230
rect 43076 24948 43128 24954
rect 43076 24890 43128 24896
rect 40776 24812 40828 24818
rect 40776 24754 40828 24760
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 42984 24812 43036 24818
rect 42984 24754 43036 24760
rect 40788 24410 40816 24754
rect 40776 24404 40828 24410
rect 40776 24346 40828 24352
rect 41984 24274 42012 24754
rect 42616 24608 42668 24614
rect 42616 24550 42668 24556
rect 41972 24268 42024 24274
rect 41972 24210 42024 24216
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 40224 23180 40276 23186
rect 40224 23122 40276 23128
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 40052 22030 40080 23054
rect 40132 22228 40184 22234
rect 40132 22170 40184 22176
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40052 21690 40080 21966
rect 40144 21962 40172 22170
rect 40132 21956 40184 21962
rect 40132 21898 40184 21904
rect 39948 21684 40000 21690
rect 39948 21626 40000 21632
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 40144 21010 40172 21898
rect 40132 21004 40184 21010
rect 40132 20946 40184 20952
rect 39764 20936 39816 20942
rect 39764 20878 39816 20884
rect 39488 20460 39540 20466
rect 39488 20402 39540 20408
rect 39500 19854 39528 20402
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 39672 19848 39724 19854
rect 39672 19790 39724 19796
rect 39684 19514 39712 19790
rect 39776 19514 39804 20878
rect 40132 20868 40184 20874
rect 40132 20810 40184 20816
rect 40144 20482 40172 20810
rect 40052 20466 40172 20482
rect 40052 20460 40184 20466
rect 40052 20454 40132 20460
rect 40052 20058 40080 20454
rect 40132 20402 40184 20408
rect 40236 20346 40264 23122
rect 40316 23112 40368 23118
rect 40316 23054 40368 23060
rect 40328 22778 40356 23054
rect 40316 22772 40368 22778
rect 40316 22714 40368 22720
rect 40420 22098 40448 24142
rect 41984 22114 42012 24210
rect 42628 24206 42656 24550
rect 42996 24410 43024 24754
rect 43272 24750 43300 26862
rect 43996 25220 44048 25226
rect 43996 25162 44048 25168
rect 43260 24744 43312 24750
rect 44008 24721 44036 25162
rect 43260 24686 43312 24692
rect 43994 24712 44050 24721
rect 42984 24404 43036 24410
rect 42984 24346 43036 24352
rect 42616 24200 42668 24206
rect 42616 24142 42668 24148
rect 42708 23724 42760 23730
rect 42708 23666 42760 23672
rect 42720 23186 42748 23666
rect 43076 23316 43128 23322
rect 43076 23258 43128 23264
rect 42708 23180 42760 23186
rect 42708 23122 42760 23128
rect 42064 22976 42116 22982
rect 42064 22918 42116 22924
rect 40408 22092 40460 22098
rect 40408 22034 40460 22040
rect 41892 22086 42012 22114
rect 41892 22030 41920 22086
rect 41880 22024 41932 22030
rect 41880 21966 41932 21972
rect 41984 21554 42012 22086
rect 42076 22030 42104 22918
rect 42064 22024 42116 22030
rect 42064 21966 42116 21972
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 41972 21548 42024 21554
rect 41972 21490 42024 21496
rect 42708 21548 42760 21554
rect 42708 21490 42760 21496
rect 40316 21412 40368 21418
rect 40316 21354 40368 21360
rect 40144 20318 40264 20346
rect 40144 20262 40172 20318
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 40040 20052 40092 20058
rect 40040 19994 40092 20000
rect 40144 19922 40172 20198
rect 40132 19916 40184 19922
rect 40132 19858 40184 19864
rect 39672 19508 39724 19514
rect 39672 19450 39724 19456
rect 39764 19508 39816 19514
rect 39764 19450 39816 19456
rect 39304 19440 39356 19446
rect 39304 19382 39356 19388
rect 38844 18420 38896 18426
rect 38844 18362 38896 18368
rect 39316 18222 39344 19382
rect 39580 19372 39632 19378
rect 39580 19314 39632 19320
rect 39592 18698 39620 19314
rect 40144 19174 40172 19858
rect 40328 19854 40356 21354
rect 40604 21146 40632 21490
rect 40592 21140 40644 21146
rect 40592 21082 40644 21088
rect 40408 21072 40460 21078
rect 40408 21014 40460 21020
rect 40420 20466 40448 21014
rect 42720 20874 42748 21490
rect 42708 20868 42760 20874
rect 42708 20810 42760 20816
rect 42524 20800 42576 20806
rect 42524 20742 42576 20748
rect 40408 20460 40460 20466
rect 40408 20402 40460 20408
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 40132 19168 40184 19174
rect 40132 19110 40184 19116
rect 41236 19168 41288 19174
rect 41236 19110 41288 19116
rect 40684 18760 40736 18766
rect 40684 18702 40736 18708
rect 39580 18692 39632 18698
rect 39580 18634 39632 18640
rect 39592 18290 39620 18634
rect 40696 18290 40724 18702
rect 41248 18358 41276 19110
rect 41236 18352 41288 18358
rect 41236 18294 41288 18300
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 40040 18284 40092 18290
rect 40040 18226 40092 18232
rect 40684 18284 40736 18290
rect 40684 18226 40736 18232
rect 39304 18216 39356 18222
rect 39304 18158 39356 18164
rect 40052 17678 40080 18226
rect 40316 18080 40368 18086
rect 40316 18022 40368 18028
rect 40328 17678 40356 18022
rect 41432 17882 41460 19994
rect 42536 19854 42564 20742
rect 42720 20602 42748 20810
rect 42800 20800 42852 20806
rect 42800 20742 42852 20748
rect 42708 20596 42760 20602
rect 42708 20538 42760 20544
rect 42708 20460 42760 20466
rect 42708 20402 42760 20408
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 42524 19848 42576 19854
rect 42524 19790 42576 19796
rect 41524 18766 41552 19790
rect 41604 19780 41656 19786
rect 41604 19722 41656 19728
rect 41616 19514 41644 19722
rect 41696 19712 41748 19718
rect 41696 19654 41748 19660
rect 41708 19514 41736 19654
rect 41604 19508 41656 19514
rect 41604 19450 41656 19456
rect 41696 19508 41748 19514
rect 41696 19450 41748 19456
rect 41512 18760 41564 18766
rect 41512 18702 41564 18708
rect 41420 17876 41472 17882
rect 41420 17818 41472 17824
rect 40040 17672 40092 17678
rect 40040 17614 40092 17620
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 38200 17196 38252 17202
rect 38200 17138 38252 17144
rect 41524 16658 41552 18702
rect 41616 18426 41644 19450
rect 42720 19446 42748 20402
rect 42812 20398 42840 20742
rect 42800 20392 42852 20398
rect 42800 20334 42852 20340
rect 42812 20058 42840 20334
rect 42984 20324 43036 20330
rect 42984 20266 43036 20272
rect 42800 20052 42852 20058
rect 42800 19994 42852 20000
rect 42996 19514 43024 20266
rect 42892 19508 42944 19514
rect 42892 19450 42944 19456
rect 42984 19508 43036 19514
rect 42984 19450 43036 19456
rect 42708 19440 42760 19446
rect 42708 19382 42760 19388
rect 42720 19242 42748 19382
rect 42708 19236 42760 19242
rect 42708 19178 42760 19184
rect 42616 19168 42668 19174
rect 42616 19110 42668 19116
rect 42628 18766 42656 19110
rect 42616 18760 42668 18766
rect 42616 18702 42668 18708
rect 42800 18692 42852 18698
rect 42800 18634 42852 18640
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 42812 17678 42840 18634
rect 42904 18290 42932 19450
rect 42996 18970 43024 19450
rect 42984 18964 43036 18970
rect 42984 18906 43036 18912
rect 42892 18284 42944 18290
rect 42892 18226 42944 18232
rect 42800 17672 42852 17678
rect 42800 17614 42852 17620
rect 38200 16652 38252 16658
rect 38200 16594 38252 16600
rect 38384 16652 38436 16658
rect 38384 16594 38436 16600
rect 41512 16652 41564 16658
rect 41512 16594 41564 16600
rect 38212 16250 38240 16594
rect 38200 16244 38252 16250
rect 38200 16186 38252 16192
rect 38212 15366 38240 16186
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38304 15026 38332 16050
rect 38016 15020 38068 15026
rect 38016 14962 38068 14968
rect 38292 15020 38344 15026
rect 38292 14962 38344 14968
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 38304 13326 38332 14962
rect 38396 14006 38424 16594
rect 38476 16516 38528 16522
rect 38476 16458 38528 16464
rect 40500 16516 40552 16522
rect 40500 16458 40552 16464
rect 38488 16046 38516 16458
rect 40132 16448 40184 16454
rect 40132 16390 40184 16396
rect 40144 16114 40172 16390
rect 40512 16250 40540 16458
rect 40500 16244 40552 16250
rect 40500 16186 40552 16192
rect 40132 16108 40184 16114
rect 40132 16050 40184 16056
rect 38476 16040 38528 16046
rect 38476 15982 38528 15988
rect 38660 16040 38712 16046
rect 38660 15982 38712 15988
rect 38844 16040 38896 16046
rect 38844 15982 38896 15988
rect 38488 15706 38516 15982
rect 38476 15700 38528 15706
rect 38476 15642 38528 15648
rect 38672 15026 38700 15982
rect 38660 15020 38712 15026
rect 38660 14962 38712 14968
rect 38476 14952 38528 14958
rect 38476 14894 38528 14900
rect 38488 14074 38516 14894
rect 38476 14068 38528 14074
rect 38476 14010 38528 14016
rect 38384 14000 38436 14006
rect 38384 13942 38436 13948
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38304 12850 38332 13262
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 37568 11150 37596 12174
rect 38292 11824 38344 11830
rect 38292 11766 38344 11772
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 11150 37872 11494
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37568 10674 37596 11086
rect 38304 10742 38332 11766
rect 38396 11694 38424 13942
rect 38672 13462 38700 14962
rect 38856 14482 38884 15982
rect 39120 15088 39172 15094
rect 39120 15030 39172 15036
rect 38844 14476 38896 14482
rect 38844 14418 38896 14424
rect 38856 13462 38884 14418
rect 39132 14414 39160 15030
rect 39488 15020 39540 15026
rect 39488 14962 39540 14968
rect 39500 14618 39528 14962
rect 39764 14952 39816 14958
rect 39764 14894 39816 14900
rect 39488 14612 39540 14618
rect 39488 14554 39540 14560
rect 39776 14414 39804 14894
rect 39120 14408 39172 14414
rect 39120 14350 39172 14356
rect 39764 14408 39816 14414
rect 39764 14350 39816 14356
rect 38660 13456 38712 13462
rect 38660 13398 38712 13404
rect 38844 13456 38896 13462
rect 38844 13398 38896 13404
rect 38672 12850 38700 13398
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38476 12776 38528 12782
rect 38476 12718 38528 12724
rect 38488 11762 38516 12718
rect 38476 11756 38528 11762
rect 38476 11698 38528 11704
rect 38384 11688 38436 11694
rect 38384 11630 38436 11636
rect 38488 11354 38516 11698
rect 38476 11348 38528 11354
rect 38476 11290 38528 11296
rect 38292 10736 38344 10742
rect 38292 10678 38344 10684
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 10266 37872 10610
rect 37832 10260 37884 10266
rect 37832 10202 37884 10208
rect 38304 10130 38332 10678
rect 38856 10130 38884 13398
rect 38936 12844 38988 12850
rect 38936 12786 38988 12792
rect 38948 10810 38976 12786
rect 39776 12782 39804 14350
rect 39948 14340 40000 14346
rect 39948 14282 40000 14288
rect 40408 14340 40460 14346
rect 40408 14282 40460 14288
rect 39960 14006 39988 14282
rect 40420 14074 40448 14282
rect 41420 14272 41472 14278
rect 41420 14214 41472 14220
rect 40408 14068 40460 14074
rect 40408 14010 40460 14016
rect 41432 14006 41460 14214
rect 39948 14000 40000 14006
rect 39948 13942 40000 13948
rect 41420 14000 41472 14006
rect 41420 13942 41472 13948
rect 40224 13796 40276 13802
rect 40224 13738 40276 13744
rect 39948 13252 40000 13258
rect 39948 13194 40000 13200
rect 40132 13252 40184 13258
rect 40132 13194 40184 13200
rect 39764 12776 39816 12782
rect 39764 12718 39816 12724
rect 39776 12238 39804 12718
rect 39960 12442 39988 13194
rect 40040 13184 40092 13190
rect 40040 13126 40092 13132
rect 40052 12918 40080 13126
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39948 12436 40000 12442
rect 39948 12378 40000 12384
rect 39764 12232 39816 12238
rect 39764 12174 39816 12180
rect 39960 11898 39988 12378
rect 40144 12170 40172 13194
rect 40132 12164 40184 12170
rect 40132 12106 40184 12112
rect 39948 11892 40000 11898
rect 39948 11834 40000 11840
rect 40144 11830 40172 12106
rect 40132 11824 40184 11830
rect 40132 11766 40184 11772
rect 40236 11694 40264 13738
rect 41144 13320 41196 13326
rect 41144 13262 41196 13268
rect 41156 12986 41184 13262
rect 41144 12980 41196 12986
rect 41144 12922 41196 12928
rect 40592 12164 40644 12170
rect 40592 12106 40644 12112
rect 40604 11898 40632 12106
rect 40592 11892 40644 11898
rect 40592 11834 40644 11840
rect 40224 11688 40276 11694
rect 40224 11630 40276 11636
rect 38936 10804 38988 10810
rect 38936 10746 38988 10752
rect 38292 10124 38344 10130
rect 38292 10066 38344 10072
rect 38844 10124 38896 10130
rect 38844 10066 38896 10072
rect 38948 10062 38976 10746
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 43088 6914 43116 23258
rect 43272 23186 43300 24686
rect 43994 24647 44050 24656
rect 43996 23656 44048 23662
rect 43996 23598 44048 23604
rect 44008 23225 44036 23598
rect 43994 23216 44050 23225
rect 43260 23180 43312 23186
rect 43994 23151 44050 23160
rect 43260 23122 43312 23128
rect 43168 22976 43220 22982
rect 43168 22918 43220 22924
rect 43180 22234 43208 22918
rect 43168 22228 43220 22234
rect 43168 22170 43220 22176
rect 43166 21720 43222 21729
rect 43166 21655 43222 21664
rect 43180 21622 43208 21655
rect 43168 21616 43220 21622
rect 43168 21558 43220 21564
rect 43272 21010 43300 23122
rect 43260 21004 43312 21010
rect 43260 20946 43312 20952
rect 43168 20392 43220 20398
rect 43168 20334 43220 20340
rect 43180 20233 43208 20334
rect 43166 20224 43222 20233
rect 43166 20159 43222 20168
rect 43272 19310 43300 20946
rect 43260 19304 43312 19310
rect 43260 19246 43312 19252
rect 43166 18728 43222 18737
rect 43166 18663 43222 18672
rect 43180 18358 43208 18663
rect 43168 18352 43220 18358
rect 43168 18294 43220 18300
rect 43168 17604 43220 17610
rect 43168 17546 43220 17552
rect 43180 17241 43208 17546
rect 43166 17232 43222 17241
rect 43166 17167 43222 17176
rect 43352 15904 43404 15910
rect 43352 15846 43404 15852
rect 43364 15745 43392 15846
rect 43350 15736 43406 15745
rect 43350 15671 43406 15680
rect 43352 14408 43404 14414
rect 43352 14350 43404 14356
rect 43364 14249 43392 14350
rect 43350 14240 43406 14249
rect 43350 14175 43406 14184
rect 43168 12776 43220 12782
rect 43166 12744 43168 12753
rect 43220 12744 43222 12753
rect 43166 12679 43222 12688
rect 43168 11688 43220 11694
rect 43168 11630 43220 11636
rect 43180 11257 43208 11630
rect 43166 11248 43222 11257
rect 43166 11183 43222 11192
rect 43168 9988 43220 9994
rect 43168 9930 43220 9936
rect 43180 9761 43208 9930
rect 43166 9752 43222 9761
rect 43166 9687 43222 9696
rect 43996 8424 44048 8430
rect 43996 8366 44048 8372
rect 44008 8265 44036 8366
rect 43994 8256 44050 8265
rect 43994 8191 44050 8200
rect 42812 6886 43116 6914
rect 42812 5710 42840 6886
rect 43166 6760 43222 6769
rect 43166 6695 43168 6704
rect 43220 6695 43222 6704
rect 43168 6666 43220 6672
rect 42800 5704 42852 5710
rect 42800 5646 42852 5652
rect 43996 5636 44048 5642
rect 43996 5578 44048 5584
rect 44008 5273 44036 5578
rect 43994 5264 44050 5273
rect 43994 5199 44050 5208
rect 37004 4140 37056 4146
rect 37004 4082 37056 4088
rect 43168 4072 43220 4078
rect 43168 4014 43220 4020
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 43180 3777 43208 4014
rect 43166 3768 43222 3777
rect 43166 3703 43222 3712
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 43168 2372 43220 2378
rect 43168 2314 43220 2320
rect 43180 2281 43208 2314
rect 43166 2272 43222 2281
rect 19574 2204 19882 2213
rect 43166 2207 43222 2216
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
<< via2 >>
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 7194 40024 7250 40080
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 5538 36216 5594 36272
rect 5538 35980 5540 36000
rect 5540 35980 5592 36000
rect 5592 35980 5594 36000
rect 5538 35944 5594 35980
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 5538 35128 5594 35184
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 10322 39888 10378 39944
rect 10690 39924 10692 39944
rect 10692 39924 10744 39944
rect 10744 39924 10746 39944
rect 10690 39888 10746 39924
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 10322 37204 10324 37224
rect 10324 37204 10376 37224
rect 10376 37204 10378 37224
rect 10322 37168 10378 37204
rect 10874 36352 10930 36408
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 12346 36624 12402 36680
rect 13450 37304 13506 37360
rect 12622 36624 12678 36680
rect 11518 29844 11574 29880
rect 11518 29824 11520 29844
rect 11520 29824 11572 29844
rect 11572 29824 11574 29844
rect 13358 37168 13414 37224
rect 13634 36624 13690 36680
rect 13358 35128 13414 35184
rect 13174 34040 13230 34096
rect 16486 38392 16542 38448
rect 15474 36624 15530 36680
rect 15658 36352 15714 36408
rect 16302 36624 16358 36680
rect 17038 37188 17094 37224
rect 17038 37168 17040 37188
rect 17040 37168 17092 37188
rect 17092 37168 17094 37188
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 18694 39344 18750 39400
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 18326 38392 18382 38448
rect 17590 35944 17646 36000
rect 17222 29180 17224 29200
rect 17224 29180 17276 29200
rect 17276 29180 17278 29200
rect 17222 29144 17278 29180
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 16946 26444 17002 26480
rect 16946 26424 16948 26444
rect 16948 26424 17000 26444
rect 17000 26424 17002 26444
rect 17222 26968 17278 27024
rect 18878 38392 18934 38448
rect 19798 38528 19854 38584
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19154 37304 19210 37360
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 18510 36216 18566 36272
rect 17774 26424 17830 26480
rect 18418 26424 18474 26480
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 18786 29844 18842 29880
rect 18786 29824 18788 29844
rect 18788 29824 18840 29844
rect 18840 29824 18842 29844
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 20994 38528 21050 38584
rect 22558 37984 22614 38040
rect 22098 36780 22154 36816
rect 22098 36760 22100 36780
rect 22100 36760 22152 36780
rect 22152 36760 22154 36780
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 18602 26288 18658 26344
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 22006 35944 22062 36000
rect 22742 37712 22798 37768
rect 22190 35944 22246 36000
rect 21914 32272 21970 32328
rect 23110 38936 23166 38992
rect 24122 40704 24178 40760
rect 21270 30252 21326 30288
rect 21270 30232 21272 30252
rect 21272 30232 21324 30252
rect 21324 30232 21326 30252
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20810 27376 20866 27432
rect 21270 27124 21326 27160
rect 21270 27104 21272 27124
rect 21272 27104 21324 27124
rect 21324 27104 21326 27124
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 21362 26832 21418 26888
rect 21638 27104 21694 27160
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 22466 23160 22522 23216
rect 23294 31764 23296 31784
rect 23296 31764 23348 31784
rect 23348 31764 23350 31784
rect 23294 31728 23350 31764
rect 23202 29552 23258 29608
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 26238 41248 26294 41304
rect 25134 35708 25136 35728
rect 25136 35708 25188 35728
rect 25188 35708 25190 35728
rect 25134 35672 25190 35708
rect 26238 39208 26294 39264
rect 25410 36760 25466 36816
rect 25962 33924 26018 33960
rect 25962 33904 25964 33924
rect 25964 33904 26016 33924
rect 26016 33904 26018 33924
rect 26422 33652 26478 33688
rect 26422 33632 26424 33652
rect 26424 33632 26476 33652
rect 26476 33632 26478 33652
rect 27250 39208 27306 39264
rect 27618 40160 27674 40216
rect 28446 41112 28502 41168
rect 28906 41248 28962 41304
rect 28722 41112 28778 41168
rect 28630 40976 28686 41032
rect 28814 41012 28816 41032
rect 28816 41012 28868 41032
rect 28868 41012 28870 41032
rect 28446 40704 28502 40760
rect 28354 40024 28410 40080
rect 26882 36236 26938 36272
rect 26882 36216 26884 36236
rect 26884 36216 26936 36236
rect 26936 36216 26938 36236
rect 26330 31728 26386 31784
rect 25686 27396 25742 27432
rect 25686 27376 25688 27396
rect 25688 27376 25740 27396
rect 25740 27376 25742 27396
rect 25410 26832 25466 26888
rect 24490 24132 24546 24168
rect 24490 24112 24492 24132
rect 24492 24112 24544 24132
rect 24544 24112 24546 24132
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 27710 36624 27766 36680
rect 28354 38392 28410 38448
rect 27986 35672 28042 35728
rect 28170 34740 28226 34776
rect 28170 34720 28172 34740
rect 28172 34720 28224 34740
rect 28224 34720 28226 34740
rect 27802 33260 27804 33280
rect 27804 33260 27856 33280
rect 27856 33260 27858 33280
rect 27802 33224 27858 33260
rect 28538 37848 28594 37904
rect 28814 40976 28870 41012
rect 28906 40724 28962 40760
rect 28906 40704 28908 40724
rect 28908 40704 28960 40724
rect 28960 40704 28962 40724
rect 28814 39924 28816 39944
rect 28816 39924 28868 39944
rect 28868 39924 28870 39944
rect 28814 39888 28870 39924
rect 28906 38936 28962 38992
rect 28078 30252 28134 30288
rect 28538 34448 28594 34504
rect 28446 33652 28502 33688
rect 28446 33632 28448 33652
rect 28448 33632 28500 33652
rect 28500 33632 28502 33652
rect 28446 33224 28502 33280
rect 28630 33088 28686 33144
rect 29642 38392 29698 38448
rect 30194 40160 30250 40216
rect 32586 41384 32642 41440
rect 29458 37168 29514 37224
rect 29090 37032 29146 37088
rect 28814 32272 28870 32328
rect 28078 30232 28080 30252
rect 28080 30232 28132 30252
rect 28132 30232 28134 30252
rect 27342 25472 27398 25528
rect 27526 25472 27582 25528
rect 28630 28464 28686 28520
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 28262 27512 28318 27568
rect 27894 26188 27896 26208
rect 27896 26188 27948 26208
rect 27948 26188 27950 26208
rect 27894 26152 27950 26188
rect 28538 24148 28540 24168
rect 28540 24148 28592 24168
rect 28592 24148 28594 24168
rect 28538 24112 28594 24148
rect 29090 26968 29146 27024
rect 32034 37204 32036 37224
rect 32036 37204 32088 37224
rect 32088 37204 32090 37224
rect 32034 37168 32090 37204
rect 32402 37712 32458 37768
rect 31482 34740 31538 34776
rect 31482 34720 31484 34740
rect 31484 34720 31536 34740
rect 31536 34720 31538 34740
rect 31022 33904 31078 33960
rect 31022 31184 31078 31240
rect 30746 29552 30802 29608
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 29918 20848 29974 20904
rect 30102 20304 30158 20360
rect 30286 26308 30342 26344
rect 30286 26288 30288 26308
rect 30288 26288 30340 26308
rect 30340 26288 30342 26308
rect 30470 26424 30526 26480
rect 31114 29688 31170 29744
rect 31298 29144 31354 29200
rect 31758 30504 31814 30560
rect 31758 29688 31814 29744
rect 32494 32544 32550 32600
rect 30746 25916 30748 25936
rect 30748 25916 30800 25936
rect 30800 25916 30802 25936
rect 30746 25880 30802 25916
rect 31390 29008 31446 29064
rect 30930 21956 30986 21992
rect 30930 21936 30932 21956
rect 30932 21936 30984 21956
rect 30984 21936 30986 21956
rect 30378 19896 30434 19952
rect 31666 28872 31722 28928
rect 31850 28484 31906 28520
rect 31850 28464 31852 28484
rect 31852 28464 31904 28484
rect 31904 28464 31906 28484
rect 31850 27512 31906 27568
rect 31206 21664 31262 21720
rect 31574 19352 31630 19408
rect 31850 26988 31906 27024
rect 31850 26968 31852 26988
rect 31852 26968 31904 26988
rect 31904 26968 31906 26988
rect 32034 27376 32090 27432
rect 32402 30096 32458 30152
rect 33046 37032 33102 37088
rect 33138 33088 33194 33144
rect 33782 39888 33838 39944
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34150 37848 34206 37904
rect 33874 37204 33876 37224
rect 33876 37204 33928 37224
rect 33928 37204 33930 37224
rect 33874 37168 33930 37204
rect 33874 34448 33930 34504
rect 33414 30368 33470 30424
rect 33138 29688 33194 29744
rect 33138 29008 33194 29064
rect 32586 27920 32642 27976
rect 32126 20984 32182 21040
rect 31850 19796 31852 19816
rect 31852 19796 31904 19816
rect 31904 19796 31906 19816
rect 31850 19760 31906 19796
rect 32586 26560 32642 26616
rect 32862 24812 32918 24848
rect 32862 24792 32864 24812
rect 32864 24792 32916 24812
rect 32916 24792 32918 24812
rect 33138 26832 33194 26888
rect 33414 29588 33416 29608
rect 33416 29588 33468 29608
rect 33468 29588 33470 29608
rect 33414 29552 33470 29588
rect 33506 27376 33562 27432
rect 33230 21936 33286 21992
rect 31758 19352 31814 19408
rect 33414 17856 33470 17912
rect 33782 33904 33838 33960
rect 33782 33768 33838 33824
rect 34150 31476 34206 31512
rect 34150 31456 34152 31476
rect 34152 31456 34204 31476
rect 34204 31456 34206 31476
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34518 30368 34574 30424
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36910 39344 36966 39400
rect 35530 38700 35532 38720
rect 35532 38700 35584 38720
rect 35584 38700 35586 38720
rect 35530 38664 35586 38700
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35070 36216 35126 36272
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35254 32272 35310 32328
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35254 31864 35310 31920
rect 35162 31764 35164 31784
rect 35164 31764 35216 31784
rect 35216 31764 35218 31784
rect 35162 31728 35218 31764
rect 35438 31220 35440 31240
rect 35440 31220 35492 31240
rect 35492 31220 35494 31240
rect 35438 31184 35494 31220
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34886 30096 34942 30152
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34702 29144 34758 29200
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34150 25880 34206 25936
rect 34518 26288 34574 26344
rect 34426 25900 34482 25936
rect 34426 25880 34428 25900
rect 34428 25880 34480 25900
rect 34480 25880 34482 25900
rect 34058 23724 34114 23760
rect 34058 23704 34060 23724
rect 34060 23704 34112 23724
rect 34112 23704 34114 23724
rect 34334 20576 34390 20632
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35898 37304 35954 37360
rect 35898 35028 35900 35048
rect 35900 35028 35952 35048
rect 35952 35028 35954 35048
rect 35898 34992 35954 35028
rect 35714 31900 35716 31920
rect 35716 31900 35768 31920
rect 35768 31900 35770 31920
rect 35714 31864 35770 31900
rect 36174 34584 36230 34640
rect 36174 33768 36230 33824
rect 35990 31764 35992 31784
rect 35992 31764 36044 31784
rect 36044 31764 36046 31784
rect 35990 31728 36046 31764
rect 36450 35028 36452 35048
rect 36452 35028 36504 35048
rect 36504 35028 36506 35048
rect 36450 34992 36506 35028
rect 37186 39208 37242 39264
rect 36910 37304 36966 37360
rect 35714 30252 35770 30288
rect 35714 30232 35716 30252
rect 35716 30232 35768 30252
rect 35768 30232 35770 30252
rect 35714 26288 35770 26344
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 36450 30096 36506 30152
rect 36634 27512 36690 27568
rect 36542 26832 36598 26888
rect 37094 34448 37150 34504
rect 36910 26968 36966 27024
rect 37370 35028 37372 35048
rect 37372 35028 37424 35048
rect 37424 35028 37426 35048
rect 37370 34992 37426 35028
rect 37462 30796 37518 30832
rect 37462 30776 37464 30796
rect 37464 30776 37516 30796
rect 37516 30776 37518 30796
rect 37278 30504 37334 30560
rect 37554 29688 37610 29744
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34978 21936 35034 21992
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35438 20884 35440 20904
rect 35440 20884 35492 20904
rect 35492 20884 35494 20904
rect 35438 20848 35494 20884
rect 35254 20460 35310 20496
rect 35254 20440 35256 20460
rect 35256 20440 35308 20460
rect 35308 20440 35310 20460
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37922 31340 37978 31376
rect 37922 31320 37924 31340
rect 37924 31320 37976 31340
rect 37976 31320 37978 31340
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38290 31592 38346 31648
rect 38290 31184 38346 31240
rect 38566 31592 38622 31648
rect 38474 31456 38530 31512
rect 38290 29008 38346 29064
rect 37830 21004 37886 21040
rect 37830 20984 37832 21004
rect 37832 20984 37884 21004
rect 37884 20984 37886 21004
rect 37186 19896 37242 19952
rect 43994 42608 44050 42664
rect 38658 26832 38714 26888
rect 38842 24248 38898 24304
rect 38934 24012 38936 24032
rect 38936 24012 38988 24032
rect 38988 24012 38990 24032
rect 38934 23976 38990 24012
rect 39026 23432 39082 23488
rect 39210 23976 39266 24032
rect 39762 35944 39818 36000
rect 43994 41112 44050 41168
rect 43994 39616 44050 39672
rect 43994 38120 44050 38176
rect 43994 36624 44050 36680
rect 43994 35148 44050 35184
rect 43994 35128 43996 35148
rect 43996 35128 44048 35148
rect 44048 35128 44050 35148
rect 43994 33632 44050 33688
rect 43166 32136 43222 32192
rect 43166 30640 43222 30696
rect 43166 29144 43222 29200
rect 38934 20304 38990 20360
rect 39118 19760 39174 19816
rect 43994 27648 44050 27704
rect 43166 26152 43222 26208
rect 43994 24656 44050 24712
rect 43994 23160 44050 23216
rect 43166 21664 43222 21720
rect 43166 20168 43222 20224
rect 43166 18672 43222 18728
rect 43166 17176 43222 17232
rect 43350 15680 43406 15736
rect 43350 14184 43406 14240
rect 43166 12724 43168 12744
rect 43168 12724 43220 12744
rect 43220 12724 43222 12744
rect 43166 12688 43222 12724
rect 43166 11192 43222 11248
rect 43166 9696 43222 9752
rect 43994 8200 44050 8256
rect 43166 6724 43222 6760
rect 43166 6704 43168 6724
rect 43168 6704 43220 6724
rect 43220 6704 43222 6724
rect 43994 5208 44050 5264
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 43166 3712 43222 3768
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 43166 2216 43222 2272
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 43989 42666 44055 42669
rect 44200 42666 45000 42696
rect 43989 42664 45000 42666
rect 43989 42608 43994 42664
rect 44050 42608 45000 42664
rect 43989 42606 45000 42608
rect 43989 42603 44055 42606
rect 44200 42576 45000 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 32581 41442 32647 41445
rect 32806 41442 32812 41444
rect 32581 41440 32812 41442
rect 32581 41384 32586 41440
rect 32642 41384 32812 41440
rect 32581 41382 32812 41384
rect 32581 41379 32647 41382
rect 32806 41380 32812 41382
rect 32876 41380 32882 41444
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 26233 41306 26299 41309
rect 28901 41306 28967 41309
rect 26233 41304 28967 41306
rect 26233 41248 26238 41304
rect 26294 41248 28906 41304
rect 28962 41248 28967 41304
rect 26233 41246 28967 41248
rect 26233 41243 26299 41246
rect 28901 41243 28967 41246
rect 28441 41170 28507 41173
rect 28717 41170 28783 41173
rect 28441 41168 28783 41170
rect 28441 41112 28446 41168
rect 28502 41112 28722 41168
rect 28778 41112 28783 41168
rect 28441 41110 28783 41112
rect 28441 41107 28507 41110
rect 28717 41107 28783 41110
rect 43989 41170 44055 41173
rect 44200 41170 45000 41200
rect 43989 41168 45000 41170
rect 43989 41112 43994 41168
rect 44050 41112 45000 41168
rect 43989 41110 45000 41112
rect 43989 41107 44055 41110
rect 44200 41080 45000 41110
rect 28625 41034 28691 41037
rect 28809 41034 28875 41037
rect 28625 41032 28875 41034
rect 28625 40976 28630 41032
rect 28686 40976 28814 41032
rect 28870 40976 28875 41032
rect 28625 40974 28875 40976
rect 28625 40971 28691 40974
rect 28809 40971 28875 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 24117 40762 24183 40765
rect 28441 40762 28507 40765
rect 28901 40762 28967 40765
rect 24117 40760 28967 40762
rect 24117 40704 24122 40760
rect 24178 40704 28446 40760
rect 28502 40704 28906 40760
rect 28962 40704 28967 40760
rect 24117 40702 28967 40704
rect 24117 40699 24183 40702
rect 28441 40699 28507 40702
rect 28901 40699 28967 40702
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 27613 40218 27679 40221
rect 30189 40218 30255 40221
rect 27613 40216 30255 40218
rect 27613 40160 27618 40216
rect 27674 40160 30194 40216
rect 30250 40160 30255 40216
rect 27613 40158 30255 40160
rect 27613 40155 27679 40158
rect 30189 40155 30255 40158
rect 7189 40082 7255 40085
rect 8150 40082 8156 40084
rect 7189 40080 8156 40082
rect 7189 40024 7194 40080
rect 7250 40024 8156 40080
rect 7189 40022 8156 40024
rect 7189 40019 7255 40022
rect 8150 40020 8156 40022
rect 8220 40020 8226 40084
rect 28349 40082 28415 40085
rect 28349 40080 28458 40082
rect 28349 40024 28354 40080
rect 28410 40024 28458 40080
rect 28349 40019 28458 40024
rect 10317 39946 10383 39949
rect 10685 39946 10751 39949
rect 10910 39946 10916 39948
rect 10317 39944 10916 39946
rect 10317 39888 10322 39944
rect 10378 39888 10690 39944
rect 10746 39888 10916 39944
rect 10317 39886 10916 39888
rect 10317 39883 10383 39886
rect 10685 39883 10751 39886
rect 10910 39884 10916 39886
rect 10980 39884 10986 39948
rect 28398 39946 28458 40019
rect 28809 39948 28875 39949
rect 28758 39946 28764 39948
rect 28398 39886 28764 39946
rect 28828 39944 28875 39948
rect 28870 39888 28875 39944
rect 28758 39884 28764 39886
rect 28828 39884 28875 39888
rect 28942 39884 28948 39948
rect 29012 39946 29018 39948
rect 33777 39946 33843 39949
rect 29012 39944 33843 39946
rect 29012 39888 33782 39944
rect 33838 39888 33843 39944
rect 29012 39886 33843 39888
rect 29012 39884 29018 39886
rect 28809 39883 28875 39884
rect 33777 39883 33843 39886
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 43989 39674 44055 39677
rect 44200 39674 45000 39704
rect 43989 39672 45000 39674
rect 43989 39616 43994 39672
rect 44050 39616 45000 39672
rect 43989 39614 45000 39616
rect 43989 39611 44055 39614
rect 44200 39584 45000 39614
rect 18689 39402 18755 39405
rect 32622 39402 32628 39404
rect 18689 39400 32628 39402
rect 18689 39344 18694 39400
rect 18750 39344 32628 39400
rect 18689 39342 32628 39344
rect 18689 39339 18755 39342
rect 32622 39340 32628 39342
rect 32692 39402 32698 39404
rect 36905 39402 36971 39405
rect 32692 39400 36971 39402
rect 32692 39344 36910 39400
rect 36966 39344 36971 39400
rect 32692 39342 36971 39344
rect 32692 39340 32698 39342
rect 36905 39339 36971 39342
rect 26233 39266 26299 39269
rect 27245 39266 27311 39269
rect 27470 39266 27476 39268
rect 26233 39264 27476 39266
rect 26233 39208 26238 39264
rect 26294 39208 27250 39264
rect 27306 39208 27476 39264
rect 26233 39206 27476 39208
rect 26233 39203 26299 39206
rect 27245 39203 27311 39206
rect 27470 39204 27476 39206
rect 27540 39204 27546 39268
rect 36670 39204 36676 39268
rect 36740 39266 36746 39268
rect 37181 39266 37247 39269
rect 36740 39264 37247 39266
rect 36740 39208 37186 39264
rect 37242 39208 37247 39264
rect 36740 39206 37247 39208
rect 36740 39204 36746 39206
rect 37181 39203 37247 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 23105 38994 23171 38997
rect 28901 38994 28967 38997
rect 23105 38992 28967 38994
rect 23105 38936 23110 38992
rect 23166 38936 28906 38992
rect 28962 38936 28967 38992
rect 23105 38934 28967 38936
rect 23105 38931 23171 38934
rect 28901 38931 28967 38934
rect 35525 38724 35591 38725
rect 35525 38720 35572 38724
rect 35636 38722 35642 38724
rect 35525 38664 35530 38720
rect 35525 38660 35572 38664
rect 35636 38662 35682 38722
rect 35636 38660 35642 38662
rect 35525 38659 35591 38660
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19793 38586 19859 38589
rect 20989 38586 21055 38589
rect 19793 38584 21055 38586
rect 19793 38528 19798 38584
rect 19854 38528 20994 38584
rect 21050 38528 21055 38584
rect 19793 38526 21055 38528
rect 19793 38523 19859 38526
rect 20989 38523 21055 38526
rect 16481 38450 16547 38453
rect 18321 38450 18387 38453
rect 16481 38448 18387 38450
rect 16481 38392 16486 38448
rect 16542 38392 18326 38448
rect 18382 38392 18387 38448
rect 16481 38390 18387 38392
rect 16481 38387 16547 38390
rect 18321 38387 18387 38390
rect 18873 38450 18939 38453
rect 28349 38450 28415 38453
rect 29637 38450 29703 38453
rect 18873 38448 29703 38450
rect 18873 38392 18878 38448
rect 18934 38392 28354 38448
rect 28410 38392 29642 38448
rect 29698 38392 29703 38448
rect 18873 38390 29703 38392
rect 18873 38387 18939 38390
rect 28349 38387 28415 38390
rect 29637 38387 29703 38390
rect 43989 38178 44055 38181
rect 44200 38178 45000 38208
rect 43989 38176 45000 38178
rect 43989 38120 43994 38176
rect 44050 38120 45000 38176
rect 43989 38118 45000 38120
rect 43989 38115 44055 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 44200 38088 45000 38118
rect 19570 38047 19886 38048
rect 22553 38042 22619 38045
rect 22553 38040 31770 38042
rect 22553 37984 22558 38040
rect 22614 37984 31770 38040
rect 22553 37982 31770 37984
rect 22553 37979 22619 37982
rect 28533 37908 28599 37909
rect 28533 37906 28580 37908
rect 28488 37904 28580 37906
rect 28488 37848 28538 37904
rect 28488 37846 28580 37848
rect 28533 37844 28580 37846
rect 28644 37844 28650 37908
rect 31710 37906 31770 37982
rect 34145 37906 34211 37909
rect 31710 37904 34211 37906
rect 31710 37848 34150 37904
rect 34206 37848 34211 37904
rect 31710 37846 34211 37848
rect 28533 37843 28599 37844
rect 34145 37843 34211 37846
rect 22737 37770 22803 37773
rect 32397 37770 32463 37773
rect 22737 37768 32463 37770
rect 22737 37712 22742 37768
rect 22798 37712 32402 37768
rect 32458 37712 32463 37768
rect 22737 37710 32463 37712
rect 22737 37707 22803 37710
rect 32397 37707 32463 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 13445 37362 13511 37365
rect 19149 37362 19215 37365
rect 13445 37360 19215 37362
rect 13445 37304 13450 37360
rect 13506 37304 19154 37360
rect 19210 37304 19215 37360
rect 13445 37302 19215 37304
rect 13445 37299 13511 37302
rect 19149 37299 19215 37302
rect 31886 37300 31892 37364
rect 31956 37362 31962 37364
rect 35893 37362 35959 37365
rect 36905 37362 36971 37365
rect 31956 37360 36971 37362
rect 31956 37304 35898 37360
rect 35954 37304 36910 37360
rect 36966 37304 36971 37360
rect 31956 37302 36971 37304
rect 31956 37300 31962 37302
rect 35893 37299 35959 37302
rect 36905 37299 36971 37302
rect 10317 37226 10383 37229
rect 13353 37226 13419 37229
rect 10317 37224 13419 37226
rect 10317 37168 10322 37224
rect 10378 37168 13358 37224
rect 13414 37168 13419 37224
rect 10317 37166 13419 37168
rect 10317 37163 10383 37166
rect 13353 37163 13419 37166
rect 17033 37226 17099 37229
rect 29453 37226 29519 37229
rect 17033 37224 29519 37226
rect 17033 37168 17038 37224
rect 17094 37168 29458 37224
rect 29514 37168 29519 37224
rect 17033 37166 29519 37168
rect 17033 37163 17099 37166
rect 29453 37163 29519 37166
rect 32029 37226 32095 37229
rect 33869 37226 33935 37229
rect 32029 37224 33935 37226
rect 32029 37168 32034 37224
rect 32090 37168 33874 37224
rect 33930 37168 33935 37224
rect 32029 37166 33935 37168
rect 32029 37163 32095 37166
rect 33869 37163 33935 37166
rect 29085 37090 29151 37093
rect 33041 37090 33107 37093
rect 29085 37088 33107 37090
rect 29085 37032 29090 37088
rect 29146 37032 33046 37088
rect 33102 37032 33107 37088
rect 29085 37030 33107 37032
rect 29085 37027 29151 37030
rect 33041 37027 33107 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 22093 36818 22159 36821
rect 25405 36818 25471 36821
rect 22093 36816 25471 36818
rect 22093 36760 22098 36816
rect 22154 36760 25410 36816
rect 25466 36760 25471 36816
rect 22093 36758 25471 36760
rect 22093 36755 22159 36758
rect 25405 36755 25471 36758
rect 12341 36682 12407 36685
rect 12617 36682 12683 36685
rect 12341 36680 12683 36682
rect 12341 36624 12346 36680
rect 12402 36624 12622 36680
rect 12678 36624 12683 36680
rect 12341 36622 12683 36624
rect 12341 36619 12407 36622
rect 12617 36619 12683 36622
rect 13629 36682 13695 36685
rect 15469 36682 15535 36685
rect 13629 36680 15535 36682
rect 13629 36624 13634 36680
rect 13690 36624 15474 36680
rect 15530 36624 15535 36680
rect 13629 36622 15535 36624
rect 13629 36619 13695 36622
rect 15469 36619 15535 36622
rect 16297 36682 16363 36685
rect 27705 36682 27771 36685
rect 16297 36680 27771 36682
rect 16297 36624 16302 36680
rect 16358 36624 27710 36680
rect 27766 36624 27771 36680
rect 16297 36622 27771 36624
rect 16297 36619 16363 36622
rect 27705 36619 27771 36622
rect 43989 36682 44055 36685
rect 44200 36682 45000 36712
rect 43989 36680 45000 36682
rect 43989 36624 43994 36680
rect 44050 36624 45000 36680
rect 43989 36622 45000 36624
rect 43989 36619 44055 36622
rect 44200 36592 45000 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 10869 36410 10935 36413
rect 15653 36410 15719 36413
rect 10869 36408 15719 36410
rect 10869 36352 10874 36408
rect 10930 36352 15658 36408
rect 15714 36352 15719 36408
rect 10869 36350 15719 36352
rect 10869 36347 10935 36350
rect 15653 36347 15719 36350
rect 5533 36274 5599 36277
rect 18505 36274 18571 36277
rect 5533 36272 18571 36274
rect 5533 36216 5538 36272
rect 5594 36216 18510 36272
rect 18566 36216 18571 36272
rect 5533 36214 18571 36216
rect 5533 36211 5599 36214
rect 18505 36211 18571 36214
rect 26877 36274 26943 36277
rect 35065 36274 35131 36277
rect 26877 36272 35131 36274
rect 26877 36216 26882 36272
rect 26938 36216 35070 36272
rect 35126 36216 35131 36272
rect 26877 36214 35131 36216
rect 26877 36211 26943 36214
rect 35065 36211 35131 36214
rect 5533 36002 5599 36005
rect 17585 36002 17651 36005
rect 5533 36000 17651 36002
rect 5533 35944 5538 36000
rect 5594 35944 17590 36000
rect 17646 35944 17651 36000
rect 5533 35942 17651 35944
rect 5533 35939 5599 35942
rect 17585 35939 17651 35942
rect 22001 36002 22067 36005
rect 22185 36002 22251 36005
rect 22001 36000 22251 36002
rect 22001 35944 22006 36000
rect 22062 35944 22190 36000
rect 22246 35944 22251 36000
rect 22001 35942 22251 35944
rect 22001 35939 22067 35942
rect 22185 35939 22251 35942
rect 39062 35940 39068 36004
rect 39132 36002 39138 36004
rect 39757 36002 39823 36005
rect 39132 36000 39823 36002
rect 39132 35944 39762 36000
rect 39818 35944 39823 36000
rect 39132 35942 39823 35944
rect 39132 35940 39138 35942
rect 39757 35939 39823 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 25129 35730 25195 35733
rect 27981 35730 28047 35733
rect 25129 35728 28047 35730
rect 25129 35672 25134 35728
rect 25190 35672 27986 35728
rect 28042 35672 28047 35728
rect 25129 35670 28047 35672
rect 25129 35667 25195 35670
rect 27981 35667 28047 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 5533 35186 5599 35189
rect 13353 35186 13419 35189
rect 5533 35184 13419 35186
rect 5533 35128 5538 35184
rect 5594 35128 13358 35184
rect 13414 35128 13419 35184
rect 5533 35126 13419 35128
rect 5533 35123 5599 35126
rect 13353 35123 13419 35126
rect 43989 35186 44055 35189
rect 44200 35186 45000 35216
rect 43989 35184 45000 35186
rect 43989 35128 43994 35184
rect 44050 35128 45000 35184
rect 43989 35126 45000 35128
rect 43989 35123 44055 35126
rect 44200 35096 45000 35126
rect 35893 35052 35959 35053
rect 35893 35050 35940 35052
rect 35848 35048 35940 35050
rect 35848 34992 35898 35048
rect 35848 34990 35940 34992
rect 35893 34988 35940 34990
rect 36004 34988 36010 35052
rect 36445 35050 36511 35053
rect 37365 35050 37431 35053
rect 36445 35048 37431 35050
rect 36445 34992 36450 35048
rect 36506 34992 37370 35048
rect 37426 34992 37431 35048
rect 36445 34990 37431 34992
rect 35893 34987 35959 34988
rect 36445 34987 36511 34990
rect 37365 34987 37431 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 28165 34778 28231 34781
rect 31477 34778 31543 34781
rect 28165 34776 31543 34778
rect 28165 34720 28170 34776
rect 28226 34720 31482 34776
rect 31538 34720 31543 34776
rect 28165 34718 31543 34720
rect 28165 34715 28231 34718
rect 31477 34715 31543 34718
rect 36169 34642 36235 34645
rect 36126 34640 36235 34642
rect 36126 34584 36174 34640
rect 36230 34584 36235 34640
rect 36126 34579 36235 34584
rect 28533 34506 28599 34509
rect 28942 34506 28948 34508
rect 28533 34504 28948 34506
rect 28533 34448 28538 34504
rect 28594 34448 28948 34504
rect 28533 34446 28948 34448
rect 28533 34443 28599 34446
rect 28942 34444 28948 34446
rect 29012 34444 29018 34508
rect 33869 34506 33935 34509
rect 36126 34506 36186 34579
rect 37089 34506 37155 34509
rect 33869 34504 37155 34506
rect 33869 34448 33874 34504
rect 33930 34448 37094 34504
rect 37150 34448 37155 34504
rect 33869 34446 37155 34448
rect 33869 34443 33935 34446
rect 37089 34443 37155 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 13169 34098 13235 34101
rect 27654 34098 27660 34100
rect 13169 34096 27660 34098
rect 13169 34040 13174 34096
rect 13230 34040 27660 34096
rect 13169 34038 27660 34040
rect 13169 34035 13235 34038
rect 27654 34036 27660 34038
rect 27724 34036 27730 34100
rect 25957 33962 26023 33965
rect 31017 33962 31083 33965
rect 33777 33962 33843 33965
rect 25957 33960 33843 33962
rect 25957 33904 25962 33960
rect 26018 33904 31022 33960
rect 31078 33904 33782 33960
rect 33838 33904 33843 33960
rect 25957 33902 33843 33904
rect 25957 33899 26023 33902
rect 31017 33899 31083 33902
rect 33777 33899 33843 33902
rect 33777 33826 33843 33829
rect 36169 33826 36235 33829
rect 33777 33824 36235 33826
rect 33777 33768 33782 33824
rect 33838 33768 36174 33824
rect 36230 33768 36235 33824
rect 33777 33766 36235 33768
rect 33777 33763 33843 33766
rect 36169 33763 36235 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 26417 33690 26483 33693
rect 28441 33690 28507 33693
rect 26417 33688 28507 33690
rect 26417 33632 26422 33688
rect 26478 33632 28446 33688
rect 28502 33632 28507 33688
rect 26417 33630 28507 33632
rect 26417 33627 26483 33630
rect 28441 33627 28507 33630
rect 43989 33690 44055 33693
rect 44200 33690 45000 33720
rect 43989 33688 45000 33690
rect 43989 33632 43994 33688
rect 44050 33632 45000 33688
rect 43989 33630 45000 33632
rect 43989 33627 44055 33630
rect 44200 33600 45000 33630
rect 27797 33282 27863 33285
rect 28441 33282 28507 33285
rect 27797 33280 28507 33282
rect 27797 33224 27802 33280
rect 27858 33224 28446 33280
rect 28502 33224 28507 33280
rect 27797 33222 28507 33224
rect 27797 33219 27863 33222
rect 28441 33219 28507 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 28625 33148 28691 33149
rect 28574 33146 28580 33148
rect 28534 33086 28580 33146
rect 28644 33144 28691 33148
rect 28686 33088 28691 33144
rect 28574 33084 28580 33086
rect 28644 33084 28691 33088
rect 32806 33084 32812 33148
rect 32876 33146 32882 33148
rect 33133 33146 33199 33149
rect 32876 33144 33199 33146
rect 32876 33088 33138 33144
rect 33194 33088 33199 33144
rect 32876 33086 33199 33088
rect 32876 33084 32882 33086
rect 28625 33083 28691 33084
rect 33133 33083 33199 33086
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 27654 32540 27660 32604
rect 27724 32602 27730 32604
rect 32489 32602 32555 32605
rect 27724 32600 32555 32602
rect 27724 32544 32494 32600
rect 32550 32544 32555 32600
rect 27724 32542 32555 32544
rect 27724 32540 27730 32542
rect 32489 32539 32555 32542
rect 21909 32330 21975 32333
rect 28809 32330 28875 32333
rect 21909 32328 28875 32330
rect 21909 32272 21914 32328
rect 21970 32272 28814 32328
rect 28870 32272 28875 32328
rect 21909 32270 28875 32272
rect 21909 32267 21975 32270
rect 28809 32267 28875 32270
rect 35249 32330 35315 32333
rect 35249 32328 35450 32330
rect 35249 32272 35254 32328
rect 35310 32272 35450 32328
rect 35249 32270 35450 32272
rect 35249 32267 35315 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 35249 31922 35315 31925
rect 35390 31922 35450 32270
rect 43161 32194 43227 32197
rect 44200 32194 45000 32224
rect 43161 32192 45000 32194
rect 43161 32136 43166 32192
rect 43222 32136 45000 32192
rect 43161 32134 45000 32136
rect 43161 32131 43227 32134
rect 44200 32104 45000 32134
rect 35709 31924 35775 31925
rect 35709 31922 35756 31924
rect 35249 31920 35450 31922
rect 35249 31864 35254 31920
rect 35310 31864 35450 31920
rect 35249 31862 35450 31864
rect 35664 31920 35756 31922
rect 35664 31864 35714 31920
rect 35664 31862 35756 31864
rect 35249 31859 35315 31862
rect 35709 31860 35756 31862
rect 35820 31860 35826 31924
rect 35709 31859 35775 31860
rect 23289 31786 23355 31789
rect 26325 31786 26391 31789
rect 23289 31784 26391 31786
rect 23289 31728 23294 31784
rect 23350 31728 26330 31784
rect 26386 31728 26391 31784
rect 23289 31726 26391 31728
rect 23289 31723 23355 31726
rect 26325 31723 26391 31726
rect 35157 31786 35223 31789
rect 35985 31786 36051 31789
rect 35157 31784 36051 31786
rect 35157 31728 35162 31784
rect 35218 31728 35990 31784
rect 36046 31728 36051 31784
rect 35157 31726 36051 31728
rect 35157 31723 35223 31726
rect 35985 31723 36051 31726
rect 38285 31650 38351 31653
rect 38561 31650 38627 31653
rect 38285 31648 38627 31650
rect 38285 31592 38290 31648
rect 38346 31592 38566 31648
rect 38622 31592 38627 31648
rect 38285 31590 38627 31592
rect 38285 31587 38351 31590
rect 38561 31587 38627 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 34145 31514 34211 31517
rect 38469 31514 38535 31517
rect 34145 31512 38535 31514
rect 34145 31456 34150 31512
rect 34206 31456 38474 31512
rect 38530 31456 38535 31512
rect 34145 31454 38535 31456
rect 34145 31451 34211 31454
rect 38469 31451 38535 31454
rect 37917 31378 37983 31381
rect 37917 31376 38026 31378
rect 37917 31320 37922 31376
rect 37978 31320 38026 31376
rect 37917 31315 38026 31320
rect 31017 31242 31083 31245
rect 35433 31242 35499 31245
rect 31017 31240 35499 31242
rect 31017 31184 31022 31240
rect 31078 31184 35438 31240
rect 35494 31184 35499 31240
rect 31017 31182 35499 31184
rect 37966 31242 38026 31315
rect 38285 31242 38351 31245
rect 37966 31240 38351 31242
rect 37966 31184 38290 31240
rect 38346 31184 38351 31240
rect 37966 31182 38351 31184
rect 31017 31179 31083 31182
rect 35433 31179 35499 31182
rect 38285 31179 38351 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 31518 30772 31524 30836
rect 31588 30834 31594 30836
rect 37457 30834 37523 30837
rect 31588 30832 37523 30834
rect 31588 30776 37462 30832
rect 37518 30776 37523 30832
rect 31588 30774 37523 30776
rect 31588 30772 31594 30774
rect 37457 30771 37523 30774
rect 43161 30698 43227 30701
rect 44200 30698 45000 30728
rect 43161 30696 45000 30698
rect 43161 30640 43166 30696
rect 43222 30640 45000 30696
rect 43161 30638 45000 30640
rect 43161 30635 43227 30638
rect 44200 30608 45000 30638
rect 31753 30562 31819 30565
rect 37273 30562 37339 30565
rect 31753 30560 37339 30562
rect 31753 30504 31758 30560
rect 31814 30504 37278 30560
rect 37334 30504 37339 30560
rect 31753 30502 37339 30504
rect 31753 30499 31819 30502
rect 37273 30499 37339 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 33409 30426 33475 30429
rect 33542 30426 33548 30428
rect 33409 30424 33548 30426
rect 33409 30368 33414 30424
rect 33470 30368 33548 30424
rect 33409 30366 33548 30368
rect 33409 30363 33475 30366
rect 33542 30364 33548 30366
rect 33612 30364 33618 30428
rect 34278 30364 34284 30428
rect 34348 30426 34354 30428
rect 34513 30426 34579 30429
rect 34348 30424 34579 30426
rect 34348 30368 34518 30424
rect 34574 30368 34579 30424
rect 34348 30366 34579 30368
rect 34348 30364 34354 30366
rect 34513 30363 34579 30366
rect 21265 30290 21331 30293
rect 28073 30290 28139 30293
rect 21265 30288 28139 30290
rect 21265 30232 21270 30288
rect 21326 30232 28078 30288
rect 28134 30232 28139 30288
rect 21265 30230 28139 30232
rect 21265 30227 21331 30230
rect 28073 30227 28139 30230
rect 35709 30292 35775 30293
rect 35709 30288 35756 30292
rect 35820 30290 35826 30292
rect 35709 30232 35714 30288
rect 35709 30228 35756 30232
rect 35820 30230 35866 30290
rect 35820 30228 35826 30230
rect 35709 30227 35775 30228
rect 32397 30154 32463 30157
rect 34881 30154 34947 30157
rect 36445 30154 36511 30157
rect 32397 30152 36511 30154
rect 32397 30096 32402 30152
rect 32458 30096 34886 30152
rect 34942 30096 36450 30152
rect 36506 30096 36511 30152
rect 32397 30094 36511 30096
rect 32397 30091 32463 30094
rect 34881 30091 34947 30094
rect 36445 30091 36511 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 11513 29882 11579 29885
rect 18781 29882 18847 29885
rect 11513 29880 18847 29882
rect 11513 29824 11518 29880
rect 11574 29824 18786 29880
rect 18842 29824 18847 29880
rect 11513 29822 18847 29824
rect 11513 29819 11579 29822
rect 18781 29819 18847 29822
rect 31109 29746 31175 29749
rect 31334 29746 31340 29748
rect 31109 29744 31340 29746
rect 31109 29688 31114 29744
rect 31170 29688 31340 29744
rect 31109 29686 31340 29688
rect 31109 29683 31175 29686
rect 31334 29684 31340 29686
rect 31404 29746 31410 29748
rect 31753 29746 31819 29749
rect 31404 29744 31819 29746
rect 31404 29688 31758 29744
rect 31814 29688 31819 29744
rect 31404 29686 31819 29688
rect 31404 29684 31410 29686
rect 31753 29683 31819 29686
rect 33133 29746 33199 29749
rect 37549 29746 37615 29749
rect 33133 29744 37615 29746
rect 33133 29688 33138 29744
rect 33194 29688 37554 29744
rect 37610 29688 37615 29744
rect 33133 29686 37615 29688
rect 33133 29683 33199 29686
rect 37549 29683 37615 29686
rect 10910 29548 10916 29612
rect 10980 29610 10986 29612
rect 23197 29610 23263 29613
rect 10980 29608 23263 29610
rect 10980 29552 23202 29608
rect 23258 29552 23263 29608
rect 10980 29550 23263 29552
rect 10980 29548 10986 29550
rect 23197 29547 23263 29550
rect 30741 29610 30807 29613
rect 33409 29610 33475 29613
rect 30741 29608 33475 29610
rect 30741 29552 30746 29608
rect 30802 29552 33414 29608
rect 33470 29552 33475 29608
rect 30741 29550 33475 29552
rect 30741 29547 30807 29550
rect 33409 29547 33475 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 8150 29140 8156 29204
rect 8220 29202 8226 29204
rect 17217 29202 17283 29205
rect 8220 29200 17283 29202
rect 8220 29144 17222 29200
rect 17278 29144 17283 29200
rect 8220 29142 17283 29144
rect 8220 29140 8226 29142
rect 17217 29139 17283 29142
rect 31293 29202 31359 29205
rect 34697 29202 34763 29205
rect 31293 29200 34763 29202
rect 31293 29144 31298 29200
rect 31354 29144 34702 29200
rect 34758 29144 34763 29200
rect 31293 29142 34763 29144
rect 31293 29139 31359 29142
rect 34697 29139 34763 29142
rect 43161 29202 43227 29205
rect 44200 29202 45000 29232
rect 43161 29200 45000 29202
rect 43161 29144 43166 29200
rect 43222 29144 45000 29200
rect 43161 29142 45000 29144
rect 43161 29139 43227 29142
rect 44200 29112 45000 29142
rect 31385 29066 31451 29069
rect 33133 29066 33199 29069
rect 38285 29066 38351 29069
rect 31385 29064 38351 29066
rect 31385 29008 31390 29064
rect 31446 29008 33138 29064
rect 33194 29008 38290 29064
rect 38346 29008 38351 29064
rect 31385 29006 38351 29008
rect 31385 29003 31451 29006
rect 33133 29003 33199 29006
rect 38285 29003 38351 29006
rect 31661 28932 31727 28933
rect 31661 28930 31708 28932
rect 31616 28928 31708 28930
rect 31616 28872 31666 28928
rect 31616 28870 31708 28872
rect 31661 28868 31708 28870
rect 31772 28868 31778 28932
rect 31661 28867 31727 28868
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 28625 28522 28691 28525
rect 28758 28522 28764 28524
rect 28625 28520 28764 28522
rect 28625 28464 28630 28520
rect 28686 28464 28764 28520
rect 28625 28462 28764 28464
rect 28625 28459 28691 28462
rect 28758 28460 28764 28462
rect 28828 28460 28834 28524
rect 31518 28460 31524 28524
rect 31588 28522 31594 28524
rect 31845 28522 31911 28525
rect 31588 28520 31911 28522
rect 31588 28464 31850 28520
rect 31906 28464 31911 28520
rect 31588 28462 31911 28464
rect 31588 28460 31594 28462
rect 31845 28459 31911 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 32581 27980 32647 27981
rect 32581 27978 32628 27980
rect 32536 27976 32628 27978
rect 32536 27920 32586 27976
rect 32536 27918 32628 27920
rect 32581 27916 32628 27918
rect 32692 27916 32698 27980
rect 32581 27915 32647 27916
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 43989 27706 44055 27709
rect 44200 27706 45000 27736
rect 43989 27704 45000 27706
rect 43989 27648 43994 27704
rect 44050 27648 45000 27704
rect 43989 27646 45000 27648
rect 43989 27643 44055 27646
rect 44200 27616 45000 27646
rect 28257 27570 28323 27573
rect 31845 27570 31911 27573
rect 28257 27568 31911 27570
rect 28257 27512 28262 27568
rect 28318 27512 31850 27568
rect 31906 27512 31911 27568
rect 28257 27510 31911 27512
rect 28257 27507 28323 27510
rect 31845 27507 31911 27510
rect 36629 27572 36695 27573
rect 36629 27568 36676 27572
rect 36740 27570 36746 27572
rect 36629 27512 36634 27568
rect 36629 27508 36676 27512
rect 36740 27510 36786 27570
rect 36740 27508 36746 27510
rect 36629 27507 36695 27508
rect 20805 27434 20871 27437
rect 25681 27434 25747 27437
rect 32029 27434 32095 27437
rect 33501 27434 33567 27437
rect 20805 27432 33567 27434
rect 20805 27376 20810 27432
rect 20866 27376 25686 27432
rect 25742 27376 32034 27432
rect 32090 27376 33506 27432
rect 33562 27376 33567 27432
rect 20805 27374 33567 27376
rect 20805 27371 20871 27374
rect 25681 27371 25747 27374
rect 32029 27371 32095 27374
rect 33501 27371 33567 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 21265 27162 21331 27165
rect 21633 27162 21699 27165
rect 21265 27160 21699 27162
rect 21265 27104 21270 27160
rect 21326 27104 21638 27160
rect 21694 27104 21699 27160
rect 21265 27102 21699 27104
rect 21265 27099 21331 27102
rect 21633 27099 21699 27102
rect 17217 27026 17283 27029
rect 29085 27026 29151 27029
rect 31845 27026 31911 27029
rect 36905 27026 36971 27029
rect 17217 27024 31770 27026
rect 17217 26968 17222 27024
rect 17278 26968 29090 27024
rect 29146 26968 31770 27024
rect 17217 26966 31770 26968
rect 17217 26963 17283 26966
rect 29085 26963 29151 26966
rect 21357 26890 21423 26893
rect 25405 26890 25471 26893
rect 21357 26888 25471 26890
rect 21357 26832 21362 26888
rect 21418 26832 25410 26888
rect 25466 26832 25471 26888
rect 21357 26830 25471 26832
rect 21357 26827 21423 26830
rect 25405 26827 25471 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 31710 26618 31770 26966
rect 31845 27024 36971 27026
rect 31845 26968 31850 27024
rect 31906 26968 36910 27024
rect 36966 26968 36971 27024
rect 31845 26966 36971 26968
rect 31845 26963 31911 26966
rect 36905 26963 36971 26966
rect 33133 26890 33199 26893
rect 36537 26890 36603 26893
rect 33133 26888 36603 26890
rect 33133 26832 33138 26888
rect 33194 26832 36542 26888
rect 36598 26832 36603 26888
rect 33133 26830 36603 26832
rect 33133 26827 33199 26830
rect 36537 26827 36603 26830
rect 38653 26892 38719 26893
rect 38653 26888 38700 26892
rect 38764 26890 38770 26892
rect 38653 26832 38658 26888
rect 38653 26828 38700 26832
rect 38764 26830 38810 26890
rect 38764 26828 38770 26830
rect 38653 26827 38719 26828
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 32581 26618 32647 26621
rect 31710 26616 32647 26618
rect 31710 26560 32586 26616
rect 32642 26560 32647 26616
rect 31710 26558 32647 26560
rect 32581 26555 32647 26558
rect 16941 26482 17007 26485
rect 17769 26482 17835 26485
rect 18413 26482 18479 26485
rect 30465 26484 30531 26485
rect 30414 26482 30420 26484
rect 16941 26480 18479 26482
rect 16941 26424 16946 26480
rect 17002 26424 17774 26480
rect 17830 26424 18418 26480
rect 18474 26424 18479 26480
rect 16941 26422 18479 26424
rect 30374 26422 30420 26482
rect 30484 26480 30531 26484
rect 30526 26424 30531 26480
rect 16941 26419 17007 26422
rect 17769 26419 17835 26422
rect 18413 26419 18479 26422
rect 30414 26420 30420 26422
rect 30484 26420 30531 26424
rect 30465 26419 30531 26420
rect 18597 26346 18663 26349
rect 24894 26346 24900 26348
rect 18597 26344 24900 26346
rect 18597 26288 18602 26344
rect 18658 26288 24900 26344
rect 18597 26286 24900 26288
rect 18597 26283 18663 26286
rect 24894 26284 24900 26286
rect 24964 26284 24970 26348
rect 30281 26346 30347 26349
rect 34513 26346 34579 26349
rect 35709 26346 35775 26349
rect 30281 26344 35775 26346
rect 30281 26288 30286 26344
rect 30342 26288 34518 26344
rect 34574 26288 35714 26344
rect 35770 26288 35775 26344
rect 30281 26286 35775 26288
rect 30281 26283 30347 26286
rect 34513 26283 34579 26286
rect 35709 26283 35775 26286
rect 27470 26148 27476 26212
rect 27540 26210 27546 26212
rect 27889 26210 27955 26213
rect 27540 26208 27955 26210
rect 27540 26152 27894 26208
rect 27950 26152 27955 26208
rect 27540 26150 27955 26152
rect 27540 26148 27546 26150
rect 27889 26147 27955 26150
rect 43161 26210 43227 26213
rect 44200 26210 45000 26240
rect 43161 26208 45000 26210
rect 43161 26152 43166 26208
rect 43222 26152 45000 26208
rect 43161 26150 45000 26152
rect 43161 26147 43227 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 44200 26120 45000 26150
rect 19570 26079 19886 26080
rect 30741 25938 30807 25941
rect 34145 25938 34211 25941
rect 34421 25938 34487 25941
rect 30741 25936 34487 25938
rect 30741 25880 30746 25936
rect 30802 25880 34150 25936
rect 34206 25880 34426 25936
rect 34482 25880 34487 25936
rect 30741 25878 34487 25880
rect 30741 25875 30807 25878
rect 34145 25875 34211 25878
rect 34421 25875 34487 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 27337 25530 27403 25533
rect 27521 25530 27587 25533
rect 27337 25528 27587 25530
rect 27337 25472 27342 25528
rect 27398 25472 27526 25528
rect 27582 25472 27587 25528
rect 27337 25470 27587 25472
rect 27337 25467 27403 25470
rect 27521 25467 27587 25470
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 32857 24850 32923 24853
rect 35934 24850 35940 24852
rect 32857 24848 35940 24850
rect 32857 24792 32862 24848
rect 32918 24792 35940 24848
rect 32857 24790 35940 24792
rect 32857 24787 32923 24790
rect 35934 24788 35940 24790
rect 36004 24788 36010 24852
rect 43989 24714 44055 24717
rect 44200 24714 45000 24744
rect 43989 24712 45000 24714
rect 43989 24656 43994 24712
rect 44050 24656 45000 24712
rect 43989 24654 45000 24656
rect 43989 24651 44055 24654
rect 44200 24624 45000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 38694 24244 38700 24308
rect 38764 24306 38770 24308
rect 38837 24306 38903 24309
rect 38764 24304 38903 24306
rect 38764 24248 38842 24304
rect 38898 24248 38903 24304
rect 38764 24246 38903 24248
rect 38764 24244 38770 24246
rect 38837 24243 38903 24246
rect 24485 24170 24551 24173
rect 28533 24170 28599 24173
rect 24485 24168 28599 24170
rect 24485 24112 24490 24168
rect 24546 24112 28538 24168
rect 28594 24112 28599 24168
rect 24485 24110 28599 24112
rect 24485 24107 24551 24110
rect 28533 24107 28599 24110
rect 38929 24034 38995 24037
rect 39205 24034 39271 24037
rect 38929 24032 39271 24034
rect 38929 23976 38934 24032
rect 38990 23976 39210 24032
rect 39266 23976 39271 24032
rect 38929 23974 39271 23976
rect 38929 23971 38995 23974
rect 39205 23971 39271 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 24894 23700 24900 23764
rect 24964 23762 24970 23764
rect 34053 23762 34119 23765
rect 24964 23760 34119 23762
rect 24964 23704 34058 23760
rect 34114 23704 34119 23760
rect 24964 23702 34119 23704
rect 24964 23700 24970 23702
rect 34053 23699 34119 23702
rect 39021 23492 39087 23493
rect 39021 23488 39068 23492
rect 39132 23490 39138 23492
rect 39021 23432 39026 23488
rect 39021 23428 39068 23432
rect 39132 23430 39178 23490
rect 39132 23428 39138 23430
rect 39021 23427 39087 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 22461 23218 22527 23221
rect 30414 23218 30420 23220
rect 22461 23216 30420 23218
rect 22461 23160 22466 23216
rect 22522 23160 30420 23216
rect 22461 23158 30420 23160
rect 22461 23155 22527 23158
rect 30414 23156 30420 23158
rect 30484 23156 30490 23220
rect 43989 23218 44055 23221
rect 44200 23218 45000 23248
rect 43989 23216 45000 23218
rect 43989 23160 43994 23216
rect 44050 23160 45000 23216
rect 43989 23158 45000 23160
rect 43989 23155 44055 23158
rect 44200 23128 45000 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 30925 21994 30991 21997
rect 33225 21994 33291 21997
rect 34973 21994 35039 21997
rect 30925 21992 35039 21994
rect 30925 21936 30930 21992
rect 30986 21936 33230 21992
rect 33286 21936 34978 21992
rect 35034 21936 35039 21992
rect 30925 21934 35039 21936
rect 30925 21931 30991 21934
rect 33225 21931 33291 21934
rect 34973 21931 35039 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 31201 21722 31267 21725
rect 32622 21722 32628 21724
rect 31201 21720 32628 21722
rect 31201 21664 31206 21720
rect 31262 21664 32628 21720
rect 31201 21662 32628 21664
rect 31201 21659 31267 21662
rect 32622 21660 32628 21662
rect 32692 21660 32698 21724
rect 43161 21722 43227 21725
rect 44200 21722 45000 21752
rect 43161 21720 45000 21722
rect 43161 21664 43166 21720
rect 43222 21664 45000 21720
rect 43161 21662 45000 21664
rect 43161 21659 43227 21662
rect 44200 21632 45000 21662
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 32121 21042 32187 21045
rect 37825 21042 37891 21045
rect 32121 21040 37891 21042
rect 32121 20984 32126 21040
rect 32182 20984 37830 21040
rect 37886 20984 37891 21040
rect 32121 20982 37891 20984
rect 32121 20979 32187 20982
rect 37825 20979 37891 20982
rect 29913 20906 29979 20909
rect 35433 20906 35499 20909
rect 29913 20904 35499 20906
rect 29913 20848 29918 20904
rect 29974 20848 35438 20904
rect 35494 20848 35499 20904
rect 29913 20846 35499 20848
rect 29913 20843 29979 20846
rect 35433 20843 35499 20846
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 34329 20636 34395 20637
rect 34278 20634 34284 20636
rect 34238 20574 34284 20634
rect 34348 20632 34395 20636
rect 34390 20576 34395 20632
rect 34278 20572 34284 20574
rect 34348 20572 34395 20576
rect 34329 20571 34395 20572
rect 35249 20498 35315 20501
rect 35566 20498 35572 20500
rect 35249 20496 35572 20498
rect 35249 20440 35254 20496
rect 35310 20440 35572 20496
rect 35249 20438 35572 20440
rect 35249 20435 35315 20438
rect 35566 20436 35572 20438
rect 35636 20436 35642 20500
rect 30097 20362 30163 20365
rect 38929 20362 38995 20365
rect 30097 20360 38995 20362
rect 30097 20304 30102 20360
rect 30158 20304 38934 20360
rect 38990 20304 38995 20360
rect 30097 20302 38995 20304
rect 30097 20299 30163 20302
rect 38929 20299 38995 20302
rect 43161 20226 43227 20229
rect 44200 20226 45000 20256
rect 43161 20224 45000 20226
rect 43161 20168 43166 20224
rect 43222 20168 45000 20224
rect 43161 20166 45000 20168
rect 43161 20163 43227 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 44200 20136 45000 20166
rect 34930 20095 35246 20096
rect 30373 19954 30439 19957
rect 31518 19954 31524 19956
rect 30373 19952 31524 19954
rect 30373 19896 30378 19952
rect 30434 19896 31524 19952
rect 30373 19894 31524 19896
rect 30373 19891 30439 19894
rect 31518 19892 31524 19894
rect 31588 19954 31594 19956
rect 37181 19954 37247 19957
rect 31588 19952 37247 19954
rect 31588 19896 37186 19952
rect 37242 19896 37247 19952
rect 31588 19894 37247 19896
rect 31588 19892 31594 19894
rect 37181 19891 37247 19894
rect 31845 19818 31911 19821
rect 39113 19818 39179 19821
rect 31845 19816 39179 19818
rect 31845 19760 31850 19816
rect 31906 19760 39118 19816
rect 39174 19760 39179 19816
rect 31845 19758 39179 19760
rect 31845 19755 31911 19758
rect 39113 19755 39179 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 31569 19410 31635 19413
rect 31753 19410 31819 19413
rect 31569 19408 31854 19410
rect 31569 19352 31574 19408
rect 31630 19352 31758 19408
rect 31814 19352 31854 19408
rect 31569 19350 31854 19352
rect 31569 19347 31635 19350
rect 31753 19347 31819 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 43161 18730 43227 18733
rect 44200 18730 45000 18760
rect 43161 18728 45000 18730
rect 43161 18672 43166 18728
rect 43222 18672 45000 18728
rect 43161 18670 45000 18672
rect 43161 18667 43227 18670
rect 44200 18640 45000 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 33409 17914 33475 17917
rect 33542 17914 33548 17916
rect 33409 17912 33548 17914
rect 33409 17856 33414 17912
rect 33470 17856 33548 17912
rect 33409 17854 33548 17856
rect 33409 17851 33475 17854
rect 33542 17852 33548 17854
rect 33612 17852 33618 17916
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 43161 17234 43227 17237
rect 44200 17234 45000 17264
rect 43161 17232 45000 17234
rect 43161 17176 43166 17232
rect 43222 17176 45000 17232
rect 43161 17174 45000 17176
rect 43161 17171 43227 17174
rect 44200 17144 45000 17174
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 43345 15738 43411 15741
rect 44200 15738 45000 15768
rect 43345 15736 45000 15738
rect 43345 15680 43350 15736
rect 43406 15680 45000 15736
rect 43345 15678 45000 15680
rect 43345 15675 43411 15678
rect 44200 15648 45000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 43345 14242 43411 14245
rect 44200 14242 45000 14272
rect 43345 14240 45000 14242
rect 43345 14184 43350 14240
rect 43406 14184 45000 14240
rect 43345 14182 45000 14184
rect 43345 14179 43411 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 44200 14152 45000 14182
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 43161 12746 43227 12749
rect 44200 12746 45000 12776
rect 43161 12744 45000 12746
rect 43161 12688 43166 12744
rect 43222 12688 45000 12744
rect 43161 12686 45000 12688
rect 43161 12683 43227 12686
rect 44200 12656 45000 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 43161 11250 43227 11253
rect 44200 11250 45000 11280
rect 43161 11248 45000 11250
rect 43161 11192 43166 11248
rect 43222 11192 45000 11248
rect 43161 11190 45000 11192
rect 43161 11187 43227 11190
rect 44200 11160 45000 11190
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 43161 9754 43227 9757
rect 44200 9754 45000 9784
rect 43161 9752 45000 9754
rect 43161 9696 43166 9752
rect 43222 9696 45000 9752
rect 43161 9694 45000 9696
rect 43161 9691 43227 9694
rect 44200 9664 45000 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 43989 8258 44055 8261
rect 44200 8258 45000 8288
rect 43989 8256 45000 8258
rect 43989 8200 43994 8256
rect 44050 8200 45000 8256
rect 43989 8198 45000 8200
rect 43989 8195 44055 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 44200 8168 45000 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 43161 6762 43227 6765
rect 44200 6762 45000 6792
rect 43161 6760 45000 6762
rect 43161 6704 43166 6760
rect 43222 6704 45000 6760
rect 43161 6702 45000 6704
rect 43161 6699 43227 6702
rect 44200 6672 45000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 43989 5266 44055 5269
rect 44200 5266 45000 5296
rect 43989 5264 45000 5266
rect 43989 5208 43994 5264
rect 44050 5208 45000 5264
rect 43989 5206 45000 5208
rect 43989 5203 44055 5206
rect 44200 5176 45000 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 43161 3770 43227 3773
rect 44200 3770 45000 3800
rect 43161 3768 45000 3770
rect 43161 3712 43166 3768
rect 43222 3712 45000 3768
rect 43161 3710 45000 3712
rect 43161 3707 43227 3710
rect 44200 3680 45000 3710
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 43161 2274 43227 2277
rect 44200 2274 45000 2304
rect 43161 2272 45000 2274
rect 43161 2216 43166 2272
rect 43222 2216 45000 2272
rect 43161 2214 45000 2216
rect 43161 2211 43227 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 44200 2184 45000 2214
rect 19570 2143 19886 2144
<< via3 >>
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 32812 41380 32876 41444
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 8156 40020 8220 40084
rect 10916 39884 10980 39948
rect 28764 39944 28828 39948
rect 28764 39888 28814 39944
rect 28814 39888 28828 39944
rect 28764 39884 28828 39888
rect 28948 39884 29012 39948
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 32628 39340 32692 39404
rect 27476 39204 27540 39268
rect 36676 39204 36740 39268
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 35572 38720 35636 38724
rect 35572 38664 35586 38720
rect 35586 38664 35636 38720
rect 35572 38660 35636 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 28580 37904 28644 37908
rect 28580 37848 28594 37904
rect 28594 37848 28644 37904
rect 28580 37844 28644 37848
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 31892 37300 31956 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 39068 35940 39132 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 35940 35048 36004 35052
rect 35940 34992 35954 35048
rect 35954 34992 36004 35048
rect 35940 34988 36004 34992
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 28948 34444 29012 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 27660 34036 27724 34100
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 28580 33144 28644 33148
rect 28580 33088 28630 33144
rect 28630 33088 28644 33144
rect 28580 33084 28644 33088
rect 32812 33084 32876 33148
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 27660 32540 27724 32604
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 35756 31920 35820 31924
rect 35756 31864 35770 31920
rect 35770 31864 35820 31920
rect 35756 31860 35820 31864
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 31524 30772 31588 30836
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 33548 30364 33612 30428
rect 34284 30364 34348 30428
rect 35756 30288 35820 30292
rect 35756 30232 35770 30288
rect 35770 30232 35820 30288
rect 35756 30228 35820 30232
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 31340 29684 31404 29748
rect 10916 29548 10980 29612
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 8156 29140 8220 29204
rect 31708 28928 31772 28932
rect 31708 28872 31722 28928
rect 31722 28872 31772 28928
rect 31708 28868 31772 28872
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 28764 28460 28828 28524
rect 31524 28460 31588 28524
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 32628 27976 32692 27980
rect 32628 27920 32642 27976
rect 32642 27920 32692 27976
rect 32628 27916 32692 27920
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 36676 27568 36740 27572
rect 36676 27512 36690 27568
rect 36690 27512 36740 27568
rect 36676 27508 36740 27512
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 38700 26888 38764 26892
rect 38700 26832 38714 26888
rect 38714 26832 38764 26888
rect 38700 26828 38764 26832
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 30420 26480 30484 26484
rect 30420 26424 30470 26480
rect 30470 26424 30484 26480
rect 30420 26420 30484 26424
rect 24900 26284 24964 26348
rect 27476 26148 27540 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 35940 24788 36004 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 38700 24244 38764 24308
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 24900 23700 24964 23764
rect 39068 23488 39132 23492
rect 39068 23432 39082 23488
rect 39082 23432 39132 23488
rect 39068 23428 39132 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 30420 23156 30484 23220
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 32628 21660 32692 21724
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 34284 20632 34348 20636
rect 34284 20576 34334 20632
rect 34334 20576 34348 20632
rect 34284 20572 34348 20576
rect 35572 20436 35636 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 31524 19892 31588 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 33548 17852 33612 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 41920 4528 42480
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 19568 42464 19888 42480
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 34928 41920 35248 42480
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 32811 41444 32877 41445
rect 32811 41380 32812 41444
rect 32876 41380 32877 41444
rect 32811 41379 32877 41380
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 8155 40084 8221 40085
rect 8155 40020 8156 40084
rect 8220 40020 8221 40084
rect 8155 40019 8221 40020
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 8158 29205 8218 40019
rect 10915 39948 10981 39949
rect 10915 39884 10916 39948
rect 10980 39884 10981 39948
rect 10915 39883 10981 39884
rect 10918 29613 10978 39883
rect 19568 39200 19888 40224
rect 28763 39948 28829 39949
rect 28763 39884 28764 39948
rect 28828 39884 28829 39948
rect 28763 39883 28829 39884
rect 28947 39948 29013 39949
rect 28947 39884 28948 39948
rect 29012 39884 29013 39948
rect 28947 39883 29013 39884
rect 27475 39268 27541 39269
rect 27475 39204 27476 39268
rect 27540 39204 27541 39268
rect 27475 39203 27541 39204
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 10915 29612 10981 29613
rect 10915 29548 10916 29612
rect 10980 29548 10981 29612
rect 10915 29547 10981 29548
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 8155 29204 8221 29205
rect 8155 29140 8156 29204
rect 8220 29140 8221 29204
rect 8155 29139 8221 29140
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 24899 26348 24965 26349
rect 24899 26284 24900 26348
rect 24964 26284 24965 26348
rect 24899 26283 24965 26284
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 24902 23765 24962 26283
rect 27478 26213 27538 39203
rect 28579 37908 28645 37909
rect 28579 37844 28580 37908
rect 28644 37844 28645 37908
rect 28579 37843 28645 37844
rect 27659 34100 27725 34101
rect 27659 34036 27660 34100
rect 27724 34036 27725 34100
rect 27659 34035 27725 34036
rect 27662 32605 27722 34035
rect 28582 33149 28642 37843
rect 28579 33148 28645 33149
rect 28579 33084 28580 33148
rect 28644 33084 28645 33148
rect 28579 33083 28645 33084
rect 27659 32604 27725 32605
rect 27659 32540 27660 32604
rect 27724 32540 27725 32604
rect 27659 32539 27725 32540
rect 28766 28525 28826 39883
rect 28950 34509 29010 39883
rect 32627 39404 32693 39405
rect 32627 39340 32628 39404
rect 32692 39340 32693 39404
rect 32627 39339 32693 39340
rect 31891 37364 31957 37365
rect 31891 37300 31892 37364
rect 31956 37300 31957 37364
rect 31891 37299 31957 37300
rect 28947 34508 29013 34509
rect 28947 34444 28948 34508
rect 29012 34444 29013 34508
rect 28947 34443 29013 34444
rect 31523 30836 31589 30837
rect 31523 30772 31524 30836
rect 31588 30772 31589 30836
rect 31523 30771 31589 30772
rect 31339 29748 31405 29749
rect 31339 29684 31340 29748
rect 31404 29684 31405 29748
rect 31339 29683 31405 29684
rect 28763 28524 28829 28525
rect 28763 28460 28764 28524
rect 28828 28460 28829 28524
rect 28763 28459 28829 28460
rect 30419 26484 30485 26485
rect 30419 26420 30420 26484
rect 30484 26420 30485 26484
rect 30419 26419 30485 26420
rect 27475 26212 27541 26213
rect 27475 26148 27476 26212
rect 27540 26148 27541 26212
rect 27475 26147 27541 26148
rect 24899 23764 24965 23765
rect 24899 23700 24900 23764
rect 24964 23700 24965 23764
rect 24899 23699 24965 23700
rect 30422 23221 30482 26419
rect 30419 23220 30485 23221
rect 30419 23156 30420 23220
rect 30484 23156 30485 23220
rect 30419 23155 30485 23156
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 31342 22110 31402 29683
rect 31526 28525 31586 30771
rect 31707 28932 31773 28933
rect 31707 28868 31708 28932
rect 31772 28930 31773 28932
rect 31894 28930 31954 37299
rect 31772 28870 31954 28930
rect 31772 28868 31773 28870
rect 31707 28867 31773 28868
rect 31523 28524 31589 28525
rect 31523 28460 31524 28524
rect 31588 28460 31589 28524
rect 31523 28459 31589 28460
rect 32630 27981 32690 39339
rect 32814 33149 32874 41379
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 36675 39268 36741 39269
rect 36675 39204 36676 39268
rect 36740 39204 36741 39268
rect 36675 39203 36741 39204
rect 35571 38724 35637 38725
rect 35571 38660 35572 38724
rect 35636 38660 35637 38724
rect 35571 38659 35637 38660
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 32811 33148 32877 33149
rect 32811 33084 32812 33148
rect 32876 33084 32877 33148
rect 32811 33083 32877 33084
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 33547 30428 33613 30429
rect 33547 30364 33548 30428
rect 33612 30364 33613 30428
rect 33547 30363 33613 30364
rect 34283 30428 34349 30429
rect 34283 30364 34284 30428
rect 34348 30364 34349 30428
rect 34283 30363 34349 30364
rect 32627 27980 32693 27981
rect 32627 27916 32628 27980
rect 32692 27916 32693 27980
rect 32627 27915 32693 27916
rect 31342 22050 31586 22110
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 31526 19957 31586 22050
rect 32630 21725 32690 27915
rect 32627 21724 32693 21725
rect 32627 21660 32628 21724
rect 32692 21660 32693 21724
rect 32627 21659 32693 21660
rect 31523 19956 31589 19957
rect 31523 19892 31524 19956
rect 31588 19892 31589 19956
rect 31523 19891 31589 19892
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 33550 17917 33610 30363
rect 34286 20637 34346 30363
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34283 20636 34349 20637
rect 34283 20572 34284 20636
rect 34348 20572 34349 20636
rect 34283 20571 34349 20572
rect 34928 20160 35248 21184
rect 35574 20501 35634 38659
rect 35939 35052 36005 35053
rect 35939 34988 35940 35052
rect 36004 34988 36005 35052
rect 35939 34987 36005 34988
rect 35755 31924 35821 31925
rect 35755 31860 35756 31924
rect 35820 31860 35821 31924
rect 35755 31859 35821 31860
rect 35758 30293 35818 31859
rect 35755 30292 35821 30293
rect 35755 30228 35756 30292
rect 35820 30228 35821 30292
rect 35755 30227 35821 30228
rect 35942 24853 36002 34987
rect 36678 27573 36738 39203
rect 39067 36004 39133 36005
rect 39067 35940 39068 36004
rect 39132 35940 39133 36004
rect 39067 35939 39133 35940
rect 36675 27572 36741 27573
rect 36675 27508 36676 27572
rect 36740 27508 36741 27572
rect 36675 27507 36741 27508
rect 38699 26892 38765 26893
rect 38699 26828 38700 26892
rect 38764 26828 38765 26892
rect 38699 26827 38765 26828
rect 35939 24852 36005 24853
rect 35939 24788 35940 24852
rect 36004 24788 36005 24852
rect 35939 24787 36005 24788
rect 38702 24309 38762 26827
rect 38699 24308 38765 24309
rect 38699 24244 38700 24308
rect 38764 24244 38765 24308
rect 38699 24243 38765 24244
rect 39070 23493 39130 35939
rect 39067 23492 39133 23493
rect 39067 23428 39068 23492
rect 39132 23428 39133 23492
rect 39067 23427 39133 23428
rect 35571 20500 35637 20501
rect 35571 20436 35572 20500
rect 35636 20436 35637 20500
rect 35571 20435 35637 20436
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 33547 17916 33613 17917
rect 33547 17852 33548 17916
rect 33612 17852 33613 17916
rect 33547 17851 33613 17852
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_453
timestamp 1676037725
transform 1 0 42780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_460 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43424 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_461
timestamp 1676037725
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp 1676037725
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_460
timestamp 1676037725
transform 1 0 43424 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_461
timestamp 1676037725
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_445 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_453
timestamp 1676037725
transform 1 0 42780 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_460
timestamp 1676037725
transform 1 0 43424 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_453
timestamp 1676037725
transform 1 0 42780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_460
timestamp 1676037725
transform 1 0 43424 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_461
timestamp 1676037725
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_453
timestamp 1676037725
transform 1 0 42780 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_460
timestamp 1676037725
transform 1 0 43424 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_461
timestamp 1676037725
transform 1 0 43516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1676037725
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_317
timestamp 1676037725
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_328
timestamp 1676037725
transform 1 0 31280 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_340
timestamp 1676037725
transform 1 0 32384 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_352
timestamp 1676037725
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1676037725
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_408
timestamp 1676037725
transform 1 0 38640 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_453
timestamp 1676037725
transform 1 0 42780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_460
timestamp 1676037725
transform 1 0 43424 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1676037725
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_304
timestamp 1676037725
transform 1 0 29072 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1676037725
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_354
timestamp 1676037725
transform 1 0 33672 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_366
timestamp 1676037725
transform 1 0 34776 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1676037725
transform 1 0 35880 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1676037725
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_412
timestamp 1676037725
transform 1 0 39008 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_424
timestamp 1676037725
transform 1 0 40112 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_436
timestamp 1676037725
transform 1 0 41216 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_271
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_283
timestamp 1676037725
transform 1 0 27140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_331
timestamp 1676037725
transform 1 0 31556 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_339
timestamp 1676037725
transform 1 0 32292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1676037725
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_383
timestamp 1676037725
transform 1 0 36340 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_395
timestamp 1676037725
transform 1 0 37444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1676037725
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_461
timestamp 1676037725
transform 1 0 43516 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_252
timestamp 1676037725
transform 1 0 24288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_263
timestamp 1676037725
transform 1 0 25300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1676037725
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_314
timestamp 1676037725
transform 1 0 29992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_328
timestamp 1676037725
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_360
timestamp 1676037725
transform 1 0 34224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_368
timestamp 1676037725
transform 1 0 34960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_386
timestamp 1676037725
transform 1 0 36616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_397
timestamp 1676037725
transform 1 0 37628 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_407
timestamp 1676037725
transform 1 0 38548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_419
timestamp 1676037725
transform 1 0 39652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_430
timestamp 1676037725
transform 1 0 40664 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_442
timestamp 1676037725
transform 1 0 41768 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_453
timestamp 1676037725
transform 1 0 42780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_460
timestamp 1676037725
transform 1 0 43424 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1676037725
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1676037725
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1676037725
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_296
timestamp 1676037725
transform 1 0 28336 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_332
timestamp 1676037725
transform 1 0 31648 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_344
timestamp 1676037725
transform 1 0 32752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1676037725
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_373
timestamp 1676037725
transform 1 0 35420 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_383
timestamp 1676037725
transform 1 0 36340 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_395
timestamp 1676037725
transform 1 0 37444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_407
timestamp 1676037725
transform 1 0 38548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_439
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_451
timestamp 1676037725
transform 1 0 42596 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_459
timestamp 1676037725
transform 1 0 43332 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_251
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_265
timestamp 1676037725
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_296
timestamp 1676037725
transform 1 0 28336 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_308
timestamp 1676037725
transform 1 0 29440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_316
timestamp 1676037725
transform 1 0 30176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_357
timestamp 1676037725
transform 1 0 33948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_366
timestamp 1676037725
transform 1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_370
timestamp 1676037725
transform 1 0 35144 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_379
timestamp 1676037725
transform 1 0 35972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_416
timestamp 1676037725
transform 1 0 39376 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_436
timestamp 1676037725
transform 1 0 41216 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_453
timestamp 1676037725
transform 1 0 42780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_460
timestamp 1676037725
transform 1 0 43424 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1676037725
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_266
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_288
timestamp 1676037725
transform 1 0 27600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1676037725
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_351
timestamp 1676037725
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_373
timestamp 1676037725
transform 1 0 35420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_383
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_391
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_415
timestamp 1676037725
transform 1 0 39284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_432
timestamp 1676037725
transform 1 0 40848 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_444
timestamp 1676037725
transform 1 0 41952 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_456
timestamp 1676037725
transform 1 0 43056 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1676037725
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_208
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1676037725
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1676037725
transform 1 0 24932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_270
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_292
timestamp 1676037725
transform 1 0 27968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_316
timestamp 1676037725
transform 1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_324
timestamp 1676037725
transform 1 0 30912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_343
timestamp 1676037725
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_353
timestamp 1676037725
transform 1 0 33580 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_364
timestamp 1676037725
transform 1 0 34592 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_386
timestamp 1676037725
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_428
timestamp 1676037725
transform 1 0 40480 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_440
timestamp 1676037725
transform 1 0 41584 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_185
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1676037725
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1676037725
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_271
timestamp 1676037725
transform 1 0 26036 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_279
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_286
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_294
timestamp 1676037725
transform 1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1676037725
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_355
timestamp 1676037725
transform 1 0 33764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_373
timestamp 1676037725
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_383
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_395
timestamp 1676037725
transform 1 0 37444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_407
timestamp 1676037725
transform 1 0 38548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_439
timestamp 1676037725
transform 1 0 41492 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_451
timestamp 1676037725
transform 1 0 42596 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_460
timestamp 1676037725
transform 1 0 43424 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1676037725
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_250
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_262
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_297
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_314
timestamp 1676037725
transform 1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_323
timestamp 1676037725
transform 1 0 30820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_346
timestamp 1676037725
transform 1 0 32936 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_359
timestamp 1676037725
transform 1 0 34132 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_371
timestamp 1676037725
transform 1 0 35236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_383
timestamp 1676037725
transform 1 0 36340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_416
timestamp 1676037725
transform 1 0 39376 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_436
timestamp 1676037725
transform 1 0 41216 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1676037725
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_320
timestamp 1676037725
transform 1 0 30544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_332
timestamp 1676037725
transform 1 0 31648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_351
timestamp 1676037725
transform 1 0 33396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1676037725
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_382
timestamp 1676037725
transform 1 0 36248 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_411
timestamp 1676037725
transform 1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_461
timestamp 1676037725
transform 1 0 43516 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1676037725
transform 1 0 22632 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_266
timestamp 1676037725
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_304
timestamp 1676037725
transform 1 0 29072 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_312
timestamp 1676037725
transform 1 0 29808 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_322
timestamp 1676037725
transform 1 0 30728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_345
timestamp 1676037725
transform 1 0 32844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_363
timestamp 1676037725
transform 1 0 34500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_367
timestamp 1676037725
transform 1 0 34868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1676037725
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_416
timestamp 1676037725
transform 1 0 39376 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_460
timestamp 1676037725
transform 1 0 43424 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_182
timestamp 1676037725
transform 1 0 17848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_216
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_224
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1676037725
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1676037725
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1676037725
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_274
timestamp 1676037725
transform 1 0 26312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_282
timestamp 1676037725
transform 1 0 27048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1676037725
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_322
timestamp 1676037725
transform 1 0 30728 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_347
timestamp 1676037725
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1676037725
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_373
timestamp 1676037725
transform 1 0 35420 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_383
timestamp 1676037725
transform 1 0 36340 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_408
timestamp 1676037725
transform 1 0 38640 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_440
timestamp 1676037725
transform 1 0 41584 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_452
timestamp 1676037725
transform 1 0 42688 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_460
timestamp 1676037725
transform 1 0 43424 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_188
timestamp 1676037725
transform 1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1676037725
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1676037725
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_292
timestamp 1676037725
transform 1 0 27968 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_319
timestamp 1676037725
transform 1 0 30452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_367
timestamp 1676037725
transform 1 0 34868 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_377
timestamp 1676037725
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_148
timestamp 1676037725
transform 1 0 14720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_158
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_174
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_186
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_207
timestamp 1676037725
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_219
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1676037725
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_273
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_292
timestamp 1676037725
transform 1 0 27968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_300
timestamp 1676037725
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_327
timestamp 1676037725
transform 1 0 31188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_347
timestamp 1676037725
transform 1 0 33028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1676037725
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_378
timestamp 1676037725
transform 1 0 35880 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_399
timestamp 1676037725
transform 1 0 37812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_411
timestamp 1676037725
transform 1 0 38916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_440
timestamp 1676037725
transform 1 0 41584 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_452
timestamp 1676037725
transform 1 0 42688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_460
timestamp 1676037725
transform 1 0 43424 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1676037725
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_187
timestamp 1676037725
transform 1 0 18308 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1676037725
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_240
timestamp 1676037725
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1676037725
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1676037725
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_355
timestamp 1676037725
transform 1 0 33764 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1676037725
transform 1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_377
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1676037725
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_412
timestamp 1676037725
transform 1 0 39008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_423
timestamp 1676037725
transform 1 0 40020 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1676037725
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_453
timestamp 1676037725
transform 1 0 42780 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_460
timestamp 1676037725
transform 1 0 43424 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1676037725
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_156
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_164
timestamp 1676037725
transform 1 0 16192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1676037725
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1676037725
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_261
timestamp 1676037725
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_268
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_280
timestamp 1676037725
transform 1 0 26864 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_296
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1676037725
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1676037725
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1676037725
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1676037725
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_375
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_381
timestamp 1676037725
transform 1 0 36156 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_397
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_409
timestamp 1676037725
transform 1 0 38732 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_417
timestamp 1676037725
transform 1 0 39468 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_441
timestamp 1676037725
transform 1 0 41676 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_458
timestamp 1676037725
transform 1 0 43240 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_139
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_151
timestamp 1676037725
transform 1 0 14996 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_191
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_202
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1676037725
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1676037725
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp 1676037725
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 1676037725
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_308
timestamp 1676037725
transform 1 0 29440 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_323
timestamp 1676037725
transform 1 0 30820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_355
timestamp 1676037725
transform 1 0 33764 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_368
timestamp 1676037725
transform 1 0 34960 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_380
timestamp 1676037725
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_402
timestamp 1676037725
transform 1 0 38088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_414
timestamp 1676037725
transform 1 0 39192 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_421
timestamp 1676037725
transform 1 0 39836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_433
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1676037725
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_460
timestamp 1676037725
transform 1 0 43424 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_156
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_168
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1676037725
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_212
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_232
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_242
timestamp 1676037725
transform 1 0 23368 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_263
timestamp 1676037725
transform 1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_270
timestamp 1676037725
transform 1 0 25944 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_282
timestamp 1676037725
transform 1 0 27048 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_299
timestamp 1676037725
transform 1 0 28612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_317
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_324
timestamp 1676037725
transform 1 0 30912 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_342
timestamp 1676037725
transform 1 0 32568 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_399
timestamp 1676037725
transform 1 0 37812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_407
timestamp 1676037725
transform 1 0 38548 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_430
timestamp 1676037725
transform 1 0 40664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_442
timestamp 1676037725
transform 1 0 41768 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_459
timestamp 1676037725
transform 1 0 43332 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 1676037725
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_177
timestamp 1676037725
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1676037725
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_255
timestamp 1676037725
transform 1 0 24564 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1676037725
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_291
timestamp 1676037725
transform 1 0 27876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_303
timestamp 1676037725
transform 1 0 28980 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_319
timestamp 1676037725
transform 1 0 30452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1676037725
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_378
timestamp 1676037725
transform 1 0 35880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_411
timestamp 1676037725
transform 1 0 38916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_420
timestamp 1676037725
transform 1 0 39744 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1676037725
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1676037725
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_453
timestamp 1676037725
transform 1 0 42780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_460
timestamp 1676037725
transform 1 0 43424 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1676037725
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_205
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_213
timestamp 1676037725
transform 1 0 20700 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_224
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_239
timestamp 1676037725
transform 1 0 23092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1676037725
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_269
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_281
timestamp 1676037725
transform 1 0 26956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_285
timestamp 1676037725
transform 1 0 27324 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_295
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_316
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_324
timestamp 1676037725
transform 1 0 30912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_344
timestamp 1676037725
transform 1 0 32752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_352
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_374
timestamp 1676037725
transform 1 0 35512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_394
timestamp 1676037725
transform 1 0 37352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_406
timestamp 1676037725
transform 1 0 38456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1676037725
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_430
timestamp 1676037725
transform 1 0 40664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_442
timestamp 1676037725
transform 1 0 41768 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_459
timestamp 1676037725
transform 1 0 43332 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_136
timestamp 1676037725
transform 1 0 13616 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_190
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_210
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_244
timestamp 1676037725
transform 1 0 23552 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_252
timestamp 1676037725
transform 1 0 24288 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_300
timestamp 1676037725
transform 1 0 28704 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_312
timestamp 1676037725
transform 1 0 29808 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_324
timestamp 1676037725
transform 1 0 30912 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1676037725
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_346
timestamp 1676037725
transform 1 0 32936 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_354
timestamp 1676037725
transform 1 0 33672 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_362
timestamp 1676037725
transform 1 0 34408 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_378
timestamp 1676037725
transform 1 0 35880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1676037725
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_402
timestamp 1676037725
transform 1 0 38088 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_416
timestamp 1676037725
transform 1 0 39376 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_428
timestamp 1676037725
transform 1 0 40480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_453
timestamp 1676037725
transform 1 0 42780 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_460
timestamp 1676037725
transform 1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1676037725
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1676037725
transform 1 0 14720 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_157
timestamp 1676037725
transform 1 0 15548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_263
timestamp 1676037725
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_275
timestamp 1676037725
transform 1 0 26404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_297
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1676037725
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_326
timestamp 1676037725
transform 1 0 31096 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_344
timestamp 1676037725
transform 1 0 32752 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_355
timestamp 1676037725
transform 1 0 33764 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_371
timestamp 1676037725
transform 1 0 35236 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_383
timestamp 1676037725
transform 1 0 36340 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_395
timestamp 1676037725
transform 1 0 37444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_407
timestamp 1676037725
transform 1 0 38548 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1676037725
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_429
timestamp 1676037725
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_441
timestamp 1676037725
transform 1 0 41676 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_458
timestamp 1676037725
transform 1 0 43240 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_140
timestamp 1676037725
transform 1 0 13984 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_152
timestamp 1676037725
transform 1 0 15088 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1676037725
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1676037725
transform 1 0 17204 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_183
timestamp 1676037725
transform 1 0 17940 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_201
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_213
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1676037725
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_250
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1676037725
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_301
timestamp 1676037725
transform 1 0 28796 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_309
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_328
timestamp 1676037725
transform 1 0 31280 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_360
timestamp 1676037725
transform 1 0 34224 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_368
timestamp 1676037725
transform 1 0 34960 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1676037725
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1676037725
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_403
timestamp 1676037725
transform 1 0 38180 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_419
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_431
timestamp 1676037725
transform 1 0 40756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_103
timestamp 1676037725
transform 1 0 10580 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_120
timestamp 1676037725
transform 1 0 12144 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1676037725
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_178
timestamp 1676037725
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_211
timestamp 1676037725
transform 1 0 20516 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1676037725
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_224
timestamp 1676037725
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_228
timestamp 1676037725
transform 1 0 22080 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_236
timestamp 1676037725
transform 1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1676037725
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_273
timestamp 1676037725
transform 1 0 26220 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_281
timestamp 1676037725
transform 1 0 26956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_332
timestamp 1676037725
transform 1 0 31648 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_344
timestamp 1676037725
transform 1 0 32752 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_371
timestamp 1676037725
transform 1 0 35236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_380
timestamp 1676037725
transform 1 0 36064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_392
timestamp 1676037725
transform 1 0 37168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_404
timestamp 1676037725
transform 1 0 38272 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1676037725
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_430
timestamp 1676037725
transform 1 0 40664 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_442
timestamp 1676037725
transform 1 0 41768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_446
timestamp 1676037725
transform 1 0 42136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_456
timestamp 1676037725
transform 1 0 43056 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_87
timestamp 1676037725
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1676037725
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_155
timestamp 1676037725
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_209
timestamp 1676037725
transform 1 0 20332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_233
timestamp 1676037725
transform 1 0 22540 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_241
timestamp 1676037725
transform 1 0 23276 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_246
timestamp 1676037725
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_257
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_267
timestamp 1676037725
transform 1 0 25668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_288
timestamp 1676037725
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_297
timestamp 1676037725
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_306
timestamp 1676037725
transform 1 0 29256 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1676037725
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_325
timestamp 1676037725
transform 1 0 31004 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1676037725
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_350
timestamp 1676037725
transform 1 0 33304 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_371
timestamp 1676037725
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_383
timestamp 1676037725
transform 1 0 36340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1676037725
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_453
timestamp 1676037725
transform 1 0 42780 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_460
timestamp 1676037725
transform 1 0 43424 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1676037725
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_104
timestamp 1676037725
transform 1 0 10672 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_128
timestamp 1676037725
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_154
timestamp 1676037725
transform 1 0 15272 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_172
timestamp 1676037725
transform 1 0 16928 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1676037725
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_205
timestamp 1676037725
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_217
timestamp 1676037725
transform 1 0 21068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_226
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_230
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1676037725
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_270
timestamp 1676037725
transform 1 0 25944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_278
timestamp 1676037725
transform 1 0 26680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_295
timestamp 1676037725
transform 1 0 28244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1676037725
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_320
timestamp 1676037725
transform 1 0 30544 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1676037725
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_341
timestamp 1676037725
transform 1 0 32476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_395
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1676037725
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_432
timestamp 1676037725
transform 1 0 40848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_460
timestamp 1676037725
transform 1 0 43424 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1676037725
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_90
timestamp 1676037725
transform 1 0 9384 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_98
timestamp 1676037725
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1676037725
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_121
timestamp 1676037725
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1676037725
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1676037725
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_182
timestamp 1676037725
transform 1 0 17848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1676037725
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_198
timestamp 1676037725
transform 1 0 19320 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_241
timestamp 1676037725
transform 1 0 23276 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_251
timestamp 1676037725
transform 1 0 24196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1676037725
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1676037725
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_300
timestamp 1676037725
transform 1 0 28704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_312
timestamp 1676037725
transform 1 0 29808 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1676037725
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_346
timestamp 1676037725
transform 1 0 32936 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_358
timestamp 1676037725
transform 1 0 34040 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_370
timestamp 1676037725
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_415
timestamp 1676037725
transform 1 0 39284 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_423
timestamp 1676037725
transform 1 0 40020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1676037725
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_460
timestamp 1676037725
transform 1 0 43424 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_123
timestamp 1676037725
transform 1 0 12420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_154
timestamp 1676037725
transform 1 0 15272 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_166
timestamp 1676037725
transform 1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1676037725
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_228
timestamp 1676037725
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1676037725
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 1676037725
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_279
timestamp 1676037725
transform 1 0 26772 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_288
timestamp 1676037725
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1676037725
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_315
timestamp 1676037725
transform 1 0 30084 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_325
timestamp 1676037725
transform 1 0 31004 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_335
timestamp 1676037725
transform 1 0 31924 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_346
timestamp 1676037725
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1676037725
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_381
timestamp 1676037725
transform 1 0 36156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_391
timestamp 1676037725
transform 1 0 37076 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_398
timestamp 1676037725
transform 1 0 37720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_410
timestamp 1676037725
transform 1 0 38824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1676037725
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_425
timestamp 1676037725
transform 1 0 40204 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_431
timestamp 1676037725
transform 1 0 40756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_443
timestamp 1676037725
transform 1 0 41860 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_451
timestamp 1676037725
transform 1 0 42596 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_460
timestamp 1676037725
transform 1 0 43424 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_126
timestamp 1676037725
transform 1 0 12696 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_138
timestamp 1676037725
transform 1 0 13800 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1676037725
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_201
timestamp 1676037725
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_210
timestamp 1676037725
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1676037725
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_297
timestamp 1676037725
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_309
timestamp 1676037725
transform 1 0 29532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_321
timestamp 1676037725
transform 1 0 30636 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1676037725
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_343
timestamp 1676037725
transform 1 0 32660 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_352
timestamp 1676037725
transform 1 0 33488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_360
timestamp 1676037725
transform 1 0 34224 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_372
timestamp 1676037725
transform 1 0 35328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_380
timestamp 1676037725
transform 1 0 36064 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1676037725
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_416
timestamp 1676037725
transform 1 0 39376 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_420
timestamp 1676037725
transform 1 0 39744 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1676037725
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1676037725
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_453
timestamp 1676037725
transform 1 0 42780 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_460
timestamp 1676037725
transform 1 0 43424 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_94
timestamp 1676037725
transform 1 0 9752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_102
timestamp 1676037725
transform 1 0 10488 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1676037725
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_127
timestamp 1676037725
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_160
timestamp 1676037725
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_168
timestamp 1676037725
transform 1 0 16560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1676037725
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_215
timestamp 1676037725
transform 1 0 20884 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_227
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_235
timestamp 1676037725
transform 1 0 22724 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_275
timestamp 1676037725
transform 1 0 26404 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_290
timestamp 1676037725
transform 1 0 27784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_315
timestamp 1676037725
transform 1 0 30084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_323
timestamp 1676037725
transform 1 0 30820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_331
timestamp 1676037725
transform 1 0 31556 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_339
timestamp 1676037725
transform 1 0 32292 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_350
timestamp 1676037725
transform 1 0 33304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_354
timestamp 1676037725
transform 1 0 33672 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1676037725
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_373
timestamp 1676037725
transform 1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_381
timestamp 1676037725
transform 1 0 36156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_391
timestamp 1676037725
transform 1 0 37076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_395
timestamp 1676037725
transform 1 0 37444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_404
timestamp 1676037725
transform 1 0 38272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1676037725
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_432
timestamp 1676037725
transform 1 0 40848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_460
timestamp 1676037725
transform 1 0 43424 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1676037725
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_82
timestamp 1676037725
transform 1 0 8648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_89
timestamp 1676037725
transform 1 0 9292 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_97
timestamp 1676037725
transform 1 0 10028 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_135
timestamp 1676037725
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_147
timestamp 1676037725
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_159
timestamp 1676037725
transform 1 0 15732 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1676037725
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1676037725
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_204
timestamp 1676037725
transform 1 0 19872 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_212
timestamp 1676037725
transform 1 0 20608 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1676037725
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1676037725
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_246
timestamp 1676037725
transform 1 0 23736 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_254
timestamp 1676037725
transform 1 0 24472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1676037725
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_302
timestamp 1676037725
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_309
timestamp 1676037725
transform 1 0 29532 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_315
timestamp 1676037725
transform 1 0 30084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1676037725
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_348
timestamp 1676037725
transform 1 0 33120 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_354
timestamp 1676037725
transform 1 0 33672 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_362
timestamp 1676037725
transform 1 0 34408 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_374
timestamp 1676037725
transform 1 0 35512 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1676037725
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_406
timestamp 1676037725
transform 1 0 38456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_418
timestamp 1676037725
transform 1 0 39560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_426
timestamp 1676037725
transform 1 0 40296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1676037725
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_460
timestamp 1676037725
transform 1 0 43424 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_61
timestamp 1676037725
transform 1 0 6716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_69
timestamp 1676037725
transform 1 0 7452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1676037725
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_93
timestamp 1676037725
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1676037725
transform 1 0 11224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_114
timestamp 1676037725
transform 1 0 11592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_131
timestamp 1676037725
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_171
timestamp 1676037725
transform 1 0 16836 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_182
timestamp 1676037725
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_228
timestamp 1676037725
transform 1 0 22080 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_236
timestamp 1676037725
transform 1 0 22816 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1676037725
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_273
timestamp 1676037725
transform 1 0 26220 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_281
timestamp 1676037725
transform 1 0 26956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_290
timestamp 1676037725
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1676037725
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_318
timestamp 1676037725
transform 1 0 30360 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_327
timestamp 1676037725
transform 1 0 31188 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_339
timestamp 1676037725
transform 1 0 32292 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_348
timestamp 1676037725
transform 1 0 33120 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1676037725
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_376
timestamp 1676037725
transform 1 0 35696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_387
timestamp 1676037725
transform 1 0 36708 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_402
timestamp 1676037725
transform 1 0 38088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_430
timestamp 1676037725
transform 1 0 40664 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_442
timestamp 1676037725
transform 1 0 41768 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_460
timestamp 1676037725
transform 1 0 43424 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_68
timestamp 1676037725
transform 1 0 7360 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_79
timestamp 1676037725
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_91
timestamp 1676037725
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1676037725
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_117
timestamp 1676037725
transform 1 0 11868 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_154
timestamp 1676037725
transform 1 0 15272 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_175
timestamp 1676037725
transform 1 0 17204 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_185
timestamp 1676037725
transform 1 0 18124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_197
timestamp 1676037725
transform 1 0 19228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_233
timestamp 1676037725
transform 1 0 22540 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1676037725
transform 1 0 23644 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_258
timestamp 1676037725
transform 1 0 24840 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_270
timestamp 1676037725
transform 1 0 25944 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1676037725
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_303
timestamp 1676037725
transform 1 0 28980 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_315
timestamp 1676037725
transform 1 0 30084 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_328
timestamp 1676037725
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_346
timestamp 1676037725
transform 1 0 32936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_354
timestamp 1676037725
transform 1 0 33672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_358
timestamp 1676037725
transform 1 0 34040 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_372
timestamp 1676037725
transform 1 0 35328 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_378
timestamp 1676037725
transform 1 0 35880 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1676037725
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_403
timestamp 1676037725
transform 1 0 38180 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_411
timestamp 1676037725
transform 1 0 38916 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_418
timestamp 1676037725
transform 1 0 39560 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_430
timestamp 1676037725
transform 1 0 40664 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_442
timestamp 1676037725
transform 1 0 41768 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_460
timestamp 1676037725
transform 1 0 43424 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_47
timestamp 1676037725
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_64
timestamp 1676037725
transform 1 0 6992 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_72
timestamp 1676037725
transform 1 0 7728 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1676037725
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_103
timestamp 1676037725
transform 1 0 10580 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_115
timestamp 1676037725
transform 1 0 11684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_150
timestamp 1676037725
transform 1 0 14904 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_173
timestamp 1676037725
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1676037725
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_217
timestamp 1676037725
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_229
timestamp 1676037725
transform 1 0 22172 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_240
timestamp 1676037725
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_257
timestamp 1676037725
transform 1 0 24748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_274
timestamp 1676037725
transform 1 0 26312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_287
timestamp 1676037725
transform 1 0 27508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_291
timestamp 1676037725
transform 1 0 27876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1676037725
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_315
timestamp 1676037725
transform 1 0 30084 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_320
timestamp 1676037725
transform 1 0 30544 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_341
timestamp 1676037725
transform 1 0 32476 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_350
timestamp 1676037725
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1676037725
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_376
timestamp 1676037725
transform 1 0 35696 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_388
timestamp 1676037725
transform 1 0 36800 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_399
timestamp 1676037725
transform 1 0 37812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_407
timestamp 1676037725
transform 1 0 38548 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1676037725
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_430
timestamp 1676037725
transform 1 0 40664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_442
timestamp 1676037725
transform 1 0 41768 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_459
timestamp 1676037725
transform 1 0 43332 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_88
timestamp 1676037725
transform 1 0 9200 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_190
timestamp 1676037725
transform 1 0 18584 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_196
timestamp 1676037725
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_202
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1676037725
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_268
timestamp 1676037725
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_287
timestamp 1676037725
transform 1 0 27508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_291
timestamp 1676037725
transform 1 0 27876 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_295
timestamp 1676037725
transform 1 0 28244 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_301
timestamp 1676037725
transform 1 0 28796 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_309
timestamp 1676037725
transform 1 0 29532 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1676037725
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_326
timestamp 1676037725
transform 1 0 31096 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_352
timestamp 1676037725
transform 1 0 33488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_360
timestamp 1676037725
transform 1 0 34224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_369
timestamp 1676037725
transform 1 0 35052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_404
timestamp 1676037725
transform 1 0 38272 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_410
timestamp 1676037725
transform 1 0 38824 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_419
timestamp 1676037725
transform 1 0 39652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_428
timestamp 1676037725
transform 1 0 40480 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_436
timestamp 1676037725
transform 1 0 41216 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_59
timestamp 1676037725
transform 1 0 6532 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_67
timestamp 1676037725
transform 1 0 7268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_115
timestamp 1676037725
transform 1 0 11684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_123
timestamp 1676037725
transform 1 0 12420 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1676037725
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_161
timestamp 1676037725
transform 1 0 15916 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_173
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1676037725
transform 1 0 18032 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_207
timestamp 1676037725
transform 1 0 20148 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_214
timestamp 1676037725
transform 1 0 20792 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_226
timestamp 1676037725
transform 1 0 21896 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_234
timestamp 1676037725
transform 1 0 22632 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_273
timestamp 1676037725
transform 1 0 26220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_282
timestamp 1676037725
transform 1 0 27048 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_294
timestamp 1676037725
transform 1 0 28152 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1676037725
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_324
timestamp 1676037725
transform 1 0 30912 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_335
timestamp 1676037725
transform 1 0 31924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_342
timestamp 1676037725
transform 1 0 32568 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_354
timestamp 1676037725
transform 1 0 33672 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1676037725
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_376
timestamp 1676037725
transform 1 0 35696 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_382
timestamp 1676037725
transform 1 0 36248 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_400
timestamp 1676037725
transform 1 0 37904 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_412
timestamp 1676037725
transform 1 0 39008 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_427
timestamp 1676037725
transform 1 0 40388 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_453
timestamp 1676037725
transform 1 0 42780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_460
timestamp 1676037725
transform 1 0 43424 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1676037725
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_89
timestamp 1676037725
transform 1 0 9292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_101
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_133
timestamp 1676037725
transform 1 0 13340 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_139
timestamp 1676037725
transform 1 0 13892 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_147
timestamp 1676037725
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_159
timestamp 1676037725
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1676037725
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_184
timestamp 1676037725
transform 1 0 18032 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1676037725
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_207
timestamp 1676037725
transform 1 0 20148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_215
timestamp 1676037725
transform 1 0 20884 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1676037725
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1676037725
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_268
timestamp 1676037725
transform 1 0 25760 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_272
timestamp 1676037725
transform 1 0 26128 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1676037725
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_289
timestamp 1676037725
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1676037725
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_312
timestamp 1676037725
transform 1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1676037725
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1676037725
transform 1 0 33672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_369
timestamp 1676037725
transform 1 0 35052 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_380
timestamp 1676037725
transform 1 0 36064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1676037725
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_419
timestamp 1676037725
transform 1 0 39652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_423
timestamp 1676037725
transform 1 0 40020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_436
timestamp 1676037725
transform 1 0 41216 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_460
timestamp 1676037725
transform 1 0 43424 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_37
timestamp 1676037725
transform 1 0 4508 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_49
timestamp 1676037725
transform 1 0 5612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_61
timestamp 1676037725
transform 1 0 6716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_70
timestamp 1676037725
transform 1 0 7544 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1676037725
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_110
timestamp 1676037725
transform 1 0 11224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_130
timestamp 1676037725
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1676037725
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_162
timestamp 1676037725
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_174
timestamp 1676037725
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1676037725
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_203
timestamp 1676037725
transform 1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1676037725
transform 1 0 20424 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_239
timestamp 1676037725
transform 1 0 23092 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_262
timestamp 1676037725
transform 1 0 25208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_275
timestamp 1676037725
transform 1 0 26404 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_283
timestamp 1676037725
transform 1 0 27140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_293
timestamp 1676037725
transform 1 0 28060 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1676037725
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_317
timestamp 1676037725
transform 1 0 30268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_336
timestamp 1676037725
transform 1 0 32016 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_344
timestamp 1676037725
transform 1 0 32752 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_353
timestamp 1676037725
transform 1 0 33580 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1676037725
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_376
timestamp 1676037725
transform 1 0 35696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_387
timestamp 1676037725
transform 1 0 36708 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_400
timestamp 1676037725
transform 1 0 37904 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_408
timestamp 1676037725
transform 1 0 38640 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1676037725
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_429
timestamp 1676037725
transform 1 0 40572 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_441
timestamp 1676037725
transform 1 0 41676 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_460
timestamp 1676037725
transform 1 0 43424 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_61
timestamp 1676037725
transform 1 0 6716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_68
timestamp 1676037725
transform 1 0 7360 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_83
timestamp 1676037725
transform 1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_94
timestamp 1676037725
transform 1 0 9752 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_106
timestamp 1676037725
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_121
timestamp 1676037725
transform 1 0 12236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_130
timestamp 1676037725
transform 1 0 13064 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_136
timestamp 1676037725
transform 1 0 13616 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_142
timestamp 1676037725
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_154
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_198
timestamp 1676037725
transform 1 0 19320 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1676037725
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_244
timestamp 1676037725
transform 1 0 23552 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_251
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_259
timestamp 1676037725
transform 1 0 24932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_268
timestamp 1676037725
transform 1 0 25760 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_330
timestamp 1676037725
transform 1 0 31464 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_345
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_365
timestamp 1676037725
transform 1 0 34684 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_377
timestamp 1676037725
transform 1 0 35788 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1676037725
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_399
timestamp 1676037725
transform 1 0 37812 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_407
timestamp 1676037725
transform 1 0 38548 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_419
timestamp 1676037725
transform 1 0 39652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_431
timestamp 1676037725
transform 1 0 40756 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_436
timestamp 1676037725
transform 1 0 41216 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_453
timestamp 1676037725
transform 1 0 42780 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_460
timestamp 1676037725
transform 1 0 43424 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_37
timestamp 1676037725
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_47
timestamp 1676037725
transform 1 0 5428 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_61
timestamp 1676037725
transform 1 0 6716 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_68
timestamp 1676037725
transform 1 0 7360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1676037725
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_93
timestamp 1676037725
transform 1 0 9660 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_99
timestamp 1676037725
transform 1 0 10212 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_107
timestamp 1676037725
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_119
timestamp 1676037725
transform 1 0 12052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_125
timestamp 1676037725
transform 1 0 12604 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1676037725
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_159
timestamp 1676037725
transform 1 0 15732 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_182
timestamp 1676037725
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_218
timestamp 1676037725
transform 1 0 21160 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_229
timestamp 1676037725
transform 1 0 22172 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_275
timestamp 1676037725
transform 1 0 26404 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_282
timestamp 1676037725
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_294
timestamp 1676037725
transform 1 0 28152 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_314
timestamp 1676037725
transform 1 0 29992 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_326
timestamp 1676037725
transform 1 0 31096 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 1676037725
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_354
timestamp 1676037725
transform 1 0 33672 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1676037725
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_379
timestamp 1676037725
transform 1 0 35972 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_387
timestamp 1676037725
transform 1 0 36708 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_396
timestamp 1676037725
transform 1 0 37536 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_407
timestamp 1676037725
transform 1 0 38548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_425
timestamp 1676037725
transform 1 0 40204 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_434
timestamp 1676037725
transform 1 0 41032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_438
timestamp 1676037725
transform 1 0 41400 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_456
timestamp 1676037725
transform 1 0 43056 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_47
timestamp 1676037725
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_73
timestamp 1676037725
transform 1 0 7820 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_84
timestamp 1676037725
transform 1 0 8832 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_121
timestamp 1676037725
transform 1 0 12236 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_134
timestamp 1676037725
transform 1 0 13432 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_145
timestamp 1676037725
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1676037725
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_204
timestamp 1676037725
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_214
timestamp 1676037725
transform 1 0 20792 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_233
timestamp 1676037725
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1676037725
transform 1 0 25760 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1676037725
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_292
timestamp 1676037725
transform 1 0 27968 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_301
timestamp 1676037725
transform 1 0 28796 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_310
timestamp 1676037725
transform 1 0 29624 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_322
timestamp 1676037725
transform 1 0 30728 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1676037725
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_355
timestamp 1676037725
transform 1 0 33764 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_363
timestamp 1676037725
transform 1 0 34500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_381
timestamp 1676037725
transform 1 0 36156 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1676037725
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_397
timestamp 1676037725
transform 1 0 37628 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_413
timestamp 1676037725
transform 1 0 39100 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_420
timestamp 1676037725
transform 1 0 39744 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_432
timestamp 1676037725
transform 1 0 40848 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_444
timestamp 1676037725
transform 1 0 41952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_460
timestamp 1676037725
transform 1 0 43424 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_48
timestamp 1676037725
transform 1 0 5520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_63
timestamp 1676037725
transform 1 0 6900 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1676037725
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_94
timestamp 1676037725
transform 1 0 9752 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_102
timestamp 1676037725
transform 1 0 10488 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_108
timestamp 1676037725
transform 1 0 11040 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_116
timestamp 1676037725
transform 1 0 11776 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_124
timestamp 1676037725
transform 1 0 12512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1676037725
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1676037725
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_206
timestamp 1676037725
transform 1 0 20056 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_214
timestamp 1676037725
transform 1 0 20792 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1676037725
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1676037725
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_274
timestamp 1676037725
transform 1 0 26312 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_280
timestamp 1676037725
transform 1 0 26864 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_286
timestamp 1676037725
transform 1 0 27416 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_294
timestamp 1676037725
transform 1 0 28152 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_332
timestamp 1676037725
transform 1 0 31648 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1676037725
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_376
timestamp 1676037725
transform 1 0 35696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_405
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_415
timestamp 1676037725
transform 1 0 39284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_439
timestamp 1676037725
transform 1 0 41492 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_451
timestamp 1676037725
transform 1 0 42596 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_460
timestamp 1676037725
transform 1 0 43424 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1676037725
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_66
timestamp 1676037725
transform 1 0 7176 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_78
timestamp 1676037725
transform 1 0 8280 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_82
timestamp 1676037725
transform 1 0 8648 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_90
timestamp 1676037725
transform 1 0 9384 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_98
timestamp 1676037725
transform 1 0 10120 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1676037725
transform 1 0 10948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_117
timestamp 1676037725
transform 1 0 11868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_129
timestamp 1676037725
transform 1 0 12972 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_139
timestamp 1676037725
transform 1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_146
timestamp 1676037725
transform 1 0 14536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1676037725
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1676037725
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_187
timestamp 1676037725
transform 1 0 18308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_195
timestamp 1676037725
transform 1 0 19044 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_214
timestamp 1676037725
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_241
timestamp 1676037725
transform 1 0 23276 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_260
timestamp 1676037725
transform 1 0 25024 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1676037725
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_303
timestamp 1676037725
transform 1 0 28980 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_322
timestamp 1676037725
transform 1 0 30728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_345
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_368
timestamp 1676037725
transform 1 0 34960 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1676037725
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_420
timestamp 1676037725
transform 1 0 39744 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_426
timestamp 1676037725
transform 1 0 40296 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_435
timestamp 1676037725
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_460
timestamp 1676037725
transform 1 0 43424 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_49
timestamp 1676037725
transform 1 0 5612 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_59
timestamp 1676037725
transform 1 0 6532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_66
timestamp 1676037725
transform 1 0 7176 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_74
timestamp 1676037725
transform 1 0 7912 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_79
timestamp 1676037725
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1676037725
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_102
timestamp 1676037725
transform 1 0 10488 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1676037725
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_129
timestamp 1676037725
transform 1 0 12972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1676037725
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1676037725
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_174
timestamp 1676037725
transform 1 0 17112 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_205
timestamp 1676037725
transform 1 0 19964 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_217
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_227
timestamp 1676037725
transform 1 0 21988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1676037725
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1676037725
transform 1 0 26036 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_275
timestamp 1676037725
transform 1 0 26404 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1676037725
transform 1 0 26956 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_288
timestamp 1676037725
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_295
timestamp 1676037725
transform 1 0 28244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_316
timestamp 1676037725
transform 1 0 30176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_329
timestamp 1676037725
transform 1 0 31372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_338
timestamp 1676037725
transform 1 0 32200 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_350
timestamp 1676037725
transform 1 0 33304 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_354
timestamp 1676037725
transform 1 0 33672 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1676037725
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_372
timestamp 1676037725
transform 1 0 35328 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_381
timestamp 1676037725
transform 1 0 36156 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_393
timestamp 1676037725
transform 1 0 37260 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_405
timestamp 1676037725
transform 1 0 38364 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_417
timestamp 1676037725
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_441
timestamp 1676037725
transform 1 0 41676 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_460
timestamp 1676037725
transform 1 0 43424 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1676037725
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_71
timestamp 1676037725
transform 1 0 7636 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_77
timestamp 1676037725
transform 1 0 8188 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_83
timestamp 1676037725
transform 1 0 8740 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_100
timestamp 1676037725
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_118
timestamp 1676037725
transform 1 0 11960 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_131
timestamp 1676037725
transform 1 0 13156 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_140
timestamp 1676037725
transform 1 0 13984 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_147
timestamp 1676037725
transform 1 0 14628 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_159
timestamp 1676037725
transform 1 0 15732 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_201
timestamp 1676037725
transform 1 0 19596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_213
timestamp 1676037725
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1676037725
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_233
timestamp 1676037725
transform 1 0 22540 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_251
timestamp 1676037725
transform 1 0 24196 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_285
timestamp 1676037725
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_291
timestamp 1676037725
transform 1 0 27876 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_345
timestamp 1676037725
transform 1 0 32844 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_355
timestamp 1676037725
transform 1 0 33764 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_372
timestamp 1676037725
transform 1 0 35328 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_378
timestamp 1676037725
transform 1 0 35880 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_387
timestamp 1676037725
transform 1 0 36708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_458
timestamp 1676037725
transform 1 0 43240 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_45
timestamp 1676037725
transform 1 0 5244 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_51
timestamp 1676037725
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_63
timestamp 1676037725
transform 1 0 6900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_76
timestamp 1676037725
transform 1 0 8096 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_92
timestamp 1676037725
transform 1 0 9568 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_104
timestamp 1676037725
transform 1 0 10672 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_110
timestamp 1676037725
transform 1 0 11224 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_118
timestamp 1676037725
transform 1 0 11960 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_128
timestamp 1676037725
transform 1 0 12880 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_149
timestamp 1676037725
transform 1 0 14812 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 1676037725
transform 1 0 15364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_162
timestamp 1676037725
transform 1 0 16008 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_170
timestamp 1676037725
transform 1 0 16744 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_184
timestamp 1676037725
transform 1 0 18032 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_208
timestamp 1676037725
transform 1 0 20240 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_220
timestamp 1676037725
transform 1 0 21344 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_228
timestamp 1676037725
transform 1 0 22080 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1676037725
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1676037725
transform 1 0 25576 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_275
timestamp 1676037725
transform 1 0 26404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_285
timestamp 1676037725
transform 1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_292
timestamp 1676037725
transform 1 0 27968 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_298
timestamp 1676037725
transform 1 0 28520 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1676037725
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1676037725
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_329
timestamp 1676037725
transform 1 0 31372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_355
timestamp 1676037725
transform 1 0 33764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1676037725
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_385
timestamp 1676037725
transform 1 0 36524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_398
timestamp 1676037725
transform 1 0 37720 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_409
timestamp 1676037725
transform 1 0 38732 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 1676037725
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_439
timestamp 1676037725
transform 1 0 41492 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_443
timestamp 1676037725
transform 1 0 41860 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_450
timestamp 1676037725
transform 1 0 42504 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_460
timestamp 1676037725
transform 1 0 43424 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_49
timestamp 1676037725
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_72
timestamp 1676037725
transform 1 0 7728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_76
timestamp 1676037725
transform 1 0 8096 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_80
timestamp 1676037725
transform 1 0 8464 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_102
timestamp 1676037725
transform 1 0 10488 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_120
timestamp 1676037725
transform 1 0 12144 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_131
timestamp 1676037725
transform 1 0 13156 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_150
timestamp 1676037725
transform 1 0 14904 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_154
timestamp 1676037725
transform 1 0 15272 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_158
timestamp 1676037725
transform 1 0 15640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1676037725
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_175
timestamp 1676037725
transform 1 0 17204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_179
timestamp 1676037725
transform 1 0 17572 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_187
timestamp 1676037725
transform 1 0 18308 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_194
timestamp 1676037725
transform 1 0 18952 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_206
timestamp 1676037725
transform 1 0 20056 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_213
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 1676037725
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_235
timestamp 1676037725
transform 1 0 22724 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_246
timestamp 1676037725
transform 1 0 23736 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_254
timestamp 1676037725
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_265
timestamp 1676037725
transform 1 0 25484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_294
timestamp 1676037725
transform 1 0 28152 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_302
timestamp 1676037725
transform 1 0 28888 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_309
timestamp 1676037725
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_322
timestamp 1676037725
transform 1 0 30728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1676037725
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_345
timestamp 1676037725
transform 1 0 32844 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_355
timestamp 1676037725
transform 1 0 33764 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_362
timestamp 1676037725
transform 1 0 34408 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_374
timestamp 1676037725
transform 1 0 35512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_386
timestamp 1676037725
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_399
timestamp 1676037725
transform 1 0 37812 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_406
timestamp 1676037725
transform 1 0 38456 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_460
timestamp 1676037725
transform 1 0 43424 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_49
timestamp 1676037725
transform 1 0 5612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_56
timestamp 1676037725
transform 1 0 6256 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_67
timestamp 1676037725
transform 1 0 7268 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_75
timestamp 1676037725
transform 1 0 8004 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_89
timestamp 1676037725
transform 1 0 9292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_103
timestamp 1676037725
transform 1 0 10580 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_117
timestamp 1676037725
transform 1 0 11868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_129
timestamp 1676037725
transform 1 0 12972 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_149
timestamp 1676037725
transform 1 0 14812 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_157
timestamp 1676037725
transform 1 0 15548 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1676037725
transform 1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_188
timestamp 1676037725
transform 1 0 18400 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_206
timestamp 1676037725
transform 1 0 20056 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_220
timestamp 1676037725
transform 1 0 21344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1676037725
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_238
timestamp 1676037725
transform 1 0 23000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_242
timestamp 1676037725
transform 1 0 23368 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1676037725
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_263
timestamp 1676037725
transform 1 0 25300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_275
timestamp 1676037725
transform 1 0 26404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_294
timestamp 1676037725
transform 1 0 28152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1676037725
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_320
timestamp 1676037725
transform 1 0 30544 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_332
timestamp 1676037725
transform 1 0 31648 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_342
timestamp 1676037725
transform 1 0 32568 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_350
timestamp 1676037725
transform 1 0 33304 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_361
timestamp 1676037725
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_383
timestamp 1676037725
transform 1 0 36340 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1676037725
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1676037725
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_410
timestamp 1676037725
transform 1 0 38824 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1676037725
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_430
timestamp 1676037725
transform 1 0 40664 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_442
timestamp 1676037725
transform 1 0 41768 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_460
timestamp 1676037725
transform 1 0 43424 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_66
timestamp 1676037725
transform 1 0 7176 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_70
timestamp 1676037725
transform 1 0 7544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_76
timestamp 1676037725
transform 1 0 8096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_91
timestamp 1676037725
transform 1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_101
timestamp 1676037725
transform 1 0 10396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_127
timestamp 1676037725
transform 1 0 12788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_131
timestamp 1676037725
transform 1 0 13156 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_138
timestamp 1676037725
transform 1 0 13800 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_146
timestamp 1676037725
transform 1 0 14536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_152
timestamp 1676037725
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_180
timestamp 1676037725
transform 1 0 17664 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_192
timestamp 1676037725
transform 1 0 18768 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_204
timestamp 1676037725
transform 1 0 19872 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 1676037725
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1676037725
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1676037725
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_252
timestamp 1676037725
transform 1 0 24288 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1676037725
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1676037725
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1676037725
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_348
timestamp 1676037725
transform 1 0 33120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_357
timestamp 1676037725
transform 1 0 33948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_375
timestamp 1676037725
transform 1 0 35604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1676037725
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_460
timestamp 1676037725
transform 1 0 43424 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_50
timestamp 1676037725
transform 1 0 5704 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_56
timestamp 1676037725
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_63
timestamp 1676037725
transform 1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_72
timestamp 1676037725
transform 1 0 7728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_76
timestamp 1676037725
transform 1 0 8096 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_101
timestamp 1676037725
transform 1 0 10396 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1676037725
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_126
timestamp 1676037725
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1676037725
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_150
timestamp 1676037725
transform 1 0 14904 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_162
timestamp 1676037725
transform 1 0 16008 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_175
timestamp 1676037725
transform 1 0 17204 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_187
timestamp 1676037725
transform 1 0 18308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_216
timestamp 1676037725
transform 1 0 20976 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_228
timestamp 1676037725
transform 1 0 22080 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_235
timestamp 1676037725
transform 1 0 22724 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1676037725
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_262
timestamp 1676037725
transform 1 0 25208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_271
timestamp 1676037725
transform 1 0 26036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_282
timestamp 1676037725
transform 1 0 27048 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_291
timestamp 1676037725
transform 1 0 27876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_299
timestamp 1676037725
transform 1 0 28612 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1676037725
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_320
timestamp 1676037725
transform 1 0 30544 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_351
timestamp 1676037725
transform 1 0 33396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 1676037725
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_380
timestamp 1676037725
transform 1 0 36064 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_394
timestamp 1676037725
transform 1 0 37352 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_406
timestamp 1676037725
transform 1 0 38456 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_410
timestamp 1676037725
transform 1 0 38824 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1676037725
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_432
timestamp 1676037725
transform 1 0 40848 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_440
timestamp 1676037725
transform 1 0 41584 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_458
timestamp 1676037725
transform 1 0 43240 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_70
timestamp 1676037725
transform 1 0 7544 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_80
timestamp 1676037725
transform 1 0 8464 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_100
timestamp 1676037725
transform 1 0 10304 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_110
timestamp 1676037725
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_122
timestamp 1676037725
transform 1 0 12328 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_131
timestamp 1676037725
transform 1 0 13156 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_147
timestamp 1676037725
transform 1 0 14628 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_176
timestamp 1676037725
transform 1 0 17296 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_187
timestamp 1676037725
transform 1 0 18308 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_199
timestamp 1676037725
transform 1 0 19412 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_208
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1676037725
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_236
timestamp 1676037725
transform 1 0 22816 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_245
timestamp 1676037725
transform 1 0 23644 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_261
timestamp 1676037725
transform 1 0 25116 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1676037725
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_286
timestamp 1676037725
transform 1 0 27416 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_298
timestamp 1676037725
transform 1 0 28520 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_303
timestamp 1676037725
transform 1 0 28980 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_312
timestamp 1676037725
transform 1 0 29808 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_319
timestamp 1676037725
transform 1 0 30452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_327
timestamp 1676037725
transform 1 0 31188 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1676037725
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_346
timestamp 1676037725
transform 1 0 32936 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_360
timestamp 1676037725
transform 1 0 34224 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_369
timestamp 1676037725
transform 1 0 35052 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_404
timestamp 1676037725
transform 1 0 38272 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_437
timestamp 1676037725
transform 1 0 41308 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_445
timestamp 1676037725
transform 1 0 42044 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_453
timestamp 1676037725
transform 1 0 42780 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_460
timestamp 1676037725
transform 1 0 43424 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_49
timestamp 1676037725
transform 1 0 5612 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_55
timestamp 1676037725
transform 1 0 6164 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_66
timestamp 1676037725
transform 1 0 7176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_79
timestamp 1676037725
transform 1 0 8372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_103
timestamp 1676037725
transform 1 0 10580 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_111
timestamp 1676037725
transform 1 0 11316 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_120
timestamp 1676037725
transform 1 0 12144 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_128
timestamp 1676037725
transform 1 0 12880 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1676037725
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_152
timestamp 1676037725
transform 1 0 15088 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_160
timestamp 1676037725
transform 1 0 15824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_170
timestamp 1676037725
transform 1 0 16744 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_183
timestamp 1676037725
transform 1 0 17940 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1676037725
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_204
timestamp 1676037725
transform 1 0 19872 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_214
timestamp 1676037725
transform 1 0 20792 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_224
timestamp 1676037725
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_236
timestamp 1676037725
transform 1 0 22816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_242
timestamp 1676037725
transform 1 0 23368 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1676037725
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_263
timestamp 1676037725
transform 1 0 25300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_275
timestamp 1676037725
transform 1 0 26404 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_279
timestamp 1676037725
transform 1 0 26772 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_287
timestamp 1676037725
transform 1 0 27508 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_291
timestamp 1676037725
transform 1 0 27876 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_299
timestamp 1676037725
transform 1 0 28612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_320
timestamp 1676037725
transform 1 0 30544 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_328
timestamp 1676037725
transform 1 0 31280 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_336
timestamp 1676037725
transform 1 0 32016 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_348
timestamp 1676037725
transform 1 0 33120 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_352
timestamp 1676037725
transform 1 0 33488 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1676037725
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_370
timestamp 1676037725
transform 1 0 35144 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_390
timestamp 1676037725
transform 1 0 36984 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_394
timestamp 1676037725
transform 1 0 37352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_403
timestamp 1676037725
transform 1 0 38180 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_418
timestamp 1676037725
transform 1 0 39560 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_431
timestamp 1676037725
transform 1 0 40756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_439
timestamp 1676037725
transform 1 0 41492 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_459
timestamp 1676037725
transform 1 0 43332 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_47
timestamp 1676037725
transform 1 0 5428 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1676037725
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_70
timestamp 1676037725
transform 1 0 7544 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_78
timestamp 1676037725
transform 1 0 8280 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_86
timestamp 1676037725
transform 1 0 9016 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1676037725
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_123
timestamp 1676037725
transform 1 0 12420 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_150
timestamp 1676037725
transform 1 0 14904 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_174
timestamp 1676037725
transform 1 0 17112 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_186
timestamp 1676037725
transform 1 0 18216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_195
timestamp 1676037725
transform 1 0 19044 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_207
timestamp 1676037725
transform 1 0 20148 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_213
timestamp 1676037725
transform 1 0 20700 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1676037725
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_231
timestamp 1676037725
transform 1 0 22356 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_244
timestamp 1676037725
transform 1 0 23552 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_252
timestamp 1676037725
transform 1 0 24288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_262
timestamp 1676037725
transform 1 0 25208 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_270
timestamp 1676037725
transform 1 0 25944 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1676037725
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_290
timestamp 1676037725
transform 1 0 27784 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_297
timestamp 1676037725
transform 1 0 28428 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_301
timestamp 1676037725
transform 1 0 28796 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_306
timestamp 1676037725
transform 1 0 29256 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_319
timestamp 1676037725
transform 1 0 30452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_327
timestamp 1676037725
transform 1 0 31188 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1676037725
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_355
timestamp 1676037725
transform 1 0 33764 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_362
timestamp 1676037725
transform 1 0 34408 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_381
timestamp 1676037725
transform 1 0 36156 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1676037725
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_404
timestamp 1676037725
transform 1 0 38272 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_415
timestamp 1676037725
transform 1 0 39284 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_427
timestamp 1676037725
transform 1 0 40388 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_439
timestamp 1676037725
transform 1 0 41492 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_460
timestamp 1676037725
transform 1 0 43424 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_66
timestamp 1676037725
transform 1 0 7176 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_78
timestamp 1676037725
transform 1 0 8280 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_92
timestamp 1676037725
transform 1 0 9568 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_100
timestamp 1676037725
transform 1 0 10304 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_106
timestamp 1676037725
transform 1 0 10856 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_120
timestamp 1676037725
transform 1 0 12144 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_132
timestamp 1676037725
transform 1 0 13248 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_161
timestamp 1676037725
transform 1 0 15916 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_167
timestamp 1676037725
transform 1 0 16468 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_175
timestamp 1676037725
transform 1 0 17204 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_182
timestamp 1676037725
transform 1 0 17848 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_205
timestamp 1676037725
transform 1 0 19964 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_210
timestamp 1676037725
transform 1 0 20424 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_219
timestamp 1676037725
transform 1 0 21252 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_231
timestamp 1676037725
transform 1 0 22356 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_240
timestamp 1676037725
transform 1 0 23184 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1676037725
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_283
timestamp 1676037725
transform 1 0 27140 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_313
timestamp 1676037725
transform 1 0 29900 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_322
timestamp 1676037725
transform 1 0 30728 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_330
timestamp 1676037725
transform 1 0 31464 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_339
timestamp 1676037725
transform 1 0 32292 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_349
timestamp 1676037725
transform 1 0 33212 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_355
timestamp 1676037725
transform 1 0 33764 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1676037725
transform 1 0 34408 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_376
timestamp 1676037725
transform 1 0 35696 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_386
timestamp 1676037725
transform 1 0 36616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_390
timestamp 1676037725
transform 1 0 36984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_399
timestamp 1676037725
transform 1 0 37812 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_407
timestamp 1676037725
transform 1 0 38548 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_412
timestamp 1676037725
transform 1 0 39008 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_440
timestamp 1676037725
transform 1 0 41584 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_452
timestamp 1676037725
transform 1 0 42688 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_460
timestamp 1676037725
transform 1 0 43424 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_35
timestamp 1676037725
transform 1 0 4324 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1676037725
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_68
timestamp 1676037725
transform 1 0 7360 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_76
timestamp 1676037725
transform 1 0 8096 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_88
timestamp 1676037725
transform 1 0 9200 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1676037725
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_124
timestamp 1676037725
transform 1 0 12512 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_130
timestamp 1676037725
transform 1 0 13064 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_152
timestamp 1676037725
transform 1 0 15088 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1676037725
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_177
timestamp 1676037725
transform 1 0 17388 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_188
timestamp 1676037725
transform 1 0 18400 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_200
timestamp 1676037725
transform 1 0 19504 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_212
timestamp 1676037725
transform 1 0 20608 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_232
timestamp 1676037725
transform 1 0 22448 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_240
timestamp 1676037725
transform 1 0 23184 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_260
timestamp 1676037725
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_272
timestamp 1676037725
transform 1 0 26128 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1676037725
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1676037725
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_341
timestamp 1676037725
transform 1 0 32476 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_354
timestamp 1676037725
transform 1 0 33672 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_376
timestamp 1676037725
transform 1 0 35696 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_388
timestamp 1676037725
transform 1 0 36800 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_412
timestamp 1676037725
transform 1 0 39008 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_424
timestamp 1676037725
transform 1 0 40112 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_436
timestamp 1676037725
transform 1 0 41216 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_460
timestamp 1676037725
transform 1 0 43424 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_54
timestamp 1676037725
transform 1 0 6072 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_67
timestamp 1676037725
transform 1 0 7268 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_79
timestamp 1676037725
transform 1 0 8372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_99
timestamp 1676037725
transform 1 0 10212 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_105
timestamp 1676037725
transform 1 0 10764 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_122
timestamp 1676037725
transform 1 0 12328 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_134
timestamp 1676037725
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_154
timestamp 1676037725
transform 1 0 15272 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_162
timestamp 1676037725
transform 1 0 16008 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_167
timestamp 1676037725
transform 1 0 16468 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1676037725
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_205
timestamp 1676037725
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_211
timestamp 1676037725
transform 1 0 20516 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_217
timestamp 1676037725
transform 1 0 21068 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_239
timestamp 1676037725
transform 1 0 23092 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_261
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_275
timestamp 1676037725
transform 1 0 26404 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_287
timestamp 1676037725
transform 1 0 27508 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_294
timestamp 1676037725
transform 1 0 28152 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1676037725
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_322
timestamp 1676037725
transform 1 0 30728 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_329
timestamp 1676037725
transform 1 0 31372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_346
timestamp 1676037725
transform 1 0 32936 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_355
timestamp 1676037725
transform 1 0 33764 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1676037725
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_371
timestamp 1676037725
transform 1 0 35236 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_382
timestamp 1676037725
transform 1 0 36248 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_394
timestamp 1676037725
transform 1 0 37352 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_402
timestamp 1676037725
transform 1 0 38088 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_408
timestamp 1676037725
transform 1 0 38640 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_430
timestamp 1676037725
transform 1 0 40664 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_442
timestamp 1676037725
transform 1 0 41768 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_460
timestamp 1676037725
transform 1 0 43424 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_87
timestamp 1676037725
transform 1 0 9108 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_91
timestamp 1676037725
transform 1 0 9476 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_101
timestamp 1676037725
transform 1 0 10396 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 1676037725
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_124
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_136
timestamp 1676037725
transform 1 0 13616 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_155
timestamp 1676037725
transform 1 0 15364 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_159
timestamp 1676037725
transform 1 0 15732 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 1676037725
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_180
timestamp 1676037725
transform 1 0 17664 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_190
timestamp 1676037725
transform 1 0 18584 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_198
timestamp 1676037725
transform 1 0 19320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_219
timestamp 1676037725
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_229
timestamp 1676037725
transform 1 0 22172 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_233
timestamp 1676037725
transform 1 0 22540 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_245
timestamp 1676037725
transform 1 0 23644 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_258
timestamp 1676037725
transform 1 0 24840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_268
timestamp 1676037725
transform 1 0 25760 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_272
timestamp 1676037725
transform 1 0 26128 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1676037725
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_292
timestamp 1676037725
transform 1 0 27968 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_304
timestamp 1676037725
transform 1 0 29072 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_320
timestamp 1676037725
transform 1 0 30544 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_333
timestamp 1676037725
transform 1 0 31740 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_348
timestamp 1676037725
transform 1 0 33120 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_357
timestamp 1676037725
transform 1 0 33948 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_366
timestamp 1676037725
transform 1 0 34776 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 1676037725
transform 1 0 36984 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_402
timestamp 1676037725
transform 1 0 38088 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_408
timestamp 1676037725
transform 1 0 38640 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_414
timestamp 1676037725
transform 1 0 39192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_423
timestamp 1676037725
transform 1 0 40020 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_446
timestamp 1676037725
transform 1 0 42136 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_453
timestamp 1676037725
transform 1 0 42780 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_460
timestamp 1676037725
transform 1 0 43424 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_47
timestamp 1676037725
transform 1 0 5428 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_64
timestamp 1676037725
transform 1 0 6992 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_76
timestamp 1676037725
transform 1 0 8096 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_103
timestamp 1676037725
transform 1 0 10580 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_115
timestamp 1676037725
transform 1 0 11684 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_138
timestamp 1676037725
transform 1 0 13800 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_170
timestamp 1676037725
transform 1 0 16744 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_202
timestamp 1676037725
transform 1 0 19688 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_214
timestamp 1676037725
transform 1 0 20792 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_218
timestamp 1676037725
transform 1 0 21160 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_240
timestamp 1676037725
transform 1 0 23184 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_246
timestamp 1676037725
transform 1 0 23736 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_275
timestamp 1676037725
transform 1 0 26404 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_292
timestamp 1676037725
transform 1 0 27968 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_306
timestamp 1676037725
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_317
timestamp 1676037725
transform 1 0 30268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_341
timestamp 1676037725
transform 1 0 32476 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_351
timestamp 1676037725
transform 1 0 33396 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_360
timestamp 1676037725
transform 1 0 34224 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_384
timestamp 1676037725
transform 1 0 36432 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_396
timestamp 1676037725
transform 1 0 37536 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_417
timestamp 1676037725
transform 1 0 39468 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_440
timestamp 1676037725
transform 1 0 41584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_446
timestamp 1676037725
transform 1 0 42136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_450
timestamp 1676037725
transform 1 0 42504 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_460
timestamp 1676037725
transform 1 0 43424 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_11
timestamp 1676037725
transform 1 0 2116 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_22
timestamp 1676037725
transform 1 0 3128 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_29
timestamp 1676037725
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_41
timestamp 1676037725
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_54
timestamp 1676037725
transform 1 0 6072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_68
timestamp 1676037725
transform 1 0 7360 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_80
timestamp 1676037725
transform 1 0 8464 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_85
timestamp 1676037725
transform 1 0 8924 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_102
timestamp 1676037725
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_138
timestamp 1676037725
transform 1 0 13800 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_141
timestamp 1676037725
transform 1 0 14076 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_152
timestamp 1676037725
transform 1 0 15088 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1676037725
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_180
timestamp 1676037725
transform 1 0 17664 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_197
timestamp 1676037725
transform 1 0 19228 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_209
timestamp 1676037725
transform 1 0 20332 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_253
timestamp 1676037725
transform 1 0 24380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_267
timestamp 1676037725
transform 1 0 25668 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_289
timestamp 1676037725
transform 1 0 27692 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_302
timestamp 1676037725
transform 1 0 28888 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_309
timestamp 1676037725
transform 1 0 29532 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_321
timestamp 1676037725
transform 1 0 30636 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1676037725
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_343
timestamp 1676037725
transform 1 0 32660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_355
timestamp 1676037725
transform 1 0 33764 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_363
timestamp 1676037725
transform 1 0 34500 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_365
timestamp 1676037725
transform 1 0 34684 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_377
timestamp 1676037725
transform 1 0 35788 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1676037725
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_421
timestamp 1676037725
transform 1 0 39836 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_433
timestamp 1676037725
transform 1 0 40940 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_439
timestamp 1676037725
transform 1 0 41492 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_446
timestamp 1676037725
transform 1 0 42136 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_460
timestamp 1676037725
transform 1 0 43424 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 43884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 43884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 43884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 43884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 43884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 43884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 43884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 43884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 43884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 43884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 43884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 43884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 43884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 43884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 43884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 43884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 43884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 43884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 43884 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 43884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 43884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 43884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 43884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 43884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 43884 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 43884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 43884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 43884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 43884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 43884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 43884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 43884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 43884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 43884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 43884 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 43884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 43884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 43884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 43884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 43884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 43884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 43884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 43884 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 43884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 43884 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 43884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 43884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 43884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 43884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 43884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 43884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 43884 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 43884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 43884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 43884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 43884 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 43884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 43884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 43884 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 34592 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34132 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1676037725
transform 1 0 32292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1676037725
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1676037725
transform -1 0 20424 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1676037725
transform 1 0 19044 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1676037725
transform 1 0 18768 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33028 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_8  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_8  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8832 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1676037725
transform 1 0 14352 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10212 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0846_
timestamp 1676037725
transform 1 0 9108 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1676037725
transform -1 0 9660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34776 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0849_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31740 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25668 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30544 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27876 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 33948 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0855_
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31280 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30084 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31832 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1676037725
transform 1 0 32384 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform -1 0 27876 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0862_
timestamp 1676037725
transform -1 0 34224 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31372 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30544 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0865_
timestamp 1676037725
transform 1 0 30820 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0866_
timestamp 1676037725
transform -1 0 24104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0867_
timestamp 1676037725
transform -1 0 30728 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_4  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0869_
timestamp 1676037725
transform -1 0 29624 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31556 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0873_
timestamp 1676037725
transform -1 0 31832 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25024 0 -1 40256
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1676037725
transform -1 0 25760 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34500 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0878_
timestamp 1676037725
transform -1 0 34408 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0879_
timestamp 1676037725
transform -1 0 28152 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0880_
timestamp 1676037725
transform 1 0 27416 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0881_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0882_
timestamp 1676037725
transform 1 0 29440 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1676037725
transform 1 0 27232 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0884_
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1676037725
transform 1 0 30176 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29992 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0887_
timestamp 1676037725
transform -1 0 30544 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1676037725
transform -1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0889_
timestamp 1676037725
transform -1 0 31740 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1676037725
transform 1 0 33764 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31832 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0892_
timestamp 1676037725
transform 1 0 36156 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1676037725
transform 1 0 42228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0894_
timestamp 1676037725
transform 1 0 32292 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0895_
timestamp 1676037725
transform -1 0 22172 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1676037725
transform -1 0 28796 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0897_
timestamp 1676037725
transform -1 0 23552 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0898_
timestamp 1676037725
transform -1 0 26404 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1676037725
transform -1 0 26680 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0900_
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0901_
timestamp 1676037725
transform 1 0 20792 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0903_
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0904_
timestamp 1676037725
transform -1 0 27876 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0905_
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1676037725
transform -1 0 28244 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30544 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0908_
timestamp 1676037725
transform -1 0 29808 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0909_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29256 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27968 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1676037725
transform -1 0 25576 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1676037725
transform 1 0 27324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0915_
timestamp 1676037725
transform 1 0 27140 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24196 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0917_
timestamp 1676037725
transform 1 0 32292 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1676037725
transform -1 0 31372 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 29716 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0920_
timestamp 1676037725
transform 1 0 22908 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28244 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1676037725
transform 1 0 29716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1676037725
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0925_
timestamp 1676037725
transform 1 0 24196 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26680 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22356 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__o22ai_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25760 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0930_
timestamp 1676037725
transform -1 0 30452 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0931_
timestamp 1676037725
transform -1 0 31740 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0932_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33672 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27968 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_4  _0936_
timestamp 1676037725
transform 1 0 21988 0 1 32640
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21988 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23276 0 -1 33728
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0939_
timestamp 1676037725
transform 1 0 27692 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1676037725
transform 1 0 33764 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 35972 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _0945_
timestamp 1676037725
transform 1 0 31924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _0946_
timestamp 1676037725
transform 1 0 31924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__a221oi_4  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0948_
timestamp 1676037725
transform -1 0 33120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0949_
timestamp 1676037725
transform -1 0 29164 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0950_
timestamp 1676037725
transform 1 0 26404 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0951_
timestamp 1676037725
transform -1 0 30544 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform -1 0 27968 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0953_
timestamp 1676037725
transform -1 0 30544 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _0954_
timestamp 1676037725
transform -1 0 30728 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29256 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1676037725
transform -1 0 30176 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _0957_
timestamp 1676037725
transform 1 0 30084 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 33488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0959_
timestamp 1676037725
transform 1 0 28152 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform -1 0 24840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1676037725
transform 1 0 34132 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1676037725
transform -1 0 36340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0963_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1676037725
transform -1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0965_
timestamp 1676037725
transform -1 0 33304 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0966_
timestamp 1676037725
transform 1 0 27140 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0967_
timestamp 1676037725
transform 1 0 25576 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0968_
timestamp 1676037725
transform -1 0 26404 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1676037725
transform 1 0 28152 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0973_
timestamp 1676037725
transform 1 0 27324 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28152 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25668 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25944 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _0978_
timestamp 1676037725
transform -1 0 23276 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0980_
timestamp 1676037725
transform -1 0 23552 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1676037725
transform -1 0 24196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0982_
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1676037725
transform -1 0 24104 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1676037725
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1676037725
transform -1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1676037725
transform 1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0990_
timestamp 1676037725
transform 1 0 14628 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0994_
timestamp 1676037725
transform -1 0 19872 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1676037725
transform -1 0 17572 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0996_
timestamp 1676037725
transform -1 0 17112 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1676037725
transform -1 0 36340 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0999_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32936 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1002_
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1003_
timestamp 1676037725
transform -1 0 27600 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1004_
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1005_
timestamp 1676037725
transform -1 0 25944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1676037725
transform -1 0 25300 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1008_
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1009_
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1676037725
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1676037725
transform 1 0 22724 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1012_
timestamp 1676037725
transform -1 0 23368 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1676037725
transform 1 0 21988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1016_
timestamp 1676037725
transform -1 0 36340 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1017_
timestamp 1676037725
transform 1 0 37352 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1676037725
transform -1 0 33120 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1019_
timestamp 1676037725
transform 1 0 33304 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1020_
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1021_
timestamp 1676037725
transform -1 0 28980 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1676037725
transform -1 0 24104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1023_
timestamp 1676037725
transform -1 0 24104 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1676037725
transform -1 0 23092 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1025_
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1026_
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1028_
timestamp 1676037725
transform 1 0 22356 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1676037725
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1676037725
transform -1 0 23460 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1031_
timestamp 1676037725
transform -1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1032_
timestamp 1676037725
transform 1 0 23184 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 1676037725
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1676037725
transform -1 0 26128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1035_
timestamp 1676037725
transform -1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _1036_
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1676037725
transform -1 0 31924 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1038_
timestamp 1676037725
transform -1 0 30544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1039_
timestamp 1676037725
transform 1 0 29624 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1040_
timestamp 1676037725
transform -1 0 27876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1676037725
transform -1 0 25944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1042_
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1676037725
transform -1 0 25116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 1676037725
transform -1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1676037725
transform 1 0 25576 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1046_
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1047_
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1048_
timestamp 1676037725
transform -1 0 21160 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1676037725
transform -1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1676037725
transform -1 0 29256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1676037725
transform 1 0 30820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1052_
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1676037725
transform -1 0 31740 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1054_
timestamp 1676037725
transform 1 0 31004 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1055_
timestamp 1676037725
transform 1 0 30636 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1056_
timestamp 1676037725
transform -1 0 27968 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1676037725
transform -1 0 21160 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 1676037725
transform 1 0 19872 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1059_
timestamp 1676037725
transform -1 0 20516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1676037725
transform 1 0 19504 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1063_
timestamp 1676037725
transform -1 0 20424 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1066_
timestamp 1676037725
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1676037725
transform 1 0 26864 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1676037725
transform 1 0 26312 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1069_
timestamp 1676037725
transform -1 0 28796 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1676037725
transform -1 0 30360 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1071_
timestamp 1676037725
transform 1 0 29716 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1072_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1073_
timestamp 1676037725
transform -1 0 21528 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1075_
timestamp 1676037725
transform -1 0 23552 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _1076_
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1077_
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21528 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _1079_
timestamp 1676037725
transform -1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1080_
timestamp 1676037725
transform -1 0 20148 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1676037725
transform 1 0 20516 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1082_
timestamp 1676037725
transform -1 0 20148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1676037725
transform -1 0 21988 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1676037725
transform 1 0 22264 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1085_
timestamp 1676037725
transform 1 0 22356 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1676037725
transform 1 0 24656 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1087_
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25760 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1089_
timestamp 1676037725
transform -1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1090_
timestamp 1676037725
transform -1 0 19688 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1676037725
transform -1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1092_
timestamp 1676037725
transform -1 0 17940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _1093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19596 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _1094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _1095_
timestamp 1676037725
transform -1 0 18952 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1096_
timestamp 1676037725
transform -1 0 18952 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _1097_
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1098_
timestamp 1676037725
transform -1 0 21252 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1099_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__o211ai_4  _1104_
timestamp 1676037725
transform -1 0 21160 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1105_
timestamp 1676037725
transform -1 0 19964 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1106_
timestamp 1676037725
transform -1 0 21528 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1676037725
transform 1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1108_
timestamp 1676037725
transform 1 0 21804 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17848 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__o211ai_4  _1110_
timestamp 1676037725
transform -1 0 18400 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1676037725
transform 1 0 30360 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1676037725
transform -1 0 31832 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1113_
timestamp 1676037725
transform 1 0 31096 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1676037725
transform -1 0 31188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1676037725
transform -1 0 31280 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1116_
timestamp 1676037725
transform 1 0 30176 0 -1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _1117_
timestamp 1676037725
transform -1 0 27600 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1676037725
transform -1 0 22540 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1120_
timestamp 1676037725
transform -1 0 21712 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1676037725
transform 1 0 19596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1122_
timestamp 1676037725
transform -1 0 17204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17388 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1676037725
transform -1 0 16928 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1126_
timestamp 1676037725
transform -1 0 16376 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1130_
timestamp 1676037725
transform -1 0 27784 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1676037725
transform -1 0 18952 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1132_
timestamp 1676037725
transform -1 0 23552 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1133_
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1676037725
transform 1 0 14352 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1676037725
transform -1 0 15548 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1138_
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1676037725
transform -1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1140_
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1141_
timestamp 1676037725
transform -1 0 15456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1676037725
transform -1 0 14720 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1143_
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1145_
timestamp 1676037725
transform 1 0 14720 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1148_
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17480 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1151_
timestamp 1676037725
transform 1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1676037725
transform -1 0 35052 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1153_
timestamp 1676037725
transform 1 0 33488 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1154_
timestamp 1676037725
transform -1 0 33764 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1155_
timestamp 1676037725
transform -1 0 35604 0 -1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _1156_
timestamp 1676037725
transform -1 0 35328 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1157_
timestamp 1676037725
transform 1 0 31188 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__o31ai_4  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_8  _1159_
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1676037725
transform 1 0 33764 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1161_
timestamp 1676037725
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1676037725
transform 1 0 31096 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1676037725
transform 1 0 34040 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1164_
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1676037725
transform 1 0 26772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1166_
timestamp 1676037725
transform -1 0 32200 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1676037725
transform -1 0 31832 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1676037725
transform -1 0 33304 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1676037725
transform 1 0 33304 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32936 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35052 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1172_
timestamp 1676037725
transform -1 0 34224 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_2  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33764 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1174_
timestamp 1676037725
transform -1 0 34408 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1676037725
transform 1 0 33856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1676037725
transform 1 0 35236 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1676037725
transform 1 0 36248 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1178_
timestamp 1676037725
transform -1 0 35420 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1676037725
transform 1 0 33764 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _1180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34960 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_2  _1181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34960 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1676037725
transform 1 0 36156 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34040 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1676037725
transform 1 0 38640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1185_
timestamp 1676037725
transform 1 0 38824 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1676037725
transform 1 0 39376 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1187_
timestamp 1676037725
transform 1 0 39376 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1188_
timestamp 1676037725
transform 1 0 38916 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1189_
timestamp 1676037725
transform -1 0 39560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1676037725
transform 1 0 40112 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1191_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1192_
timestamp 1676037725
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1193_
timestamp 1676037725
transform 1 0 39652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1676037725
transform 1 0 40296 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp 1676037725
transform 1 0 40204 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1196_
timestamp 1676037725
transform 1 0 38824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1197_
timestamp 1676037725
transform 1 0 39836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1676037725
transform -1 0 40664 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1199_
timestamp 1676037725
transform 1 0 40204 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1200_
timestamp 1676037725
transform 1 0 38916 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1676037725
transform 1 0 40848 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1202_
timestamp 1676037725
transform 1 0 40020 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1676037725
transform 1 0 40112 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1676037725
transform -1 0 41216 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1205_
timestamp 1676037725
transform 1 0 34592 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1676037725
transform -1 0 38548 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1676037725
transform 1 0 35236 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1209_
timestamp 1676037725
transform -1 0 38364 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1210_
timestamp 1676037725
transform 1 0 36800 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1676037725
transform 1 0 37628 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1676037725
transform -1 0 39100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1676037725
transform -1 0 39744 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1676037725
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1216_
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1676037725
transform 1 0 38088 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1218_
timestamp 1676037725
transform -1 0 36708 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1220_
timestamp 1676037725
transform 1 0 37904 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1676037725
transform -1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1676037725
transform 1 0 38548 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1223_
timestamp 1676037725
transform 1 0 36708 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1224_
timestamp 1676037725
transform 1 0 37444 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1225_
timestamp 1676037725
transform 1 0 40020 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1226_
timestamp 1676037725
transform 1 0 36616 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1227_
timestamp 1676037725
transform 1 0 37444 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1228_
timestamp 1676037725
transform -1 0 39008 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1676037725
transform 1 0 38640 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1230_
timestamp 1676037725
transform -1 0 39284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1231_
timestamp 1676037725
transform 1 0 36248 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1232_
timestamp 1676037725
transform 1 0 37076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1676037725
transform 1 0 38364 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1676037725
transform 1 0 38732 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1676037725
transform 1 0 39560 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1236_
timestamp 1676037725
transform 1 0 35788 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1676037725
transform 1 0 36248 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp 1676037725
transform 1 0 37444 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1676037725
transform 1 0 22172 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1240_
timestamp 1676037725
transform -1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1676037725
transform -1 0 18952 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1676037725
transform 1 0 11684 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1243_
timestamp 1676037725
transform -1 0 7544 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1244_
timestamp 1676037725
transform 1 0 9108 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1245_
timestamp 1676037725
transform -1 0 15272 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1246_
timestamp 1676037725
transform -1 0 14904 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1247_
timestamp 1676037725
transform -1 0 11040 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1676037725
transform 1 0 6532 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1676037725
transform 1 0 6440 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1250_
timestamp 1676037725
transform 1 0 6532 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1676037725
transform 1 0 5704 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1252_
timestamp 1676037725
transform -1 0 6072 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _1253_
timestamp 1676037725
transform -1 0 7176 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1254_
timestamp 1676037725
transform 1 0 7544 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1676037725
transform 1 0 10396 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1256_
timestamp 1676037725
transform 1 0 9752 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _1257_
timestamp 1676037725
transform -1 0 12144 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1258_
timestamp 1676037725
transform 1 0 13524 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1676037725
transform 1 0 7912 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10396 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1261_
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1676037725
transform 1 0 32384 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1264_
timestamp 1676037725
transform -1 0 22816 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 1676037725
transform -1 0 22540 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1267_
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1268_
timestamp 1676037725
transform 1 0 14260 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1269_
timestamp 1676037725
transform -1 0 9292 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1270_
timestamp 1676037725
transform 1 0 12696 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1676037725
transform 1 0 14628 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1676037725
transform 1 0 17756 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1676037725
transform -1 0 20700 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1676037725
transform -1 0 10304 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1676037725
transform 1 0 16008 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1676037725
transform -1 0 8464 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1277_
timestamp 1676037725
transform 1 0 12052 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1676037725
transform -1 0 8372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1279_
timestamp 1676037725
transform 1 0 15456 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1280_
timestamp 1676037725
transform 1 0 14444 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1676037725
transform -1 0 24104 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1676037725
transform 1 0 28704 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1283_
timestamp 1676037725
transform -1 0 26312 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1676037725
transform 1 0 23184 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1285_
timestamp 1676037725
transform -1 0 26036 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1676037725
transform -1 0 25208 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1676037725
transform -1 0 25116 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1288_
timestamp 1676037725
transform 1 0 17480 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1289_
timestamp 1676037725
transform 1 0 27324 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1290_
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1676037725
transform 1 0 15364 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1676037725
transform -1 0 19872 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1294_
timestamp 1676037725
transform 1 0 12328 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1676037725
transform -1 0 17204 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1676037725
transform 1 0 14260 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1297_
timestamp 1676037725
transform 1 0 19596 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1676037725
transform -1 0 24288 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1676037725
transform -1 0 8096 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1676037725
transform -1 0 6256 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1301_
timestamp 1676037725
transform 1 0 12696 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1676037725
transform 1 0 14260 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1676037725
transform -1 0 18952 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1676037725
transform 1 0 20148 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1305_
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1306_
timestamp 1676037725
transform -1 0 13156 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1307_
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1676037725
transform 1 0 16836 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1309_
timestamp 1676037725
transform -1 0 16744 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1676037725
transform -1 0 13708 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_2  _1312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1313_
timestamp 1676037725
transform 1 0 26128 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1314_
timestamp 1676037725
transform 1 0 14260 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1315_
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19688 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 1676037725
transform -1 0 18308 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19044 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1676037725
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1676037725
transform 1 0 15456 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1321_
timestamp 1676037725
transform -1 0 11224 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1322_
timestamp 1676037725
transform -1 0 7728 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1676037725
transform 1 0 7084 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1324_
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1325_
timestamp 1676037725
transform -1 0 11960 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1326_
timestamp 1676037725
transform -1 0 9568 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1327_
timestamp 1676037725
transform -1 0 9476 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1329_
timestamp 1676037725
transform -1 0 17664 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1676037725
transform -1 0 13800 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1331_
timestamp 1676037725
transform -1 0 13800 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1332_
timestamp 1676037725
transform 1 0 13800 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1333_
timestamp 1676037725
transform 1 0 15732 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1334_
timestamp 1676037725
transform 1 0 27508 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27232 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1337_
timestamp 1676037725
transform 1 0 27140 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1338_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1339_
timestamp 1676037725
transform 1 0 24380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1676037725
transform 1 0 20792 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1676037725
transform 1 0 16192 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1676037725
transform 1 0 17020 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1344_
timestamp 1676037725
transform 1 0 15272 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1676037725
transform 1 0 22908 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1676037725
transform 1 0 18676 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1676037725
transform -1 0 21712 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1348_
timestamp 1676037725
transform 1 0 19412 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1676037725
transform 1 0 20148 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1350_
timestamp 1676037725
transform -1 0 27048 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1676037725
transform -1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1353_
timestamp 1676037725
transform 1 0 20792 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1676037725
transform -1 0 29072 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1355_
timestamp 1676037725
transform 1 0 28520 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1356_
timestamp 1676037725
transform -1 0 28980 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1676037725
transform -1 0 23736 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1676037725
transform 1 0 23460 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1676037725
transform -1 0 17112 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1676037725
transform 1 0 23552 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1361_
timestamp 1676037725
transform 1 0 16560 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29164 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1676037725
transform 1 0 29716 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1676037725
transform 1 0 23092 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1365_
timestamp 1676037725
transform 1 0 26864 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1366_
timestamp 1676037725
transform 1 0 24564 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1367_
timestamp 1676037725
transform 1 0 29348 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1368_
timestamp 1676037725
transform 1 0 34132 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _1369_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _1370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 36340 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_4  _1371_
timestamp 1676037725
transform 1 0 34868 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1372_
timestamp 1676037725
transform 1 0 35696 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1676037725
transform -1 0 34408 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1374_
timestamp 1676037725
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1375_
timestamp 1676037725
transform 1 0 34500 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1376_
timestamp 1676037725
transform -1 0 33396 0 1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1377_
timestamp 1676037725
transform 1 0 34868 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_4  _1378_
timestamp 1676037725
transform 1 0 30268 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1676037725
transform -1 0 35512 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1381_
timestamp 1676037725
transform 1 0 37444 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1382_
timestamp 1676037725
transform 1 0 35144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1383_
timestamp 1676037725
transform 1 0 33948 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1676037725
transform 1 0 38824 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1385_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1386_
timestamp 1676037725
transform -1 0 40664 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1387_
timestamp 1676037725
transform 1 0 37076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_
timestamp 1676037725
transform -1 0 37352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1389_
timestamp 1676037725
transform -1 0 38088 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1390_
timestamp 1676037725
transform 1 0 39008 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1391_
timestamp 1676037725
transform -1 0 38456 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1392_
timestamp 1676037725
transform -1 0 40756 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1676037725
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1394_
timestamp 1676037725
transform -1 0 38180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1395_
timestamp 1676037725
transform -1 0 40664 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 1676037725
transform 1 0 38548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1397_
timestamp 1676037725
transform -1 0 38272 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1398_
timestamp 1676037725
transform -1 0 39560 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1399_
timestamp 1676037725
transform 1 0 38640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1400_
timestamp 1676037725
transform -1 0 38272 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1676037725
transform -1 0 39376 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1402_
timestamp 1676037725
transform 1 0 38824 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1403_
timestamp 1676037725
transform -1 0 38180 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1404_
timestamp 1676037725
transform -1 0 40664 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1405_
timestamp 1676037725
transform -1 0 36064 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1406_
timestamp 1676037725
transform 1 0 34868 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1676037725
transform -1 0 36800 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1676037725
transform -1 0 36708 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 1676037725
transform 1 0 38732 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1410_
timestamp 1676037725
transform -1 0 39652 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1676037725
transform -1 0 40572 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 1676037725
transform 1 0 37904 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1413_
timestamp 1676037725
transform 1 0 40296 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 1676037725
transform 1 0 39100 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1676037725
transform 1 0 40388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 1676037725
transform 1 0 40020 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1417_
timestamp 1676037725
transform 1 0 40940 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 1676037725
transform 1 0 38916 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1676037725
transform 1 0 40112 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 1676037725
transform 1 0 38824 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1421_
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1676037725
transform 1 0 38916 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1676037725
transform 1 0 40020 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 33488 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _1425_
timestamp 1676037725
transform -1 0 33672 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 1676037725
transform 1 0 36064 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1676037725
transform 1 0 35052 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1676037725
transform 1 0 36064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1429_
timestamp 1676037725
transform 1 0 35328 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1676037725
transform 1 0 33488 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1431_
timestamp 1676037725
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1432_
timestamp 1676037725
transform -1 0 37168 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1676037725
transform -1 0 39100 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1436_
timestamp 1676037725
transform -1 0 38272 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 1676037725
transform -1 0 32936 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _1439_
timestamp 1676037725
transform 1 0 33488 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 1676037725
transform 1 0 32752 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1676037725
transform 1 0 32936 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1442_
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _1443_
timestamp 1676037725
transform -1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1444_
timestamp 1676037725
transform -1 0 34040 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1445_
timestamp 1676037725
transform -1 0 37720 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 1676037725
transform -1 0 35420 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1676037725
transform 1 0 35420 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1448_
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1676037725
transform 1 0 33764 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1450_
timestamp 1676037725
transform -1 0 37076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1451_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 36984 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1676037725
transform 1 0 34408 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1453_
timestamp 1676037725
transform 1 0 36064 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1454_
timestamp 1676037725
transform -1 0 35696 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _1455_
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27968 0 1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _1457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1458_
timestamp 1676037725
transform 1 0 27416 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1461_
timestamp 1676037725
transform 1 0 27048 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1462_
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1463_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1676037725
transform -1 0 30268 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1466_
timestamp 1676037725
transform -1 0 30452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1676037725
transform 1 0 30452 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1676037725
transform -1 0 28336 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1469_
timestamp 1676037725
transform -1 0 29256 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1470_
timestamp 1676037725
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1471_
timestamp 1676037725
transform 1 0 28428 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27784 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1676037725
transform 1 0 25852 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1474_
timestamp 1676037725
transform 1 0 28704 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1475_
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1676037725
transform 1 0 31188 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1477_
timestamp 1676037725
transform 1 0 31464 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1478_
timestamp 1676037725
transform 1 0 32936 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1479_
timestamp 1676037725
transform -1 0 31832 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1676037725
transform 1 0 33304 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1482_
timestamp 1676037725
transform 1 0 27968 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1676037725
transform -1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1676037725
transform 1 0 28796 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1485_
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31832 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1676037725
transform 1 0 32752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1676037725
transform 1 0 30912 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1676037725
transform 1 0 28428 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1490_
timestamp 1676037725
transform -1 0 30084 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1491_
timestamp 1676037725
transform -1 0 30544 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1492_
timestamp 1676037725
transform -1 0 31188 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1676037725
transform 1 0 32844 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1494_
timestamp 1676037725
transform -1 0 29808 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 1676037725
transform 1 0 27784 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1676037725
transform 1 0 29256 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1497_
timestamp 1676037725
transform 1 0 28336 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28980 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1676037725
transform -1 0 29256 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1500_
timestamp 1676037725
transform -1 0 31832 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1676037725
transform 1 0 22724 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1676037725
transform -1 0 40664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1676037725
transform 1 0 37812 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1676037725
transform -1 0 40480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1676037725
transform 1 0 37720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1676037725
transform 1 0 29900 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1509_
timestamp 1676037725
transform -1 0 33304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1510_
timestamp 1676037725
transform 1 0 26128 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1676037725
transform -1 0 34408 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1512_
timestamp 1676037725
transform 1 0 28244 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1513_
timestamp 1676037725
transform -1 0 28980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1676037725
transform 1 0 26956 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1515_
timestamp 1676037725
transform 1 0 26496 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1516_
timestamp 1676037725
transform 1 0 27508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1517_
timestamp 1676037725
transform -1 0 33764 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1518_
timestamp 1676037725
transform 1 0 33212 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1676037725
transform 1 0 34132 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1676037725
transform 1 0 41216 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1676037725
transform 1 0 42504 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1676037725
transform 1 0 42228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1676037725
transform 1 0 42596 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1676037725
transform 1 0 42596 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1676037725
transform 1 0 42596 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1527_
timestamp 1676037725
transform -1 0 18860 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1528_
timestamp 1676037725
transform -1 0 18584 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1529_
timestamp 1676037725
transform 1 0 17664 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1530_
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1676037725
transform 1 0 17756 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1676037725
transform 1 0 17296 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1676037725
transform 1 0 16192 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 1676037725
transform 1 0 23184 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1536_
timestamp 1676037725
transform -1 0 23184 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1537_
timestamp 1676037725
transform 1 0 23000 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1539_
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1540_
timestamp 1676037725
transform 1 0 25668 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1676037725
transform 1 0 25760 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1676037725
transform 1 0 24564 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1676037725
transform 1 0 22908 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1545_
timestamp 1676037725
transform 1 0 20884 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1676037725
transform 1 0 20700 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1676037725
transform 1 0 15824 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1676037725
transform 1 0 17940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1676037725
transform -1 0 17572 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1676037725
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1676037725
transform -1 0 15916 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1555_
timestamp 1676037725
transform 1 0 22908 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1556_
timestamp 1676037725
transform -1 0 23552 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1676037725
transform -1 0 23644 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1676037725
transform 1 0 23920 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1676037725
transform -1 0 21528 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1560_
timestamp 1676037725
transform 1 0 18032 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19044 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 1676037725
transform 1 0 11868 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1564_
timestamp 1676037725
transform 1 0 13340 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1565_
timestamp 1676037725
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1566_
timestamp 1676037725
transform -1 0 18768 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1676037725
transform -1 0 19596 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1568_
timestamp 1676037725
transform -1 0 18400 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1676037725
transform 1 0 6532 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1676037725
transform 1 0 5244 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1676037725
transform 1 0 9568 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1676037725
transform 1 0 14260 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1676037725
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1574_
timestamp 1676037725
transform 1 0 16836 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1676037725
transform 1 0 8372 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1676037725
transform 1 0 12972 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1676037725
transform -1 0 18492 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1578_
timestamp 1676037725
transform 1 0 17020 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1579_
timestamp 1676037725
transform -1 0 9016 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1580_
timestamp 1676037725
transform -1 0 8740 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1581_
timestamp 1676037725
transform -1 0 10488 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1676037725
transform -1 0 8832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1583_
timestamp 1676037725
transform -1 0 8648 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1676037725
transform -1 0 7728 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1586_
timestamp 1676037725
transform 1 0 6624 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1676037725
transform 1 0 10580 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1588_
timestamp 1676037725
transform -1 0 10948 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1676037725
transform 1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1590_
timestamp 1676037725
transform 1 0 8004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1591_
timestamp 1676037725
transform -1 0 9660 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1592_
timestamp 1676037725
transform 1 0 7268 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1593_
timestamp 1676037725
transform -1 0 7636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 1676037725
transform 1 0 6532 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1595_
timestamp 1676037725
transform -1 0 34408 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1596_
timestamp 1676037725
transform -1 0 10580 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1598_
timestamp 1676037725
transform -1 0 7820 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1599_
timestamp 1676037725
transform -1 0 7176 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1600_
timestamp 1676037725
transform 1 0 20240 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1676037725
transform -1 0 19964 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1602_
timestamp 1676037725
transform -1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1676037725
transform 1 0 6992 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1604_
timestamp 1676037725
transform 1 0 6072 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1676037725
transform 1 0 4600 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 1676037725
transform -1 0 9660 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1676037725
transform 1 0 9752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1676037725
transform 1 0 9108 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1609_
timestamp 1676037725
transform 1 0 6256 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1610_
timestamp 1676037725
transform 1 0 4876 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1676037725
transform -1 0 7268 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1612_
timestamp 1676037725
transform 1 0 5796 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1676037725
transform 1 0 10764 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1614_
timestamp 1676037725
transform -1 0 13616 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1615_
timestamp 1676037725
transform -1 0 11592 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1616_
timestamp 1676037725
transform 1 0 17480 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1617_
timestamp 1676037725
transform 1 0 6348 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1618_
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1619_
timestamp 1676037725
transform -1 0 5796 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1676037725
transform 1 0 4968 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1676037725
transform 1 0 4784 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp 1676037725
transform -1 0 7360 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1676037725
transform -1 0 7268 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1624_
timestamp 1676037725
transform -1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1626_
timestamp 1676037725
transform 1 0 9108 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1627_
timestamp 1676037725
transform 1 0 10672 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1676037725
transform -1 0 15272 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1630_
timestamp 1676037725
transform -1 0 9384 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1676037725
transform -1 0 8648 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1676037725
transform -1 0 8648 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1676037725
transform 1 0 11684 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 1676037725
transform 1 0 9844 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1676037725
transform 1 0 10580 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1636_
timestamp 1676037725
transform -1 0 13892 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1637_
timestamp 1676037725
transform -1 0 10856 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1638_
timestamp 1676037725
transform 1 0 12788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1639_
timestamp 1676037725
transform 1 0 9108 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1640_
timestamp 1676037725
transform -1 0 8740 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1641_
timestamp 1676037725
transform -1 0 11868 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1642_
timestamp 1676037725
transform 1 0 9844 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1643_
timestamp 1676037725
transform 1 0 10304 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1676037725
transform -1 0 12880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1645_
timestamp 1676037725
transform 1 0 9476 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1646_
timestamp 1676037725
transform 1 0 11684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1676037725
transform 1 0 10212 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1676037725
transform -1 0 9292 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1676037725
transform -1 0 9752 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1676037725
transform 1 0 10304 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1651_
timestamp 1676037725
transform 1 0 7728 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1652_
timestamp 1676037725
transform 1 0 11684 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1676037725
transform 1 0 14260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1676037725
transform 1 0 13800 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1676037725
transform 1 0 12052 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp 1676037725
transform 1 0 12788 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1657_
timestamp 1676037725
transform 1 0 11960 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1658_
timestamp 1676037725
transform -1 0 12788 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1676037725
transform 1 0 13156 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1676037725
transform -1 0 20056 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1676037725
transform 1 0 17664 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1663_
timestamp 1676037725
transform -1 0 36248 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1664_
timestamp 1676037725
transform 1 0 34868 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1676037725
transform 1 0 42596 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1676037725
transform 1 0 42596 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1676037725
transform 1 0 42596 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1676037725
transform 1 0 42596 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1676037725
transform 1 0 42596 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1676037725
transform 1 0 42596 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1676037725
transform 1 0 42596 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1673_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1676037725
transform 1 0 30452 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1676037725
transform 1 0 24472 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1676037725
transform 1 0 35512 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1676037725
transform 1 0 35420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1676037725
transform 1 0 35512 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1676037725
transform 1 0 35052 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1682_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1676037725
transform 1 0 40020 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1676037725
transform -1 0 40572 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1676037725
transform -1 0 39560 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1676037725
transform 1 0 37812 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1676037725
transform -1 0 31832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1676037725
transform -1 0 19688 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1676037725
transform 1 0 22264 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1676037725
transform -1 0 22448 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1676037725
transform 1 0 23828 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1676037725
transform 1 0 31556 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1697_
timestamp 1676037725
transform 1 0 17112 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21252 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21160 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1701_
timestamp 1676037725
transform -1 0 32476 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1676037725
transform 1 0 30084 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1676037725
transform 1 0 25208 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1676037725
transform 1 0 32476 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1676037725
transform 1 0 33028 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1676037725
transform 1 0 32292 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1676037725
transform 1 0 32384 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1676037725
transform 1 0 28704 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1676037725
transform 1 0 27324 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1676037725
transform 1 0 37444 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1676037725
transform 1 0 37536 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11960 0 1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1719_
timestamp 1676037725
transform 1 0 12144 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1721_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1722_
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1723_
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1724_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1725_
timestamp 1676037725
transform 1 0 23920 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1726_
timestamp 1676037725
transform 1 0 17020 0 1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1727_
timestamp 1676037725
transform 1 0 15732 0 1 22848
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1676037725
transform 1 0 10764 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1676037725
transform 1 0 10672 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 32752 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1731_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1732_
timestamp 1676037725
transform 1 0 36248 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1733_
timestamp 1676037725
transform 1 0 40020 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1734_
timestamp 1676037725
transform -1 0 42136 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1735_
timestamp 1676037725
transform -1 0 42136 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1736_
timestamp 1676037725
transform -1 0 42136 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1737_
timestamp 1676037725
transform -1 0 42044 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1676037725
transform -1 0 36800 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1676037725
transform -1 0 41492 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1676037725
transform 1 0 40020 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1741_
timestamp 1676037725
transform 1 0 39008 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1742_
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1743_
timestamp 1676037725
transform 1 0 40020 0 1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1744_
timestamp 1676037725
transform 1 0 40020 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1745_
timestamp 1676037725
transform 1 0 37904 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1676037725
transform -1 0 33764 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1676037725
transform 1 0 40664 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1676037725
transform 1 0 41768 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1676037725
transform 1 0 41860 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1676037725
transform 1 0 41768 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1676037725
transform 1 0 41952 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1676037725
transform 1 0 41952 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1676037725
transform 1 0 41860 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1754_
timestamp 1676037725
transform 1 0 15456 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1676037725
transform 1 0 20608 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1676037725
transform 1 0 24840 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1676037725
transform 1 0 22540 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1676037725
transform 1 0 20608 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1759_
timestamp 1676037725
transform -1 0 15824 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1760_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1676037725
transform 1 0 5520 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1676037725
transform 1 0 4600 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1676037725
transform 1 0 9108 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1676037725
transform 1 0 13892 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1676037725
transform 1 0 10856 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1676037725
transform -1 0 16744 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1676037725
transform 1 0 7636 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1676037725
transform 1 0 12328 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1770_
timestamp 1676037725
transform 1 0 16836 0 1 40256
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1676037725
transform 1 0 5244 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1676037725
transform 1 0 34224 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1676037725
transform 1 0 19320 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1676037725
transform 1 0 3956 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1676037725
transform 1 0 4048 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1676037725
transform 1 0 4140 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1676037725
transform -1 0 17112 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1778_
timestamp 1676037725
transform 1 0 4232 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1779_
timestamp 1676037725
transform 1 0 4048 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1780_
timestamp 1676037725
transform 1 0 4140 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1676037725
transform 1 0 5520 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1676037725
transform 1 0 14536 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1676037725
transform 1 0 10212 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1784_
timestamp 1676037725
transform 1 0 14444 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1785_
timestamp 1676037725
transform 1 0 7636 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1676037725
transform 1 0 9200 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1788_
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1789_
timestamp 1676037725
transform 1 0 11316 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1676037725
transform 1 0 9660 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1676037725
transform -1 0 9384 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1676037725
transform 1 0 9752 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1676037725
transform 1 0 7176 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1676037725
transform 1 0 12052 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1676037725
transform 1 0 11684 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1676037725
transform -1 0 15272 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1800_
timestamp 1676037725
transform 1 0 18124 0 -1 32640
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1676037725
transform 1 0 18124 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1676037725
transform 1 0 16836 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1676037725
transform 1 0 35512 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1806_
timestamp 1676037725
transform 1 0 34868 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1807_
timestamp 1676037725
transform -1 0 37904 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1808_
timestamp 1676037725
transform 1 0 41860 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1809_
timestamp 1676037725
transform 1 0 41492 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1810_
timestamp 1676037725
transform 1 0 41860 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1811_
timestamp 1676037725
transform 1 0 41860 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1812_
timestamp 1676037725
transform 1 0 41676 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1813_
timestamp 1676037725
transform 1 0 41768 0 1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1814_
timestamp 1676037725
transform 1 0 41860 0 1 40256
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1676037725
transform 1 0 30084 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1676037725
transform 1 0 34960 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1676037725
transform 1 0 35144 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1676037725
transform 1 0 28520 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1676037725
transform 1 0 26496 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1676037725
transform 1 0 27600 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1676037725
transform 1 0 39744 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1676037725
transform -1 0 41584 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1676037725
transform 1 0 39744 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1676037725
transform 1 0 37536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1676037725
transform -1 0 33028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26404 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12696 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform -1 0 11776 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform -1 0 17848 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform -1 0 12972 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform -1 0 12972 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform 1 0 17480 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform -1 0 18032 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform -1 0 30728 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform -1 0 30268 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform -1 0 35880 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform 1 0 34776 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform 1 0 37076 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 35972 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform -1 0 36432 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 37904 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42688 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 39560 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1676037725
transform -1 0 21896 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1676037725
transform -1 0 35696 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  fanout44
timestamp 1676037725
transform -1 0 30452 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout45
timestamp 1676037725
transform -1 0 25116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout46
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 1676037725
transform -1 0 16284 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1676037725
transform 1 0 11592 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1676037725
transform -1 0 31096 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1676037725
transform 1 0 36432 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1676037725
transform -1 0 10396 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout52
timestamp 1676037725
transform -1 0 35052 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout53
timestamp 1676037725
transform -1 0 9936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout54
timestamp 1676037725
transform -1 0 26680 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1676037725
transform 1 0 28980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout56
timestamp 1676037725
transform -1 0 13340 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout57
timestamp 1676037725
transform 1 0 18032 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 1676037725
transform 1 0 17480 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout59
timestamp 1676037725
transform 1 0 15824 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1676037725
transform -1 0 16468 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout61
timestamp 1676037725
transform 1 0 34868 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout62
timestamp 1676037725
transform 1 0 11684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout63
timestamp 1676037725
transform 1 0 19044 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout65
timestamp 1676037725
transform -1 0 25392 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout66
timestamp 1676037725
transform 1 0 26680 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout67
timestamp 1676037725
transform -1 0 31004 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1676037725
transform 1 0 28520 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout69
timestamp 1676037725
transform -1 0 36616 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout70
timestamp 1676037725
transform 1 0 37444 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout72
timestamp 1676037725
transform -1 0 33764 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout73
timestamp 1676037725
transform 1 0 11868 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout74
timestamp 1676037725
transform -1 0 31372 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout75
timestamp 1676037725
transform 1 0 33856 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout76
timestamp 1676037725
transform 1 0 33120 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 1676037725
transform 1 0 32660 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout78
timestamp 1676037725
transform -1 0 33672 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout79
timestamp 1676037725
transform -1 0 33212 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout80
timestamp 1676037725
transform -1 0 34408 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout81
timestamp 1676037725
transform -1 0 18032 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout82
timestamp 1676037725
transform 1 0 27140 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1676037725
transform 1 0 27140 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1676037725
transform 1 0 28704 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout85
timestamp 1676037725
transform 1 0 25208 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout86
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout87
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout88
timestamp 1676037725
transform -1 0 30268 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout89
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout90
timestamp 1676037725
transform -1 0 30636 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout91
timestamp 1676037725
transform 1 0 23092 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1676037725
transform 1 0 2300 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1676037725
transform -1 0 6072 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input4
timestamp 1676037725
transform -1 0 12604 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input5
timestamp 1676037725
transform 1 0 18032 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1676037725
transform 1 0 20700 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  input7
timestamp 1676037725
transform 1 0 24564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input8
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input11
timestamp 1676037725
transform 1 0 42596 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 41584 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 42872 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 42872 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 42872 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 42872 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1676037725
transform 1 0 42872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1676037725
transform 1 0 42872 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1676037725
transform 1 0 42872 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1676037725
transform 1 0 42872 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1676037725
transform 1 0 42872 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1676037725
transform 1 0 42872 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1676037725
transform 1 0 42872 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1676037725
transform 1 0 42872 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1676037725
transform 1 0 42872 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1676037725
transform 1 0 42872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1676037725
transform 1 0 41952 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp 1676037725
transform 1 0 42872 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp 1676037725
transform 1 0 42872 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp 1676037725
transform 1 0 42872 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp 1676037725
transform 1 0 42872 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp 1676037725
transform 1 0 42872 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp 1676037725
transform 1 0 42872 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp 1676037725
transform 1 0 42872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp 1676037725
transform 1 0 42872 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp 1676037725
transform 1 0 42872 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp 1676037725
transform 1 0 42872 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_92 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_93
timestamp 1676037725
transform 1 0 43148 0 -1 16320
box -38 -48 314 592
<< labels >>
flabel metal2 s 39026 44200 39082 45000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 2226 44200 2282 45000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 5906 44200 5962 45000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 9586 44200 9642 45000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 13266 44200 13322 45000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 16946 44200 17002 45000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 20626 44200 20682 45000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 24306 44200 24362 45000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 27986 44200 28042 45000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 31666 44200 31722 45000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 35346 44200 35402 45000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 44200 42576 45000 42696 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal3 s 44200 2184 45000 2304 0 FreeSans 480 0 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal3 s 44200 17144 45000 17264 0 FreeSans 480 0 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal3 s 44200 18640 45000 18760 0 FreeSans 480 0 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal3 s 44200 20136 45000 20256 0 FreeSans 480 0 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal3 s 44200 21632 45000 21752 0 FreeSans 480 0 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal3 s 44200 23128 45000 23248 0 FreeSans 480 0 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal3 s 44200 24624 45000 24744 0 FreeSans 480 0 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal3 s 44200 26120 45000 26240 0 FreeSans 480 0 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal3 s 44200 27616 45000 27736 0 FreeSans 480 0 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal3 s 44200 29112 45000 29232 0 FreeSans 480 0 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal3 s 44200 30608 45000 30728 0 FreeSans 480 0 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal3 s 44200 3680 45000 3800 0 FreeSans 480 0 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal3 s 44200 32104 45000 32224 0 FreeSans 480 0 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal3 s 44200 33600 45000 33720 0 FreeSans 480 0 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal3 s 44200 35096 45000 35216 0 FreeSans 480 0 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal3 s 44200 36592 45000 36712 0 FreeSans 480 0 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal3 s 44200 38088 45000 38208 0 FreeSans 480 0 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal3 s 44200 39584 45000 39704 0 FreeSans 480 0 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal3 s 44200 41080 45000 41200 0 FreeSans 480 0 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal3 s 44200 5176 45000 5296 0 FreeSans 480 0 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal3 s 44200 6672 45000 6792 0 FreeSans 480 0 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal3 s 44200 8168 45000 8288 0 FreeSans 480 0 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal3 s 44200 9664 45000 9784 0 FreeSans 480 0 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal3 s 44200 11160 45000 11280 0 FreeSans 480 0 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal3 s 44200 12656 45000 12776 0 FreeSans 480 0 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal3 s 44200 14152 45000 14272 0 FreeSans 480 0 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal3 s 44200 15648 45000 15768 0 FreeSans 480 0 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 42706 44200 42762 45000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 42480 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 42480 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 42480 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 45000
<< end >>
