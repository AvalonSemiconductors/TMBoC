magic
tech sky130B
magscale 1 2
timestamp 1680007197
<< viali >>
rect 8585 15657 8619 15691
rect 9321 15453 9355 15487
rect 10241 15453 10275 15487
rect 9137 15385 9171 15419
rect 10057 15385 10091 15419
rect 10333 15113 10367 15147
rect 9597 12801 9631 12835
rect 10241 12801 10275 12835
rect 10057 12665 10091 12699
rect 4068 11781 4102 11815
rect 7297 11781 7331 11815
rect 6561 11713 6595 11747
rect 7481 11713 7515 11747
rect 3801 11645 3835 11679
rect 6653 11645 6687 11679
rect 7665 11645 7699 11679
rect 5181 11509 5215 11543
rect 4261 11305 4295 11339
rect 5641 11101 5675 11135
rect 6101 11101 6135 11135
rect 5396 11033 5430 11067
rect 6193 11033 6227 11067
rect 5089 10761 5123 10795
rect 6745 10761 6779 10795
rect 7205 10693 7239 10727
rect 3709 10625 3743 10659
rect 3976 10625 4010 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 6561 10557 6595 10591
rect 6653 10557 6687 10591
rect 6285 10217 6319 10251
rect 7481 10217 7515 10251
rect 6193 10013 6227 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 6009 9469 6043 9503
rect 7021 9469 7055 9503
rect 5733 9401 5767 9435
rect 6653 9401 6687 9435
rect 5549 9333 5583 9367
rect 6561 9333 6595 9367
rect 5457 9129 5491 9163
rect 5365 9061 5399 9095
rect 10057 9061 10091 9095
rect 6193 8993 6227 9027
rect 3341 8925 3375 8959
rect 5917 8925 5951 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 4997 8857 5031 8891
rect 9597 8857 9631 8891
rect 10241 8857 10275 8891
rect 3249 8789 3283 8823
rect 6653 8789 6687 8823
rect 5641 8585 5675 8619
rect 5850 8517 5884 8551
rect 3065 8449 3099 8483
rect 3332 8449 3366 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 7021 8449 7055 8483
rect 7205 8449 7239 8483
rect 5365 8381 5399 8415
rect 5733 8381 5767 8415
rect 4445 8245 4479 8279
rect 6009 8245 6043 8279
rect 2789 8041 2823 8075
rect 7113 8041 7147 8075
rect 6653 7905 6687 7939
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 3341 7701 3375 7735
rect 5273 7701 5307 7735
rect 3065 7497 3099 7531
rect 6561 7497 6595 7531
rect 5181 7429 5215 7463
rect 4353 7361 4387 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 5273 7293 5307 7327
rect 5457 7293 5491 7327
rect 4813 7157 4847 7191
rect 5365 6953 5399 6987
rect 3985 6817 4019 6851
rect 4252 6749 4286 6783
rect 6377 6749 6411 6783
rect 6469 6613 6503 6647
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 6745 6069 6779 6103
rect 5365 5865 5399 5899
rect 6837 5865 6871 5899
rect 7481 5865 7515 5899
rect 6561 5797 6595 5831
rect 8493 5729 8527 5763
rect 3985 5661 4019 5695
rect 6377 5661 6411 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 8309 5661 8343 5695
rect 4252 5593 4286 5627
rect 7297 5593 7331 5627
rect 7497 5593 7531 5627
rect 10057 5593 10091 5627
rect 10241 5593 10275 5627
rect 7665 5525 7699 5559
rect 8125 5525 8159 5559
rect 9597 5525 9631 5559
rect 4905 5321 4939 5355
rect 7757 5321 7791 5355
rect 3525 5185 3559 5219
rect 3792 5185 3826 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 7941 5185 7975 5219
rect 8033 5185 8067 5219
rect 5641 4981 5675 5015
rect 6653 4981 6687 5015
rect 6377 4777 6411 4811
rect 6561 4777 6595 4811
rect 3985 4709 4019 4743
rect 5641 4709 5675 4743
rect 3157 4573 3191 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 6193 4505 6227 4539
rect 6409 4505 6443 4539
rect 3065 4437 3099 4471
rect 4169 4437 4203 4471
rect 6561 4233 6595 4267
rect 2421 4097 2455 4131
rect 3332 4097 3366 4131
rect 5273 4097 5307 4131
rect 6929 4097 6963 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 2513 4029 2547 4063
rect 3065 4029 3099 4063
rect 5365 4029 5399 4063
rect 5457 4029 5491 4063
rect 6837 4029 6871 4063
rect 4905 3961 4939 3995
rect 7389 3961 7423 3995
rect 4445 3893 4479 3927
rect 6745 3893 6779 3927
rect 4353 3689 4387 3723
rect 4261 3621 4295 3655
rect 7297 3621 7331 3655
rect 4445 3553 4479 3587
rect 4997 3553 5031 3587
rect 5457 3553 5491 3587
rect 5549 3553 5583 3587
rect 6352 3553 6386 3587
rect 6469 3553 6503 3587
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 2421 3485 2455 3519
rect 2973 3485 3007 3519
rect 3157 3485 3191 3519
rect 4169 3485 4203 3519
rect 7665 3485 7699 3519
rect 10149 3485 10183 3519
rect 3249 3417 3283 3451
rect 7573 3417 7607 3451
rect 2237 3349 2271 3383
rect 5181 3349 5215 3383
rect 6193 3349 6227 3383
rect 7481 3349 7515 3383
rect 7849 3349 7883 3383
rect 5917 3145 5951 3179
rect 6745 3145 6779 3179
rect 6837 3145 6871 3179
rect 2053 3077 2087 3111
rect 2789 3077 2823 3111
rect 4353 3077 4387 3111
rect 5825 3009 5859 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 9873 3009 9907 3043
rect 10149 2941 10183 2975
rect 1869 2873 1903 2907
rect 6561 2805 6595 2839
rect 9413 2805 9447 2839
rect 10057 2533 10091 2567
rect 2053 2397 2087 2431
rect 3249 2397 3283 2431
rect 4721 2397 4755 2431
rect 5917 2397 5951 2431
rect 6653 2397 6687 2431
rect 7849 2397 7883 2431
rect 9137 2397 9171 2431
rect 1777 2329 1811 2363
rect 3065 2329 3099 2363
rect 4445 2329 4479 2363
rect 5641 2329 5675 2363
rect 6929 2329 6963 2363
rect 8125 2329 8159 2363
rect 9413 2329 9447 2363
rect 10241 2329 10275 2363
<< metal1 >>
rect 1104 15802 10856 15824
rect 1104 15750 2169 15802
rect 2221 15750 2233 15802
rect 2285 15750 2297 15802
rect 2349 15750 2361 15802
rect 2413 15750 2425 15802
rect 2477 15750 4607 15802
rect 4659 15750 4671 15802
rect 4723 15750 4735 15802
rect 4787 15750 4799 15802
rect 4851 15750 4863 15802
rect 4915 15750 7045 15802
rect 7097 15750 7109 15802
rect 7161 15750 7173 15802
rect 7225 15750 7237 15802
rect 7289 15750 7301 15802
rect 7353 15750 9483 15802
rect 9535 15750 9547 15802
rect 9599 15750 9611 15802
rect 9663 15750 9675 15802
rect 9727 15750 9739 15802
rect 9791 15750 10856 15802
rect 1104 15728 10856 15750
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15688 8631 15691
rect 8938 15688 8944 15700
rect 8619 15660 8944 15688
rect 8619 15657 8631 15660
rect 8573 15651 8631 15657
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 8996 15456 9321 15484
rect 8996 15444 9002 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15484 10287 15487
rect 10318 15484 10324 15496
rect 10275 15456 10324 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10318 15444 10324 15456
rect 10376 15484 10382 15496
rect 11054 15484 11060 15496
rect 10376 15456 11060 15484
rect 10376 15444 10382 15456
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 9122 15376 9128 15428
rect 9180 15376 9186 15428
rect 9858 15376 9864 15428
rect 9916 15416 9922 15428
rect 10045 15419 10103 15425
rect 10045 15416 10057 15419
rect 9916 15388 10057 15416
rect 9916 15376 9922 15388
rect 10045 15385 10057 15388
rect 10091 15385 10103 15419
rect 10045 15379 10103 15385
rect 1104 15258 11016 15280
rect 1104 15206 3388 15258
rect 3440 15206 3452 15258
rect 3504 15206 3516 15258
rect 3568 15206 3580 15258
rect 3632 15206 3644 15258
rect 3696 15206 5826 15258
rect 5878 15206 5890 15258
rect 5942 15206 5954 15258
rect 6006 15206 6018 15258
rect 6070 15206 6082 15258
rect 6134 15206 8264 15258
rect 8316 15206 8328 15258
rect 8380 15206 8392 15258
rect 8444 15206 8456 15258
rect 8508 15206 8520 15258
rect 8572 15206 10702 15258
rect 10754 15206 10766 15258
rect 10818 15206 10830 15258
rect 10882 15206 10894 15258
rect 10946 15206 10958 15258
rect 11010 15206 11016 15258
rect 1104 15184 11016 15206
rect 10318 15104 10324 15156
rect 10376 15104 10382 15156
rect 1104 14714 10856 14736
rect 1104 14662 2169 14714
rect 2221 14662 2233 14714
rect 2285 14662 2297 14714
rect 2349 14662 2361 14714
rect 2413 14662 2425 14714
rect 2477 14662 4607 14714
rect 4659 14662 4671 14714
rect 4723 14662 4735 14714
rect 4787 14662 4799 14714
rect 4851 14662 4863 14714
rect 4915 14662 7045 14714
rect 7097 14662 7109 14714
rect 7161 14662 7173 14714
rect 7225 14662 7237 14714
rect 7289 14662 7301 14714
rect 7353 14662 9483 14714
rect 9535 14662 9547 14714
rect 9599 14662 9611 14714
rect 9663 14662 9675 14714
rect 9727 14662 9739 14714
rect 9791 14662 10856 14714
rect 1104 14640 10856 14662
rect 1104 14170 11016 14192
rect 1104 14118 3388 14170
rect 3440 14118 3452 14170
rect 3504 14118 3516 14170
rect 3568 14118 3580 14170
rect 3632 14118 3644 14170
rect 3696 14118 5826 14170
rect 5878 14118 5890 14170
rect 5942 14118 5954 14170
rect 6006 14118 6018 14170
rect 6070 14118 6082 14170
rect 6134 14118 8264 14170
rect 8316 14118 8328 14170
rect 8380 14118 8392 14170
rect 8444 14118 8456 14170
rect 8508 14118 8520 14170
rect 8572 14118 10702 14170
rect 10754 14118 10766 14170
rect 10818 14118 10830 14170
rect 10882 14118 10894 14170
rect 10946 14118 10958 14170
rect 11010 14118 11016 14170
rect 1104 14096 11016 14118
rect 1104 13626 10856 13648
rect 1104 13574 2169 13626
rect 2221 13574 2233 13626
rect 2285 13574 2297 13626
rect 2349 13574 2361 13626
rect 2413 13574 2425 13626
rect 2477 13574 4607 13626
rect 4659 13574 4671 13626
rect 4723 13574 4735 13626
rect 4787 13574 4799 13626
rect 4851 13574 4863 13626
rect 4915 13574 7045 13626
rect 7097 13574 7109 13626
rect 7161 13574 7173 13626
rect 7225 13574 7237 13626
rect 7289 13574 7301 13626
rect 7353 13574 9483 13626
rect 9535 13574 9547 13626
rect 9599 13574 9611 13626
rect 9663 13574 9675 13626
rect 9727 13574 9739 13626
rect 9791 13574 10856 13626
rect 1104 13552 10856 13574
rect 1104 13082 11016 13104
rect 1104 13030 3388 13082
rect 3440 13030 3452 13082
rect 3504 13030 3516 13082
rect 3568 13030 3580 13082
rect 3632 13030 3644 13082
rect 3696 13030 5826 13082
rect 5878 13030 5890 13082
rect 5942 13030 5954 13082
rect 6006 13030 6018 13082
rect 6070 13030 6082 13082
rect 6134 13030 8264 13082
rect 8316 13030 8328 13082
rect 8380 13030 8392 13082
rect 8444 13030 8456 13082
rect 8508 13030 8520 13082
rect 8572 13030 10702 13082
rect 10754 13030 10766 13082
rect 10818 13030 10830 13082
rect 10882 13030 10894 13082
rect 10946 13030 10958 13082
rect 11010 13030 11016 13082
rect 1104 13008 11016 13030
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10226 12832 10232 12844
rect 9631 12804 10232 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 7466 12656 7472 12708
rect 7524 12696 7530 12708
rect 10045 12699 10103 12705
rect 10045 12696 10057 12699
rect 7524 12668 10057 12696
rect 7524 12656 7530 12668
rect 10045 12665 10057 12668
rect 10091 12665 10103 12699
rect 10045 12659 10103 12665
rect 1104 12538 10856 12560
rect 1104 12486 2169 12538
rect 2221 12486 2233 12538
rect 2285 12486 2297 12538
rect 2349 12486 2361 12538
rect 2413 12486 2425 12538
rect 2477 12486 4607 12538
rect 4659 12486 4671 12538
rect 4723 12486 4735 12538
rect 4787 12486 4799 12538
rect 4851 12486 4863 12538
rect 4915 12486 7045 12538
rect 7097 12486 7109 12538
rect 7161 12486 7173 12538
rect 7225 12486 7237 12538
rect 7289 12486 7301 12538
rect 7353 12486 9483 12538
rect 9535 12486 9547 12538
rect 9599 12486 9611 12538
rect 9663 12486 9675 12538
rect 9727 12486 9739 12538
rect 9791 12486 10856 12538
rect 1104 12464 10856 12486
rect 1104 11994 11016 12016
rect 1104 11942 3388 11994
rect 3440 11942 3452 11994
rect 3504 11942 3516 11994
rect 3568 11942 3580 11994
rect 3632 11942 3644 11994
rect 3696 11942 5826 11994
rect 5878 11942 5890 11994
rect 5942 11942 5954 11994
rect 6006 11942 6018 11994
rect 6070 11942 6082 11994
rect 6134 11942 8264 11994
rect 8316 11942 8328 11994
rect 8380 11942 8392 11994
rect 8444 11942 8456 11994
rect 8508 11942 8520 11994
rect 8572 11942 10702 11994
rect 10754 11942 10766 11994
rect 10818 11942 10830 11994
rect 10882 11942 10894 11994
rect 10946 11942 10958 11994
rect 11010 11942 11016 11994
rect 1104 11920 11016 11942
rect 4056 11815 4114 11821
rect 4056 11781 4068 11815
rect 4102 11812 4114 11815
rect 7285 11815 7343 11821
rect 7285 11812 7297 11815
rect 4102 11784 7297 11812
rect 4102 11781 4114 11784
rect 4056 11775 4114 11781
rect 7285 11781 7297 11784
rect 7331 11781 7343 11815
rect 7285 11775 7343 11781
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 3786 11636 3792 11688
rect 3844 11636 3850 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 6687 11648 7665 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7653 11645 7665 11648
rect 7699 11676 7711 11679
rect 7742 11676 7748 11688
rect 7699 11648 7748 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5626 11540 5632 11552
rect 5215 11512 5632 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 6822 11540 6828 11552
rect 5684 11512 6828 11540
rect 5684 11500 5690 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 1104 11450 10856 11472
rect 1104 11398 2169 11450
rect 2221 11398 2233 11450
rect 2285 11398 2297 11450
rect 2349 11398 2361 11450
rect 2413 11398 2425 11450
rect 2477 11398 4607 11450
rect 4659 11398 4671 11450
rect 4723 11398 4735 11450
rect 4787 11398 4799 11450
rect 4851 11398 4863 11450
rect 4915 11398 7045 11450
rect 7097 11398 7109 11450
rect 7161 11398 7173 11450
rect 7225 11398 7237 11450
rect 7289 11398 7301 11450
rect 7353 11398 9483 11450
rect 9535 11398 9547 11450
rect 9599 11398 9611 11450
rect 9663 11398 9675 11450
rect 9727 11398 9739 11450
rect 9791 11398 10856 11450
rect 1104 11376 10856 11398
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 6546 11336 6552 11348
rect 4295 11308 6552 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 5552 11172 6132 11200
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 5552 11132 5580 11172
rect 6104 11141 6132 11172
rect 3844 11104 5580 11132
rect 5629 11135 5687 11141
rect 3844 11092 3850 11104
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 5384 11067 5442 11073
rect 5384 11033 5396 11067
rect 5430 11064 5442 11067
rect 5534 11064 5540 11076
rect 5430 11036 5540 11064
rect 5430 11033 5442 11036
rect 5384 11027 5442 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5644 11064 5672 11095
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 5644 11036 6193 11064
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6181 11027 6239 11033
rect 1104 10906 11016 10928
rect 1104 10854 3388 10906
rect 3440 10854 3452 10906
rect 3504 10854 3516 10906
rect 3568 10854 3580 10906
rect 3632 10854 3644 10906
rect 3696 10854 5826 10906
rect 5878 10854 5890 10906
rect 5942 10854 5954 10906
rect 6006 10854 6018 10906
rect 6070 10854 6082 10906
rect 6134 10854 8264 10906
rect 8316 10854 8328 10906
rect 8380 10854 8392 10906
rect 8444 10854 8456 10906
rect 8508 10854 8520 10906
rect 8572 10854 10702 10906
rect 10754 10854 10766 10906
rect 10818 10854 10830 10906
rect 10882 10854 10894 10906
rect 10946 10854 10958 10906
rect 11010 10854 11016 10906
rect 1104 10832 11016 10854
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 6454 10792 6460 10804
rect 5123 10764 6460 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 6454 10752 6460 10764
rect 6512 10792 6518 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6512 10764 6745 10792
rect 6512 10752 6518 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 7193 10727 7251 10733
rect 7193 10724 7205 10727
rect 5592 10696 7205 10724
rect 5592 10684 5598 10696
rect 7193 10693 7205 10696
rect 7239 10693 7251 10727
rect 7193 10687 7251 10693
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 3786 10656 3792 10668
rect 3743 10628 3792 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 3964 10659 4022 10665
rect 3964 10625 3976 10659
rect 4010 10656 4022 10659
rect 6730 10656 6736 10668
rect 4010 10628 6736 10656
rect 4010 10625 4022 10628
rect 3964 10619 4022 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6880 10628 6929 10656
rect 6880 10616 6886 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 9122 10656 9128 10668
rect 7064 10628 9128 10656
rect 7064 10616 7070 10628
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6328 10560 6561 10588
rect 6328 10548 6334 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 1104 10362 10856 10384
rect 1104 10310 2169 10362
rect 2221 10310 2233 10362
rect 2285 10310 2297 10362
rect 2349 10310 2361 10362
rect 2413 10310 2425 10362
rect 2477 10310 4607 10362
rect 4659 10310 4671 10362
rect 4723 10310 4735 10362
rect 4787 10310 4799 10362
rect 4851 10310 4863 10362
rect 4915 10310 7045 10362
rect 7097 10310 7109 10362
rect 7161 10310 7173 10362
rect 7225 10310 7237 10362
rect 7289 10310 7301 10362
rect 7353 10310 9483 10362
rect 9535 10310 9547 10362
rect 9599 10310 9611 10362
rect 9663 10310 9675 10362
rect 9727 10310 9739 10362
rect 9791 10310 10856 10362
rect 1104 10288 10856 10310
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6638 10248 6644 10260
rect 6319 10220 6644 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 6788 10220 7481 10248
rect 6788 10208 6794 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6362 10044 6368 10056
rect 6227 10016 6368 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 4580 9472 6009 9500
rect 4580 9460 4586 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 5718 9392 5724 9444
rect 5776 9392 5782 9444
rect 6012 9432 6040 9463
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6236 9472 7021 9500
rect 6236 9460 6242 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 6362 9432 6368 9444
rect 6012 9404 6368 9432
rect 6362 9392 6368 9404
rect 6420 9432 6426 9444
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6420 9404 6653 9432
rect 6420 9392 6426 9404
rect 6641 9401 6653 9404
rect 6687 9401 6699 9435
rect 6641 9395 6699 9401
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5408 9336 5549 9364
rect 5408 9324 5414 9336
rect 5537 9333 5549 9336
rect 5583 9364 5595 9367
rect 6086 9364 6092 9376
rect 5583 9336 6092 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6270 9160 6276 9172
rect 5491 9132 6276 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5353 9095 5411 9101
rect 5353 9092 5365 9095
rect 5040 9064 5365 9092
rect 5040 9052 5046 9064
rect 5353 9061 5365 9064
rect 5399 9092 5411 9095
rect 5718 9092 5724 9104
rect 5399 9064 5724 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 5718 9052 5724 9064
rect 5776 9052 5782 9104
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 7708 9064 10057 9092
rect 7708 9052 7714 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6546 9024 6552 9036
rect 6227 8996 6552 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8956 3387 8959
rect 3786 8956 3792 8968
rect 3375 8928 3792 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 4985 8891 5043 8897
rect 4985 8857 4997 8891
rect 5031 8888 5043 8891
rect 5074 8888 5080 8900
rect 5031 8860 5080 8888
rect 5031 8857 5043 8860
rect 4985 8851 5043 8857
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 5920 8888 5948 8919
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6362 8888 6368 8900
rect 5920 8860 6368 8888
rect 6362 8848 6368 8860
rect 6420 8848 6426 8900
rect 9585 8891 9643 8897
rect 9585 8857 9597 8891
rect 9631 8888 9643 8891
rect 10226 8888 10232 8900
rect 9631 8860 10232 8888
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3108 8792 3249 8820
rect 3108 8780 3114 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6604 8792 6653 8820
rect 6604 8780 6610 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6641 8783 6699 8789
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5132 8588 5641 8616
rect 5132 8576 5138 8588
rect 5629 8585 5641 8588
rect 5675 8616 5687 8619
rect 6178 8616 6184 8628
rect 5675 8588 6184 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 5838 8551 5896 8557
rect 5838 8548 5850 8551
rect 5776 8520 5850 8548
rect 5776 8508 5782 8520
rect 5838 8517 5850 8520
rect 5884 8517 5896 8551
rect 6914 8548 6920 8560
rect 5838 8511 5896 8517
rect 6748 8520 6920 8548
rect 3050 8440 3056 8492
rect 3108 8440 3114 8492
rect 6748 8489 6776 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 3320 8483 3378 8489
rect 3320 8449 3332 8483
rect 3366 8480 3378 8483
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 3366 8452 6561 8480
rect 3366 8449 3378 8452
rect 3320 8443 3378 8449
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6880 8452 7021 8480
rect 6880 8440 6886 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 7374 8480 7380 8492
rect 7239 8452 7380 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 5350 8372 5356 8424
rect 5408 8372 5414 8424
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 6638 8412 6644 8424
rect 5767 8384 6644 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 6638 8372 6644 8384
rect 6696 8412 6702 8424
rect 9858 8412 9864 8424
rect 6696 8384 9864 8412
rect 6696 8372 6702 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4522 8276 4528 8288
rect 4479 8248 4528 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 5994 8236 6000 8288
rect 6052 8236 6058 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7374 8072 7380 8084
rect 7147 8044 7380 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 2792 7936 2820 8032
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 6454 8004 6460 8016
rect 6328 7976 6460 8004
rect 6328 7964 6334 7976
rect 6454 7964 6460 7976
rect 6512 8004 6518 8016
rect 6512 7976 6960 8004
rect 6512 7964 6518 7976
rect 2792 7908 4016 7936
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3108 7840 3433 7868
rect 3108 7828 3114 7840
rect 3421 7837 3433 7840
rect 3467 7868 3479 7871
rect 3786 7868 3792 7880
rect 3467 7840 3792 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 3988 7877 4016 7908
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6052 7908 6653 7936
rect 6052 7896 6058 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 6454 7868 6460 7880
rect 6411 7840 6460 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6932 7877 6960 7976
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3878 7732 3884 7744
rect 3375 7704 3884 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 4396 7704 5273 7732
rect 4396 7692 4402 7704
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 3050 7488 3056 7540
rect 3108 7488 3114 7540
rect 6362 7488 6368 7540
rect 6420 7528 6426 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6420 7500 6561 7528
rect 6420 7488 6426 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 5166 7420 5172 7472
rect 5224 7460 5230 7472
rect 5224 7432 6684 7460
rect 5224 7420 5230 7432
rect 6656 7404 6684 7432
rect 4338 7352 4344 7404
rect 4396 7352 4402 7404
rect 5718 7392 5724 7404
rect 5276 7364 5724 7392
rect 5276 7336 5304 7364
rect 5718 7352 5724 7364
rect 5776 7392 5782 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5776 7364 6561 7392
rect 5776 7352 5782 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6696 7364 6745 7392
rect 6696 7352 6702 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5442 7284 5448 7336
rect 5500 7284 5506 7336
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4304 7160 4813 7188
rect 4304 7148 4310 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 4801 7151 4859 7157
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5353 6987 5411 6993
rect 5353 6984 5365 6987
rect 5316 6956 5365 6984
rect 5316 6944 5322 6956
rect 5353 6953 5365 6956
rect 5399 6953 5411 6987
rect 5353 6947 5411 6953
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3936 6820 3985 6848
rect 3936 6808 3942 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4246 6789 4252 6792
rect 4240 6780 4252 6789
rect 4207 6752 4252 6780
rect 4240 6743 4252 6752
rect 4246 6740 4252 6743
rect 4304 6740 4310 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5684 6752 6377 6780
rect 5684 6740 5690 6752
rect 6365 6749 6377 6752
rect 6411 6780 6423 6783
rect 6638 6780 6644 6792
rect 6411 6752 6644 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6546 6644 6552 6656
rect 6503 6616 6552 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6328 6276 6561 6304
rect 6328 6264 6334 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 6914 6304 6920 6316
rect 6788 6276 6920 6304
rect 6788 6264 6794 6276
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 6730 6060 6736 6112
rect 6788 6060 6794 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5132 5868 5365 5896
rect 5132 5856 5138 5868
rect 5353 5865 5365 5868
rect 5399 5896 5411 5899
rect 6362 5896 6368 5908
rect 5399 5868 6368 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 6822 5856 6828 5908
rect 6880 5856 6886 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 7742 5896 7748 5908
rect 7515 5868 7748 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 6730 5828 6736 5840
rect 6595 5800 6736 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 4580 5664 6377 5692
rect 4580 5652 4586 5664
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 6748 5692 6776 5788
rect 7760 5760 7788 5856
rect 8018 5760 8024 5772
rect 7760 5732 8024 5760
rect 8018 5720 8024 5732
rect 8076 5760 8082 5772
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8076 5732 8493 5760
rect 8076 5720 8082 5732
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 8481 5723 8539 5729
rect 8297 5695 8355 5701
rect 6748 5664 7420 5692
rect 4240 5627 4298 5633
rect 4240 5593 4252 5627
rect 4286 5624 4298 5627
rect 7190 5624 7196 5636
rect 4286 5596 7196 5624
rect 4286 5593 4298 5596
rect 4240 5587 4298 5593
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 7282 5584 7288 5636
rect 7340 5584 7346 5636
rect 7392 5624 7420 5664
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 7485 5627 7543 5633
rect 7485 5624 7497 5627
rect 7392 5596 7497 5624
rect 7485 5593 7497 5596
rect 7531 5593 7543 5627
rect 8312 5624 8340 5655
rect 10045 5627 10103 5633
rect 10045 5624 10057 5627
rect 8312 5596 10057 5624
rect 7485 5587 7543 5593
rect 10045 5593 10057 5596
rect 10091 5593 10103 5627
rect 10045 5587 10103 5593
rect 10226 5584 10232 5636
rect 10284 5584 10290 5636
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 7834 5556 7840 5568
rect 7699 5528 7840 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 9585 5559 9643 5565
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 10244 5556 10272 5584
rect 9631 5528 10272 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 4982 5352 4988 5364
rect 4939 5324 4988 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 4982 5312 4988 5324
rect 5040 5352 5046 5364
rect 6822 5352 6828 5364
rect 5040 5324 6828 5352
rect 5040 5312 5046 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7248 5324 7757 5352
rect 7248 5312 7254 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 3970 5284 3976 5296
rect 3528 5256 3976 5284
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3528 5225 3556 5256
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 8110 5284 8116 5296
rect 4126 5256 8116 5284
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3200 5188 3525 5216
rect 3200 5176 3206 5188
rect 3513 5185 3525 5188
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 3780 5219 3838 5225
rect 3780 5185 3792 5219
rect 3826 5216 3838 5219
rect 4126 5216 4154 5256
rect 8110 5244 8116 5256
rect 8168 5244 8174 5296
rect 3826 5188 4154 5216
rect 5813 5219 5871 5225
rect 3826 5185 3838 5188
rect 3780 5179 3838 5185
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5828 5148 5856 5179
rect 5994 5176 6000 5228
rect 6052 5176 6058 5228
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6362 5216 6368 5228
rect 6144 5188 6368 5216
rect 6144 5176 6150 5188
rect 6362 5176 6368 5188
rect 6420 5216 6426 5228
rect 6730 5216 6736 5228
rect 6420 5188 6736 5216
rect 6420 5176 6426 5188
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6880 5188 6929 5216
rect 6880 5176 6886 5188
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 6546 5148 6552 5160
rect 5828 5120 6552 5148
rect 6546 5108 6552 5120
rect 6604 5148 6610 5160
rect 7282 5148 7288 5160
rect 6604 5120 7288 5148
rect 6604 5108 6610 5120
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6270 5080 6276 5092
rect 6052 5052 6276 5080
rect 6052 5040 6058 5052
rect 6270 5040 6276 5052
rect 6328 5040 6334 5092
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6914 5012 6920 5024
rect 6687 4984 6920 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 6365 4811 6423 4817
rect 6365 4777 6377 4811
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 3973 4743 4031 4749
rect 3973 4740 3985 4743
rect 2556 4712 3985 4740
rect 2556 4700 2562 4712
rect 3973 4709 3985 4712
rect 4019 4709 4031 4743
rect 3973 4703 4031 4709
rect 5629 4743 5687 4749
rect 5629 4709 5641 4743
rect 5675 4740 5687 4743
rect 6380 4740 6408 4771
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 6512 4780 6561 4808
rect 6512 4768 6518 4780
rect 6549 4777 6561 4780
rect 6595 4777 6607 4811
rect 6549 4771 6607 4777
rect 7374 4740 7380 4752
rect 5675 4712 7380 4740
rect 5675 4709 5687 4712
rect 5629 4703 5687 4709
rect 7374 4700 7380 4712
rect 7432 4700 7438 4752
rect 4264 4644 6316 4672
rect 4264 4616 4292 4644
rect 3142 4564 3148 4616
rect 3200 4564 3206 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4154 4604 4160 4616
rect 4019 4576 4160 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5534 4604 5540 4616
rect 5040 4576 5540 4604
rect 5040 4564 5046 4576
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6086 4604 6092 4616
rect 5767 4576 6092 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6178 4536 6184 4548
rect 6052 4508 6184 4536
rect 6052 4496 6058 4508
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 6288 4536 6316 4644
rect 6397 4539 6455 4545
rect 6397 4536 6409 4539
rect 6288 4508 6409 4536
rect 6397 4505 6409 4508
rect 6443 4536 6455 4539
rect 6914 4536 6920 4548
rect 6443 4508 6920 4536
rect 6443 4505 6455 4508
rect 6397 4499 6455 4505
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 2958 4428 2964 4480
rect 3016 4468 3022 4480
rect 3053 4471 3111 4477
rect 3053 4468 3065 4471
rect 3016 4440 3065 4468
rect 3016 4428 3022 4440
rect 3053 4437 3065 4440
rect 3099 4437 3111 4471
rect 3053 4431 3111 4437
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4522 4468 4528 4480
rect 4203 4440 4528 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 5500 4236 6561 4264
rect 5500 4224 5506 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4128 2838 4140
rect 3142 4128 3148 4140
rect 2832 4100 3148 4128
rect 2832 4088 2838 4100
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3320 4131 3378 4137
rect 3320 4097 3332 4131
rect 3366 4128 3378 4131
rect 3366 4100 4936 4128
rect 3366 4097 3378 4100
rect 3320 4091 3378 4097
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 3053 4063 3111 4069
rect 3053 4060 3065 4063
rect 2547 4032 3065 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 3053 4029 3065 4032
rect 3099 4029 3111 4063
rect 3053 4023 3111 4029
rect 4908 4001 4936 4100
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 5684 4100 6929 4128
rect 5684 4088 5690 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 5166 4020 5172 4072
rect 5224 4060 5230 4072
rect 5353 4063 5411 4069
rect 5353 4060 5365 4063
rect 5224 4032 5365 4060
rect 5224 4020 5230 4032
rect 5353 4029 5365 4032
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4029 5503 4063
rect 5445 4023 5503 4029
rect 4893 3995 4951 4001
rect 4893 3961 4905 3995
rect 4939 3961 4951 3995
rect 5460 3992 5488 4023
rect 6822 4020 6828 4072
rect 6880 4020 6886 4072
rect 6932 4060 6960 4091
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7576 4060 7604 4091
rect 6932 4032 7604 4060
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 5460 3964 7389 3992
rect 4893 3955 4951 3961
rect 7377 3961 7389 3964
rect 7423 3961 7435 3995
rect 7377 3955 7435 3961
rect 4430 3884 4436 3936
rect 4488 3884 4494 3936
rect 6730 3884 6736 3936
rect 6788 3884 6794 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 4212 3692 4353 3720
rect 4212 3680 4218 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 4341 3683 4399 3689
rect 4246 3612 4252 3664
rect 4304 3612 4310 3664
rect 7098 3652 7104 3664
rect 6472 3624 7104 3652
rect 6472 3596 6500 3624
rect 7098 3612 7104 3624
rect 7156 3652 7162 3664
rect 7285 3655 7343 3661
rect 7285 3652 7297 3655
rect 7156 3624 7297 3652
rect 7156 3612 7162 3624
rect 7285 3621 7297 3624
rect 7331 3621 7343 3655
rect 7285 3615 7343 3621
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4488 3556 4997 3584
rect 4488 3544 4494 3556
rect 4985 3553 4997 3556
rect 5031 3584 5043 3587
rect 5258 3584 5264 3596
rect 5031 3556 5264 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5442 3544 5448 3596
rect 5500 3544 5506 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5626 3584 5632 3596
rect 5583 3556 5632 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6178 3544 6184 3596
rect 6236 3584 6242 3596
rect 6340 3587 6398 3593
rect 6340 3584 6352 3587
rect 6236 3556 6352 3584
rect 6236 3544 6242 3556
rect 6340 3553 6352 3556
rect 6386 3553 6398 3587
rect 6340 3547 6398 3553
rect 6454 3544 6460 3596
rect 6512 3544 6518 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6730 3584 6736 3596
rect 6595 3556 6736 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 6972 3556 7788 3584
rect 6972 3544 6978 3556
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 2774 3516 2780 3528
rect 2455 3488 2780 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 2958 3476 2964 3528
rect 3016 3476 3022 3528
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4246 3516 4252 3528
rect 4203 3488 4252 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2096 3352 2237 3380
rect 2096 3340 2102 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 3160 3380 3188 3479
rect 4246 3476 4252 3488
rect 4304 3516 4310 3528
rect 4522 3516 4528 3528
rect 4304 3488 4528 3516
rect 4304 3476 4310 3488
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5460 3516 5488 3544
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 5460 3488 5534 3516
rect 3234 3408 3240 3460
rect 3292 3408 3298 3460
rect 5506 3448 5534 3488
rect 6196 3488 6592 3516
rect 6196 3448 6224 3488
rect 5506 3420 6224 3448
rect 6564 3448 6592 3488
rect 6886 3488 7665 3516
rect 6886 3448 6914 3488
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 6564 3420 6914 3448
rect 7561 3451 7619 3457
rect 7561 3417 7573 3451
rect 7607 3448 7619 3451
rect 7760 3448 7788 3556
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 7607 3420 7788 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 5166 3380 5172 3392
rect 3160 3352 5172 3380
rect 2225 3343 2283 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 6178 3340 6184 3392
rect 6236 3340 6242 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 6328 3352 7481 3380
rect 6328 3340 6334 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 7837 3383 7895 3389
rect 7837 3349 7849 3383
rect 7883 3380 7895 3383
rect 9122 3380 9128 3392
rect 7883 3352 9128 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6730 3176 6736 3188
rect 5951 3148 6736 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6822 3136 6828 3188
rect 6880 3136 6886 3188
rect 2038 3068 2044 3120
rect 2096 3068 2102 3120
rect 2774 3068 2780 3120
rect 2832 3068 2838 3120
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 5166 3068 5172 3120
rect 5224 3108 5230 3120
rect 5224 3080 9904 3108
rect 5224 3068 5230 3080
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5500 3012 5825 3040
rect 5500 3000 5506 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6932 2972 6960 3003
rect 7098 3000 7104 3052
rect 7156 3000 7162 3052
rect 9876 3049 9904 3080
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 6328 2944 6960 2972
rect 10137 2975 10195 2981
rect 6328 2932 6334 2944
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 11330 2972 11336 2984
rect 10183 2944 11336 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 1762 2864 1768 2916
rect 1820 2904 1826 2916
rect 1857 2907 1915 2913
rect 1857 2904 1869 2907
rect 1820 2876 1869 2904
rect 1820 2864 1826 2876
rect 1857 2873 1869 2876
rect 1903 2873 1915 2907
rect 1857 2867 1915 2873
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2836 6607 2839
rect 6638 2836 6644 2848
rect 6595 2808 6644 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 10226 2836 10232 2848
rect 9447 2808 10232 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 7926 2524 7932 2576
rect 7984 2564 7990 2576
rect 10045 2567 10103 2573
rect 10045 2564 10057 2567
rect 7984 2536 10057 2564
rect 7984 2524 7990 2536
rect 10045 2533 10057 2536
rect 10091 2533 10103 2567
rect 10045 2527 10103 2533
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2498 2428 2504 2440
rect 2087 2400 2504 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4304 2400 4721 2428
rect 4304 2388 4310 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6178 2428 6184 2440
rect 5951 2400 6184 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 624 2332 1777 2360
rect 624 2320 630 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 3016 2332 3065 2360
rect 3016 2320 3022 2332
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4433 2363 4491 2369
rect 4433 2360 4445 2363
rect 4212 2332 4445 2360
rect 4212 2320 4218 2332
rect 4433 2329 4445 2332
rect 4479 2329 4491 2363
rect 4433 2323 4491 2329
rect 5534 2320 5540 2372
rect 5592 2360 5598 2372
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 5592 2332 5641 2360
rect 5592 2320 5598 2332
rect 5629 2329 5641 2332
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 6917 2363 6975 2369
rect 6917 2360 6929 2363
rect 6604 2332 6929 2360
rect 6604 2320 6610 2332
rect 6917 2329 6929 2332
rect 6963 2329 6975 2363
rect 6917 2323 6975 2329
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7800 2332 8125 2360
rect 7800 2320 7806 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8996 2332 9413 2360
rect 8996 2320 9002 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 10226 2320 10232 2372
rect 10284 2320 10290 2372
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
<< via1 >>
rect 2169 15750 2221 15802
rect 2233 15750 2285 15802
rect 2297 15750 2349 15802
rect 2361 15750 2413 15802
rect 2425 15750 2477 15802
rect 4607 15750 4659 15802
rect 4671 15750 4723 15802
rect 4735 15750 4787 15802
rect 4799 15750 4851 15802
rect 4863 15750 4915 15802
rect 7045 15750 7097 15802
rect 7109 15750 7161 15802
rect 7173 15750 7225 15802
rect 7237 15750 7289 15802
rect 7301 15750 7353 15802
rect 9483 15750 9535 15802
rect 9547 15750 9599 15802
rect 9611 15750 9663 15802
rect 9675 15750 9727 15802
rect 9739 15750 9791 15802
rect 8944 15648 8996 15700
rect 8944 15444 8996 15496
rect 10324 15444 10376 15496
rect 11060 15444 11112 15496
rect 9128 15419 9180 15428
rect 9128 15385 9137 15419
rect 9137 15385 9171 15419
rect 9171 15385 9180 15419
rect 9128 15376 9180 15385
rect 9864 15376 9916 15428
rect 3388 15206 3440 15258
rect 3452 15206 3504 15258
rect 3516 15206 3568 15258
rect 3580 15206 3632 15258
rect 3644 15206 3696 15258
rect 5826 15206 5878 15258
rect 5890 15206 5942 15258
rect 5954 15206 6006 15258
rect 6018 15206 6070 15258
rect 6082 15206 6134 15258
rect 8264 15206 8316 15258
rect 8328 15206 8380 15258
rect 8392 15206 8444 15258
rect 8456 15206 8508 15258
rect 8520 15206 8572 15258
rect 10702 15206 10754 15258
rect 10766 15206 10818 15258
rect 10830 15206 10882 15258
rect 10894 15206 10946 15258
rect 10958 15206 11010 15258
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 2169 14662 2221 14714
rect 2233 14662 2285 14714
rect 2297 14662 2349 14714
rect 2361 14662 2413 14714
rect 2425 14662 2477 14714
rect 4607 14662 4659 14714
rect 4671 14662 4723 14714
rect 4735 14662 4787 14714
rect 4799 14662 4851 14714
rect 4863 14662 4915 14714
rect 7045 14662 7097 14714
rect 7109 14662 7161 14714
rect 7173 14662 7225 14714
rect 7237 14662 7289 14714
rect 7301 14662 7353 14714
rect 9483 14662 9535 14714
rect 9547 14662 9599 14714
rect 9611 14662 9663 14714
rect 9675 14662 9727 14714
rect 9739 14662 9791 14714
rect 3388 14118 3440 14170
rect 3452 14118 3504 14170
rect 3516 14118 3568 14170
rect 3580 14118 3632 14170
rect 3644 14118 3696 14170
rect 5826 14118 5878 14170
rect 5890 14118 5942 14170
rect 5954 14118 6006 14170
rect 6018 14118 6070 14170
rect 6082 14118 6134 14170
rect 8264 14118 8316 14170
rect 8328 14118 8380 14170
rect 8392 14118 8444 14170
rect 8456 14118 8508 14170
rect 8520 14118 8572 14170
rect 10702 14118 10754 14170
rect 10766 14118 10818 14170
rect 10830 14118 10882 14170
rect 10894 14118 10946 14170
rect 10958 14118 11010 14170
rect 2169 13574 2221 13626
rect 2233 13574 2285 13626
rect 2297 13574 2349 13626
rect 2361 13574 2413 13626
rect 2425 13574 2477 13626
rect 4607 13574 4659 13626
rect 4671 13574 4723 13626
rect 4735 13574 4787 13626
rect 4799 13574 4851 13626
rect 4863 13574 4915 13626
rect 7045 13574 7097 13626
rect 7109 13574 7161 13626
rect 7173 13574 7225 13626
rect 7237 13574 7289 13626
rect 7301 13574 7353 13626
rect 9483 13574 9535 13626
rect 9547 13574 9599 13626
rect 9611 13574 9663 13626
rect 9675 13574 9727 13626
rect 9739 13574 9791 13626
rect 3388 13030 3440 13082
rect 3452 13030 3504 13082
rect 3516 13030 3568 13082
rect 3580 13030 3632 13082
rect 3644 13030 3696 13082
rect 5826 13030 5878 13082
rect 5890 13030 5942 13082
rect 5954 13030 6006 13082
rect 6018 13030 6070 13082
rect 6082 13030 6134 13082
rect 8264 13030 8316 13082
rect 8328 13030 8380 13082
rect 8392 13030 8444 13082
rect 8456 13030 8508 13082
rect 8520 13030 8572 13082
rect 10702 13030 10754 13082
rect 10766 13030 10818 13082
rect 10830 13030 10882 13082
rect 10894 13030 10946 13082
rect 10958 13030 11010 13082
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 7472 12656 7524 12708
rect 2169 12486 2221 12538
rect 2233 12486 2285 12538
rect 2297 12486 2349 12538
rect 2361 12486 2413 12538
rect 2425 12486 2477 12538
rect 4607 12486 4659 12538
rect 4671 12486 4723 12538
rect 4735 12486 4787 12538
rect 4799 12486 4851 12538
rect 4863 12486 4915 12538
rect 7045 12486 7097 12538
rect 7109 12486 7161 12538
rect 7173 12486 7225 12538
rect 7237 12486 7289 12538
rect 7301 12486 7353 12538
rect 9483 12486 9535 12538
rect 9547 12486 9599 12538
rect 9611 12486 9663 12538
rect 9675 12486 9727 12538
rect 9739 12486 9791 12538
rect 3388 11942 3440 11994
rect 3452 11942 3504 11994
rect 3516 11942 3568 11994
rect 3580 11942 3632 11994
rect 3644 11942 3696 11994
rect 5826 11942 5878 11994
rect 5890 11942 5942 11994
rect 5954 11942 6006 11994
rect 6018 11942 6070 11994
rect 6082 11942 6134 11994
rect 8264 11942 8316 11994
rect 8328 11942 8380 11994
rect 8392 11942 8444 11994
rect 8456 11942 8508 11994
rect 8520 11942 8572 11994
rect 10702 11942 10754 11994
rect 10766 11942 10818 11994
rect 10830 11942 10882 11994
rect 10894 11942 10946 11994
rect 10958 11942 11010 11994
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 7748 11636 7800 11688
rect 5632 11500 5684 11552
rect 6828 11500 6880 11552
rect 2169 11398 2221 11450
rect 2233 11398 2285 11450
rect 2297 11398 2349 11450
rect 2361 11398 2413 11450
rect 2425 11398 2477 11450
rect 4607 11398 4659 11450
rect 4671 11398 4723 11450
rect 4735 11398 4787 11450
rect 4799 11398 4851 11450
rect 4863 11398 4915 11450
rect 7045 11398 7097 11450
rect 7109 11398 7161 11450
rect 7173 11398 7225 11450
rect 7237 11398 7289 11450
rect 7301 11398 7353 11450
rect 9483 11398 9535 11450
rect 9547 11398 9599 11450
rect 9611 11398 9663 11450
rect 9675 11398 9727 11450
rect 9739 11398 9791 11450
rect 6552 11296 6604 11348
rect 3792 11092 3844 11144
rect 5540 11024 5592 11076
rect 3388 10854 3440 10906
rect 3452 10854 3504 10906
rect 3516 10854 3568 10906
rect 3580 10854 3632 10906
rect 3644 10854 3696 10906
rect 5826 10854 5878 10906
rect 5890 10854 5942 10906
rect 5954 10854 6006 10906
rect 6018 10854 6070 10906
rect 6082 10854 6134 10906
rect 8264 10854 8316 10906
rect 8328 10854 8380 10906
rect 8392 10854 8444 10906
rect 8456 10854 8508 10906
rect 8520 10854 8572 10906
rect 10702 10854 10754 10906
rect 10766 10854 10818 10906
rect 10830 10854 10882 10906
rect 10894 10854 10946 10906
rect 10958 10854 11010 10906
rect 6460 10752 6512 10804
rect 5540 10684 5592 10736
rect 3792 10616 3844 10668
rect 6736 10616 6788 10668
rect 6828 10616 6880 10668
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 9128 10616 9180 10668
rect 6276 10548 6328 10600
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 2169 10310 2221 10362
rect 2233 10310 2285 10362
rect 2297 10310 2349 10362
rect 2361 10310 2413 10362
rect 2425 10310 2477 10362
rect 4607 10310 4659 10362
rect 4671 10310 4723 10362
rect 4735 10310 4787 10362
rect 4799 10310 4851 10362
rect 4863 10310 4915 10362
rect 7045 10310 7097 10362
rect 7109 10310 7161 10362
rect 7173 10310 7225 10362
rect 7237 10310 7289 10362
rect 7301 10310 7353 10362
rect 9483 10310 9535 10362
rect 9547 10310 9599 10362
rect 9611 10310 9663 10362
rect 9675 10310 9727 10362
rect 9739 10310 9791 10362
rect 6644 10208 6696 10260
rect 6736 10208 6788 10260
rect 6368 10004 6420 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 4528 9460 4580 9512
rect 5724 9435 5776 9444
rect 5724 9401 5733 9435
rect 5733 9401 5767 9435
rect 5767 9401 5776 9435
rect 5724 9392 5776 9401
rect 6184 9460 6236 9512
rect 6368 9392 6420 9444
rect 5356 9324 5408 9376
rect 6092 9324 6144 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 6276 9120 6328 9172
rect 4988 9052 5040 9104
rect 5724 9052 5776 9104
rect 7656 9052 7708 9104
rect 6552 8984 6604 9036
rect 3792 8916 3844 8968
rect 5080 8848 5132 8900
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 6368 8848 6420 8900
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 3056 8780 3108 8832
rect 6552 8780 6604 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 5080 8576 5132 8628
rect 6184 8576 6236 8628
rect 5724 8508 5776 8560
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 6920 8508 6972 8560
rect 6828 8440 6880 8492
rect 7380 8440 7432 8492
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 6644 8372 6696 8424
rect 9864 8372 9916 8424
rect 4528 8236 4580 8288
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 7380 8032 7432 8084
rect 6276 7964 6328 8016
rect 6460 7964 6512 8016
rect 3056 7828 3108 7880
rect 3792 7828 3844 7880
rect 6000 7896 6052 7948
rect 6460 7828 6512 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 3884 7692 3936 7744
rect 4344 7692 4396 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 6368 7488 6420 7540
rect 5172 7463 5224 7472
rect 5172 7429 5181 7463
rect 5181 7429 5215 7463
rect 5215 7429 5224 7463
rect 5172 7420 5224 7429
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 5724 7352 5776 7404
rect 6644 7352 6696 7404
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 4252 7148 4304 7200
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 5264 6944 5316 6996
rect 3884 6808 3936 6860
rect 4252 6783 4304 6792
rect 4252 6749 4286 6783
rect 4286 6749 4304 6783
rect 4252 6740 4304 6749
rect 5632 6740 5684 6792
rect 6644 6740 6696 6792
rect 6552 6604 6604 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 6276 6264 6328 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 6920 6264 6972 6316
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 5080 5856 5132 5908
rect 6368 5856 6420 5908
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 7748 5856 7800 5908
rect 6736 5788 6788 5840
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4528 5652 4580 5704
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 8024 5720 8076 5772
rect 7196 5584 7248 5636
rect 7288 5627 7340 5636
rect 7288 5593 7297 5627
rect 7297 5593 7331 5627
rect 7331 5593 7340 5627
rect 7288 5584 7340 5593
rect 10232 5627 10284 5636
rect 10232 5593 10241 5627
rect 10241 5593 10275 5627
rect 10275 5593 10284 5627
rect 10232 5584 10284 5593
rect 7840 5516 7892 5568
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 4988 5312 5040 5364
rect 6828 5312 6880 5364
rect 7196 5312 7248 5364
rect 3148 5176 3200 5228
rect 3976 5244 4028 5296
rect 8116 5244 8168 5296
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 6092 5176 6144 5228
rect 6368 5176 6420 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 6828 5176 6880 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 6552 5108 6604 5160
rect 7288 5108 7340 5160
rect 6000 5040 6052 5092
rect 6276 5040 6328 5092
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6920 4972 6972 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 2504 4700 2556 4752
rect 6460 4768 6512 4820
rect 7380 4700 7432 4752
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 4160 4564 4212 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4988 4564 5040 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6092 4564 6144 4616
rect 6000 4496 6052 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 6920 4496 6972 4548
rect 2964 4428 3016 4480
rect 4528 4428 4580 4480
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 5448 4224 5500 4276
rect 2780 4088 2832 4140
rect 3148 4088 3200 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5632 4088 5684 4140
rect 5172 4020 5224 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 4160 3680 4212 3732
rect 4252 3655 4304 3664
rect 4252 3621 4261 3655
rect 4261 3621 4295 3655
rect 4295 3621 4304 3655
rect 4252 3612 4304 3621
rect 7104 3612 7156 3664
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5264 3544 5316 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5632 3544 5684 3596
rect 6184 3544 6236 3596
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 6736 3544 6788 3596
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 6920 3544 6972 3596
rect 2780 3476 2832 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 2044 3340 2096 3392
rect 4252 3476 4304 3528
rect 4528 3476 4580 3528
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 6276 3340 6328 3392
rect 9128 3340 9180 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 6736 3179 6788 3188
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 5172 3068 5224 3120
rect 5448 3000 5500 3052
rect 6276 2932 6328 2984
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 11336 2932 11388 2984
rect 1768 2864 1820 2916
rect 6644 2796 6696 2848
rect 10232 2796 10284 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 7932 2524 7984 2576
rect 2504 2388 2556 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4252 2388 4304 2440
rect 6184 2388 6236 2440
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 572 2320 624 2372
rect 2964 2320 3016 2372
rect 4160 2320 4212 2372
rect 5540 2320 5592 2372
rect 6552 2320 6604 2372
rect 7748 2320 7800 2372
rect 8944 2320 8996 2372
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
<< metal2 >>
rect 2962 17354 3018 18000
rect 2792 17326 3018 17354
rect 2169 15804 2477 15813
rect 2169 15802 2175 15804
rect 2231 15802 2255 15804
rect 2311 15802 2335 15804
rect 2391 15802 2415 15804
rect 2471 15802 2477 15804
rect 2231 15750 2233 15802
rect 2413 15750 2415 15802
rect 2169 15748 2175 15750
rect 2231 15748 2255 15750
rect 2311 15748 2335 15750
rect 2391 15748 2415 15750
rect 2471 15748 2477 15750
rect 2169 15739 2477 15748
rect 2169 14716 2477 14725
rect 2169 14714 2175 14716
rect 2231 14714 2255 14716
rect 2311 14714 2335 14716
rect 2391 14714 2415 14716
rect 2471 14714 2477 14716
rect 2231 14662 2233 14714
rect 2413 14662 2415 14714
rect 2169 14660 2175 14662
rect 2231 14660 2255 14662
rect 2311 14660 2335 14662
rect 2391 14660 2415 14662
rect 2471 14660 2477 14662
rect 2169 14651 2477 14660
rect 2169 13628 2477 13637
rect 2169 13626 2175 13628
rect 2231 13626 2255 13628
rect 2311 13626 2335 13628
rect 2391 13626 2415 13628
rect 2471 13626 2477 13628
rect 2231 13574 2233 13626
rect 2413 13574 2415 13626
rect 2169 13572 2175 13574
rect 2231 13572 2255 13574
rect 2311 13572 2335 13574
rect 2391 13572 2415 13574
rect 2471 13572 2477 13574
rect 2169 13563 2477 13572
rect 2169 12540 2477 12549
rect 2169 12538 2175 12540
rect 2231 12538 2255 12540
rect 2311 12538 2335 12540
rect 2391 12538 2415 12540
rect 2471 12538 2477 12540
rect 2231 12486 2233 12538
rect 2413 12486 2415 12538
rect 2169 12484 2175 12486
rect 2231 12484 2255 12486
rect 2311 12484 2335 12486
rect 2391 12484 2415 12486
rect 2471 12484 2477 12486
rect 2169 12475 2477 12484
rect 2169 11452 2477 11461
rect 2169 11450 2175 11452
rect 2231 11450 2255 11452
rect 2311 11450 2335 11452
rect 2391 11450 2415 11452
rect 2471 11450 2477 11452
rect 2231 11398 2233 11450
rect 2413 11398 2415 11450
rect 2169 11396 2175 11398
rect 2231 11396 2255 11398
rect 2311 11396 2335 11398
rect 2391 11396 2415 11398
rect 2471 11396 2477 11398
rect 2169 11387 2477 11396
rect 2169 10364 2477 10373
rect 2169 10362 2175 10364
rect 2231 10362 2255 10364
rect 2311 10362 2335 10364
rect 2391 10362 2415 10364
rect 2471 10362 2477 10364
rect 2231 10310 2233 10362
rect 2413 10310 2415 10362
rect 2169 10308 2175 10310
rect 2231 10308 2255 10310
rect 2311 10308 2335 10310
rect 2391 10308 2415 10310
rect 2471 10308 2477 10310
rect 2169 10299 2477 10308
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2792 8090 2820 17326
rect 2962 17200 3018 17326
rect 8942 17200 8998 18000
rect 4607 15804 4915 15813
rect 4607 15802 4613 15804
rect 4669 15802 4693 15804
rect 4749 15802 4773 15804
rect 4829 15802 4853 15804
rect 4909 15802 4915 15804
rect 4669 15750 4671 15802
rect 4851 15750 4853 15802
rect 4607 15748 4613 15750
rect 4669 15748 4693 15750
rect 4749 15748 4773 15750
rect 4829 15748 4853 15750
rect 4909 15748 4915 15750
rect 4607 15739 4915 15748
rect 7045 15804 7353 15813
rect 7045 15802 7051 15804
rect 7107 15802 7131 15804
rect 7187 15802 7211 15804
rect 7267 15802 7291 15804
rect 7347 15802 7353 15804
rect 7107 15750 7109 15802
rect 7289 15750 7291 15802
rect 7045 15748 7051 15750
rect 7107 15748 7131 15750
rect 7187 15748 7211 15750
rect 7267 15748 7291 15750
rect 7347 15748 7353 15750
rect 7045 15739 7353 15748
rect 8956 15706 8984 17200
rect 11058 16008 11114 16017
rect 11058 15943 11114 15952
rect 9483 15804 9791 15813
rect 9483 15802 9489 15804
rect 9545 15802 9569 15804
rect 9625 15802 9649 15804
rect 9705 15802 9729 15804
rect 9785 15802 9791 15804
rect 9545 15750 9547 15802
rect 9727 15750 9729 15802
rect 9483 15748 9489 15750
rect 9545 15748 9569 15750
rect 9625 15748 9649 15750
rect 9705 15748 9729 15750
rect 9785 15748 9791 15750
rect 9483 15739 9791 15748
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8956 15502 8984 15642
rect 11072 15502 11100 15943
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 3388 15260 3696 15269
rect 3388 15258 3394 15260
rect 3450 15258 3474 15260
rect 3530 15258 3554 15260
rect 3610 15258 3634 15260
rect 3690 15258 3696 15260
rect 3450 15206 3452 15258
rect 3632 15206 3634 15258
rect 3388 15204 3394 15206
rect 3450 15204 3474 15206
rect 3530 15204 3554 15206
rect 3610 15204 3634 15206
rect 3690 15204 3696 15206
rect 3388 15195 3696 15204
rect 5826 15260 6134 15269
rect 5826 15258 5832 15260
rect 5888 15258 5912 15260
rect 5968 15258 5992 15260
rect 6048 15258 6072 15260
rect 6128 15258 6134 15260
rect 5888 15206 5890 15258
rect 6070 15206 6072 15258
rect 5826 15204 5832 15206
rect 5888 15204 5912 15206
rect 5968 15204 5992 15206
rect 6048 15204 6072 15206
rect 6128 15204 6134 15206
rect 5826 15195 6134 15204
rect 8264 15260 8572 15269
rect 8264 15258 8270 15260
rect 8326 15258 8350 15260
rect 8406 15258 8430 15260
rect 8486 15258 8510 15260
rect 8566 15258 8572 15260
rect 8326 15206 8328 15258
rect 8508 15206 8510 15258
rect 8264 15204 8270 15206
rect 8326 15204 8350 15206
rect 8406 15204 8430 15206
rect 8486 15204 8510 15206
rect 8566 15204 8572 15206
rect 8264 15195 8572 15204
rect 4607 14716 4915 14725
rect 4607 14714 4613 14716
rect 4669 14714 4693 14716
rect 4749 14714 4773 14716
rect 4829 14714 4853 14716
rect 4909 14714 4915 14716
rect 4669 14662 4671 14714
rect 4851 14662 4853 14714
rect 4607 14660 4613 14662
rect 4669 14660 4693 14662
rect 4749 14660 4773 14662
rect 4829 14660 4853 14662
rect 4909 14660 4915 14662
rect 4607 14651 4915 14660
rect 7045 14716 7353 14725
rect 7045 14714 7051 14716
rect 7107 14714 7131 14716
rect 7187 14714 7211 14716
rect 7267 14714 7291 14716
rect 7347 14714 7353 14716
rect 7107 14662 7109 14714
rect 7289 14662 7291 14714
rect 7045 14660 7051 14662
rect 7107 14660 7131 14662
rect 7187 14660 7211 14662
rect 7267 14660 7291 14662
rect 7347 14660 7353 14662
rect 7045 14651 7353 14660
rect 3388 14172 3696 14181
rect 3388 14170 3394 14172
rect 3450 14170 3474 14172
rect 3530 14170 3554 14172
rect 3610 14170 3634 14172
rect 3690 14170 3696 14172
rect 3450 14118 3452 14170
rect 3632 14118 3634 14170
rect 3388 14116 3394 14118
rect 3450 14116 3474 14118
rect 3530 14116 3554 14118
rect 3610 14116 3634 14118
rect 3690 14116 3696 14118
rect 3388 14107 3696 14116
rect 5826 14172 6134 14181
rect 5826 14170 5832 14172
rect 5888 14170 5912 14172
rect 5968 14170 5992 14172
rect 6048 14170 6072 14172
rect 6128 14170 6134 14172
rect 5888 14118 5890 14170
rect 6070 14118 6072 14170
rect 5826 14116 5832 14118
rect 5888 14116 5912 14118
rect 5968 14116 5992 14118
rect 6048 14116 6072 14118
rect 6128 14116 6134 14118
rect 5826 14107 6134 14116
rect 8264 14172 8572 14181
rect 8264 14170 8270 14172
rect 8326 14170 8350 14172
rect 8406 14170 8430 14172
rect 8486 14170 8510 14172
rect 8566 14170 8572 14172
rect 8326 14118 8328 14170
rect 8508 14118 8510 14170
rect 8264 14116 8270 14118
rect 8326 14116 8350 14118
rect 8406 14116 8430 14118
rect 8486 14116 8510 14118
rect 8566 14116 8572 14118
rect 8264 14107 8572 14116
rect 4607 13628 4915 13637
rect 4607 13626 4613 13628
rect 4669 13626 4693 13628
rect 4749 13626 4773 13628
rect 4829 13626 4853 13628
rect 4909 13626 4915 13628
rect 4669 13574 4671 13626
rect 4851 13574 4853 13626
rect 4607 13572 4613 13574
rect 4669 13572 4693 13574
rect 4749 13572 4773 13574
rect 4829 13572 4853 13574
rect 4909 13572 4915 13574
rect 4607 13563 4915 13572
rect 7045 13628 7353 13637
rect 7045 13626 7051 13628
rect 7107 13626 7131 13628
rect 7187 13626 7211 13628
rect 7267 13626 7291 13628
rect 7347 13626 7353 13628
rect 7107 13574 7109 13626
rect 7289 13574 7291 13626
rect 7045 13572 7051 13574
rect 7107 13572 7131 13574
rect 7187 13572 7211 13574
rect 7267 13572 7291 13574
rect 7347 13572 7353 13574
rect 7045 13563 7353 13572
rect 3388 13084 3696 13093
rect 3388 13082 3394 13084
rect 3450 13082 3474 13084
rect 3530 13082 3554 13084
rect 3610 13082 3634 13084
rect 3690 13082 3696 13084
rect 3450 13030 3452 13082
rect 3632 13030 3634 13082
rect 3388 13028 3394 13030
rect 3450 13028 3474 13030
rect 3530 13028 3554 13030
rect 3610 13028 3634 13030
rect 3690 13028 3696 13030
rect 3388 13019 3696 13028
rect 5826 13084 6134 13093
rect 5826 13082 5832 13084
rect 5888 13082 5912 13084
rect 5968 13082 5992 13084
rect 6048 13082 6072 13084
rect 6128 13082 6134 13084
rect 5888 13030 5890 13082
rect 6070 13030 6072 13082
rect 5826 13028 5832 13030
rect 5888 13028 5912 13030
rect 5968 13028 5992 13030
rect 6048 13028 6072 13030
rect 6128 13028 6134 13030
rect 5826 13019 6134 13028
rect 8264 13084 8572 13093
rect 8264 13082 8270 13084
rect 8326 13082 8350 13084
rect 8406 13082 8430 13084
rect 8486 13082 8510 13084
rect 8566 13082 8572 13084
rect 8326 13030 8328 13082
rect 8508 13030 8510 13082
rect 8264 13028 8270 13030
rect 8326 13028 8350 13030
rect 8406 13028 8430 13030
rect 8486 13028 8510 13030
rect 8566 13028 8572 13030
rect 8264 13019 8572 13028
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 4607 12540 4915 12549
rect 4607 12538 4613 12540
rect 4669 12538 4693 12540
rect 4749 12538 4773 12540
rect 4829 12538 4853 12540
rect 4909 12538 4915 12540
rect 4669 12486 4671 12538
rect 4851 12486 4853 12538
rect 4607 12484 4613 12486
rect 4669 12484 4693 12486
rect 4749 12484 4773 12486
rect 4829 12484 4853 12486
rect 4909 12484 4915 12486
rect 4607 12475 4915 12484
rect 7045 12540 7353 12549
rect 7045 12538 7051 12540
rect 7107 12538 7131 12540
rect 7187 12538 7211 12540
rect 7267 12538 7291 12540
rect 7347 12538 7353 12540
rect 7107 12486 7109 12538
rect 7289 12486 7291 12538
rect 7045 12484 7051 12486
rect 7107 12484 7131 12486
rect 7187 12484 7211 12486
rect 7267 12484 7291 12486
rect 7347 12484 7353 12486
rect 7045 12475 7353 12484
rect 3388 11996 3696 12005
rect 3388 11994 3394 11996
rect 3450 11994 3474 11996
rect 3530 11994 3554 11996
rect 3610 11994 3634 11996
rect 3690 11994 3696 11996
rect 3450 11942 3452 11994
rect 3632 11942 3634 11994
rect 3388 11940 3394 11942
rect 3450 11940 3474 11942
rect 3530 11940 3554 11942
rect 3610 11940 3634 11942
rect 3690 11940 3696 11942
rect 3388 11931 3696 11940
rect 5826 11996 6134 12005
rect 5826 11994 5832 11996
rect 5888 11994 5912 11996
rect 5968 11994 5992 11996
rect 6048 11994 6072 11996
rect 6128 11994 6134 11996
rect 5888 11942 5890 11994
rect 6070 11942 6072 11994
rect 5826 11940 5832 11942
rect 5888 11940 5912 11942
rect 5968 11940 5992 11942
rect 6048 11940 6072 11942
rect 6128 11940 6134 11942
rect 5826 11931 6134 11940
rect 7484 11762 7512 12650
rect 8264 11996 8572 12005
rect 8264 11994 8270 11996
rect 8326 11994 8350 11996
rect 8406 11994 8430 11996
rect 8486 11994 8510 11996
rect 8566 11994 8572 11996
rect 8326 11942 8328 11994
rect 8508 11942 8510 11994
rect 8264 11940 8270 11942
rect 8326 11940 8350 11942
rect 8406 11940 8430 11942
rect 8486 11940 8510 11942
rect 8566 11940 8572 11942
rect 8264 11931 8572 11940
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 11150 3832 11630
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 4607 11452 4915 11461
rect 4607 11450 4613 11452
rect 4669 11450 4693 11452
rect 4749 11450 4773 11452
rect 4829 11450 4853 11452
rect 4909 11450 4915 11452
rect 4669 11398 4671 11450
rect 4851 11398 4853 11450
rect 4607 11396 4613 11398
rect 4669 11396 4693 11398
rect 4749 11396 4773 11398
rect 4829 11396 4853 11398
rect 4909 11396 4915 11398
rect 4607 11387 4915 11396
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3388 10908 3696 10917
rect 3388 10906 3394 10908
rect 3450 10906 3474 10908
rect 3530 10906 3554 10908
rect 3610 10906 3634 10908
rect 3690 10906 3696 10908
rect 3450 10854 3452 10906
rect 3632 10854 3634 10906
rect 3388 10852 3394 10854
rect 3450 10852 3474 10854
rect 3530 10852 3554 10854
rect 3610 10852 3634 10854
rect 3690 10852 3696 10854
rect 3388 10843 3696 10852
rect 3804 10674 3832 11086
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10742 5580 11018
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3804 8974 3832 10610
rect 4607 10364 4915 10373
rect 4607 10362 4613 10364
rect 4669 10362 4693 10364
rect 4749 10362 4773 10364
rect 4829 10362 4853 10364
rect 4909 10362 4915 10364
rect 4669 10310 4671 10362
rect 4851 10310 4853 10362
rect 4607 10308 4613 10310
rect 4669 10308 4693 10310
rect 4749 10308 4773 10310
rect 4829 10308 4853 10310
rect 4909 10308 4915 10310
rect 4607 10299 4915 10308
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8498 3096 8774
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3804 7886 3832 8910
rect 4540 8294 4568 9454
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3068 7546 3096 7822
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 3896 6866 3924 7686
rect 4356 7410 4384 7686
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 4264 6798 4292 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3988 5302 4016 5646
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 3126 2084 3334
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 584 800 612 2314
rect 1780 800 1808 2858
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2516 2446 2544 4694
rect 3160 4622 3188 5170
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 3534 2820 4082
rect 2976 3534 3004 4422
rect 3160 4146 3188 4558
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 4172 3738 4200 4558
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3670 4292 4558
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 2792 3126 2820 3470
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3252 2446 3280 3402
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 4264 2446 4292 3470
rect 4356 3126 4384 7346
rect 4540 5710 4568 8230
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 4486 4568 5646
rect 5000 5370 5028 9046
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5092 8634 5120 8842
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5092 5914 5120 8570
rect 5368 8430 5396 9318
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 5000 4622 5028 5306
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4448 3602 4476 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4540 3534 4568 4422
rect 5184 4078 5212 7414
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5276 7002 5304 7278
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5460 4282 5488 7278
rect 5644 6798 5672 11494
rect 6564 11354 6592 11698
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5826 10908 6134 10917
rect 5826 10906 5832 10908
rect 5888 10906 5912 10908
rect 5968 10906 5992 10908
rect 6048 10906 6072 10908
rect 6128 10906 6134 10908
rect 5888 10854 5890 10906
rect 6070 10854 6072 10906
rect 5826 10852 5832 10854
rect 5888 10852 5912 10854
rect 5968 10852 5992 10854
rect 6048 10852 6072 10854
rect 6128 10852 6134 10854
rect 5826 10843 6134 10852
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5736 9110 5764 9386
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 6104 8974 6132 9318
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 6196 8634 6224 9454
rect 6288 9178 6316 10542
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9450 6408 9998
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6288 8974 6316 9114
rect 6472 8974 6500 10746
rect 6840 10674 6868 11494
rect 7045 11452 7353 11461
rect 7045 11450 7051 11452
rect 7107 11450 7131 11452
rect 7187 11450 7211 11452
rect 7267 11450 7291 11452
rect 7347 11450 7353 11452
rect 7107 11398 7109 11450
rect 7289 11398 7291 11450
rect 7045 11396 7051 11398
rect 7107 11396 7131 11398
rect 7187 11396 7211 11398
rect 7267 11396 7291 11398
rect 7347 11396 7353 11398
rect 7045 11387 7353 11396
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6828 10668 6880 10674
rect 7012 10668 7064 10674
rect 6828 10610 6880 10616
rect 6932 10628 7012 10656
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10266 6684 10542
rect 6748 10266 6776 10610
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9042 6592 9318
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5736 7410 5764 8502
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7954 6040 8230
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 6288 6322 6316 7958
rect 6380 7546 6408 8842
rect 6472 8022 6500 8910
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6564 7886 6592 8774
rect 6932 8566 6960 10628
rect 7012 10610 7064 10616
rect 7045 10364 7353 10373
rect 7045 10362 7051 10364
rect 7107 10362 7131 10364
rect 7187 10362 7211 10364
rect 7267 10362 7291 10364
rect 7347 10362 7353 10364
rect 7107 10310 7109 10362
rect 7289 10310 7291 10362
rect 7045 10308 7051 10310
rect 7107 10308 7131 10310
rect 7187 10308 7211 10310
rect 7267 10308 7291 10310
rect 7347 10308 7353 10310
rect 7045 10299 7353 10308
rect 7760 10062 7788 11630
rect 8264 10908 8572 10917
rect 8264 10906 8270 10908
rect 8326 10906 8350 10908
rect 8406 10906 8430 10908
rect 8486 10906 8510 10908
rect 8566 10906 8572 10908
rect 8326 10854 8328 10906
rect 8508 10854 8510 10906
rect 8264 10852 8270 10854
rect 8326 10852 8350 10854
rect 8406 10852 8430 10854
rect 8486 10852 8510 10854
rect 8566 10852 8572 10854
rect 8264 10843 8572 10852
rect 9140 10674 9168 15370
rect 9483 14716 9791 14725
rect 9483 14714 9489 14716
rect 9545 14714 9569 14716
rect 9625 14714 9649 14716
rect 9705 14714 9729 14716
rect 9785 14714 9791 14716
rect 9545 14662 9547 14714
rect 9727 14662 9729 14714
rect 9483 14660 9489 14662
rect 9545 14660 9569 14662
rect 9625 14660 9649 14662
rect 9705 14660 9729 14662
rect 9785 14660 9791 14662
rect 9483 14651 9791 14660
rect 9483 13628 9791 13637
rect 9483 13626 9489 13628
rect 9545 13626 9569 13628
rect 9625 13626 9649 13628
rect 9705 13626 9729 13628
rect 9785 13626 9791 13628
rect 9545 13574 9547 13626
rect 9727 13574 9729 13626
rect 9483 13572 9489 13574
rect 9545 13572 9569 13574
rect 9625 13572 9649 13574
rect 9705 13572 9729 13574
rect 9785 13572 9791 13574
rect 9483 13563 9791 13572
rect 9483 12540 9791 12549
rect 9483 12538 9489 12540
rect 9545 12538 9569 12540
rect 9625 12538 9649 12540
rect 9705 12538 9729 12540
rect 9785 12538 9791 12540
rect 9545 12486 9547 12538
rect 9727 12486 9729 12538
rect 9483 12484 9489 12486
rect 9545 12484 9569 12486
rect 9625 12484 9649 12486
rect 9705 12484 9729 12486
rect 9785 12484 9791 12486
rect 9483 12475 9791 12484
rect 9483 11452 9791 11461
rect 9483 11450 9489 11452
rect 9545 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9791 11452
rect 9545 11398 9547 11450
rect 9727 11398 9729 11450
rect 9483 11396 9489 11398
rect 9545 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9791 11398
rect 9483 11387 9791 11396
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9483 10364 9791 10373
rect 9483 10362 9489 10364
rect 9545 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9791 10364
rect 9545 10310 9547 10362
rect 9727 10310 9729 10362
rect 9483 10308 9489 10310
rect 9545 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9791 10310
rect 9483 10299 9791 10308
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7668 9110 7696 9998
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6472 7290 6500 7822
rect 6656 7410 6684 8366
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6472 7262 6592 7290
rect 6564 6662 6592 7262
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6012 5098 6040 5170
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5552 4154 5580 4558
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5460 4126 5580 4154
rect 5644 4146 5672 4966
rect 6012 4554 6040 5034
rect 6104 4622 6132 5170
rect 6288 5098 6316 6258
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6380 5234 6408 5850
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6472 4826 6500 5646
rect 6564 5166 6592 6598
rect 6656 5710 6684 6734
rect 6748 6322 6776 7822
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5846 6776 6054
rect 6840 5914 6868 8434
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7392 8090 7420 8434
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 5632 4140 5684 4146
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 5276 3602 5304 4082
rect 5460 3602 5488 4126
rect 5632 4082 5684 4088
rect 5644 3602 5672 4082
rect 6196 3602 6224 4490
rect 6656 4154 6684 5646
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6840 5234 6868 5306
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6564 4126 6684 4154
rect 6748 4154 6776 5170
rect 6932 5030 6960 6258
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 7760 5914 7788 9998
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 9876 8430 9904 15370
rect 10336 15162 10364 15438
rect 10702 15260 11010 15269
rect 10702 15258 10708 15260
rect 10764 15258 10788 15260
rect 10844 15258 10868 15260
rect 10924 15258 10948 15260
rect 11004 15258 11010 15260
rect 10764 15206 10766 15258
rect 10946 15206 10948 15258
rect 10702 15204 10708 15206
rect 10764 15204 10788 15206
rect 10844 15204 10868 15206
rect 10924 15204 10948 15206
rect 11004 15204 11010 15206
rect 10702 15195 11010 15204
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10702 14172 11010 14181
rect 10702 14170 10708 14172
rect 10764 14170 10788 14172
rect 10844 14170 10868 14172
rect 10924 14170 10948 14172
rect 11004 14170 11010 14172
rect 10764 14118 10766 14170
rect 10946 14118 10948 14170
rect 10702 14116 10708 14118
rect 10764 14116 10788 14118
rect 10844 14116 10868 14118
rect 10924 14116 10948 14118
rect 11004 14116 11010 14118
rect 10702 14107 11010 14116
rect 10702 13084 11010 13093
rect 10702 13082 10708 13084
rect 10764 13082 10788 13084
rect 10844 13082 10868 13084
rect 10924 13082 10948 13084
rect 11004 13082 11010 13084
rect 10764 13030 10766 13082
rect 10946 13030 10948 13082
rect 10702 13028 10708 13030
rect 10764 13028 10788 13030
rect 10844 13028 10868 13030
rect 10924 13028 10948 13030
rect 11004 13028 11010 13030
rect 10702 13019 11010 13028
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10244 12481 10272 12786
rect 10230 12472 10286 12481
rect 10230 12407 10286 12416
rect 10702 11996 11010 12005
rect 10702 11994 10708 11996
rect 10764 11994 10788 11996
rect 10844 11994 10868 11996
rect 10924 11994 10948 11996
rect 11004 11994 11010 11996
rect 10764 11942 10766 11994
rect 10946 11942 10948 11994
rect 10702 11940 10708 11942
rect 10764 11940 10788 11942
rect 10844 11940 10868 11942
rect 10924 11940 10948 11942
rect 11004 11940 11010 11942
rect 10702 11931 11010 11940
rect 10702 10908 11010 10917
rect 10702 10906 10708 10908
rect 10764 10906 10788 10908
rect 10844 10906 10868 10908
rect 10924 10906 10948 10908
rect 11004 10906 11010 10908
rect 10764 10854 10766 10906
rect 10946 10854 10948 10906
rect 10702 10852 10708 10854
rect 10764 10852 10788 10854
rect 10844 10852 10868 10854
rect 10924 10852 10948 10854
rect 11004 10852 11010 10854
rect 10702 10843 11010 10852
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 10230 8936 10286 8945
rect 10230 8871 10232 8880
rect 10284 8871 10286 8880
rect 10232 8842 10284 8848
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7208 5370 7236 5578
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7300 5166 7328 5578
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4554 6960 4966
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6748 4126 6868 4154
rect 7392 4146 7420 4694
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 6184 3596 6236 3602
rect 6460 3596 6512 3602
rect 6236 3556 6316 3584
rect 6184 3538 6236 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 3126 5212 3334
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5460 3058 5488 3538
rect 6288 3398 6316 3556
rect 6564 3584 6592 4126
rect 6840 4078 6868 4126
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3602 6776 3878
rect 6840 3602 6868 4014
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 6512 3556 6592 3584
rect 6736 3596 6788 3602
rect 6460 3538 6512 3544
rect 6736 3538 6788 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 6196 2446 6224 3334
rect 6288 2990 6316 3334
rect 6748 3194 6776 3538
rect 6840 3482 6868 3538
rect 6932 3482 6960 3538
rect 6840 3454 6960 3482
rect 6840 3194 6868 3454
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7116 3058 7144 3606
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2446 6684 2790
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7852 2446 7880 5510
rect 8036 5234 8064 5714
rect 10230 5672 10286 5681
rect 10230 5607 10232 5616
rect 10284 5607 10286 5616
rect 10232 5578 10284 5584
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8128 5302 8156 5510
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7944 2582 7972 5170
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 9140 2446 9168 3334
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 2976 800 3004 2314
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 4172 800 4200 2314
rect 5552 898 5580 2314
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 5368 870 5580 898
rect 5368 800 5396 870
rect 6564 800 6592 2314
rect 7760 800 7788 2314
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8956 800 8984 2314
rect 10152 800 10180 3470
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10244 2378 10272 2790
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10244 1873 10272 2314
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 10230 1864 10286 1873
rect 10230 1799 10286 1808
rect 11348 800 11376 2926
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
rect 11334 0 11390 800
<< via2 >>
rect 2175 15802 2231 15804
rect 2255 15802 2311 15804
rect 2335 15802 2391 15804
rect 2415 15802 2471 15804
rect 2175 15750 2221 15802
rect 2221 15750 2231 15802
rect 2255 15750 2285 15802
rect 2285 15750 2297 15802
rect 2297 15750 2311 15802
rect 2335 15750 2349 15802
rect 2349 15750 2361 15802
rect 2361 15750 2391 15802
rect 2415 15750 2425 15802
rect 2425 15750 2471 15802
rect 2175 15748 2231 15750
rect 2255 15748 2311 15750
rect 2335 15748 2391 15750
rect 2415 15748 2471 15750
rect 2175 14714 2231 14716
rect 2255 14714 2311 14716
rect 2335 14714 2391 14716
rect 2415 14714 2471 14716
rect 2175 14662 2221 14714
rect 2221 14662 2231 14714
rect 2255 14662 2285 14714
rect 2285 14662 2297 14714
rect 2297 14662 2311 14714
rect 2335 14662 2349 14714
rect 2349 14662 2361 14714
rect 2361 14662 2391 14714
rect 2415 14662 2425 14714
rect 2425 14662 2471 14714
rect 2175 14660 2231 14662
rect 2255 14660 2311 14662
rect 2335 14660 2391 14662
rect 2415 14660 2471 14662
rect 2175 13626 2231 13628
rect 2255 13626 2311 13628
rect 2335 13626 2391 13628
rect 2415 13626 2471 13628
rect 2175 13574 2221 13626
rect 2221 13574 2231 13626
rect 2255 13574 2285 13626
rect 2285 13574 2297 13626
rect 2297 13574 2311 13626
rect 2335 13574 2349 13626
rect 2349 13574 2361 13626
rect 2361 13574 2391 13626
rect 2415 13574 2425 13626
rect 2425 13574 2471 13626
rect 2175 13572 2231 13574
rect 2255 13572 2311 13574
rect 2335 13572 2391 13574
rect 2415 13572 2471 13574
rect 2175 12538 2231 12540
rect 2255 12538 2311 12540
rect 2335 12538 2391 12540
rect 2415 12538 2471 12540
rect 2175 12486 2221 12538
rect 2221 12486 2231 12538
rect 2255 12486 2285 12538
rect 2285 12486 2297 12538
rect 2297 12486 2311 12538
rect 2335 12486 2349 12538
rect 2349 12486 2361 12538
rect 2361 12486 2391 12538
rect 2415 12486 2425 12538
rect 2425 12486 2471 12538
rect 2175 12484 2231 12486
rect 2255 12484 2311 12486
rect 2335 12484 2391 12486
rect 2415 12484 2471 12486
rect 2175 11450 2231 11452
rect 2255 11450 2311 11452
rect 2335 11450 2391 11452
rect 2415 11450 2471 11452
rect 2175 11398 2221 11450
rect 2221 11398 2231 11450
rect 2255 11398 2285 11450
rect 2285 11398 2297 11450
rect 2297 11398 2311 11450
rect 2335 11398 2349 11450
rect 2349 11398 2361 11450
rect 2361 11398 2391 11450
rect 2415 11398 2425 11450
rect 2425 11398 2471 11450
rect 2175 11396 2231 11398
rect 2255 11396 2311 11398
rect 2335 11396 2391 11398
rect 2415 11396 2471 11398
rect 2175 10362 2231 10364
rect 2255 10362 2311 10364
rect 2335 10362 2391 10364
rect 2415 10362 2471 10364
rect 2175 10310 2221 10362
rect 2221 10310 2231 10362
rect 2255 10310 2285 10362
rect 2285 10310 2297 10362
rect 2297 10310 2311 10362
rect 2335 10310 2349 10362
rect 2349 10310 2361 10362
rect 2361 10310 2391 10362
rect 2415 10310 2425 10362
rect 2425 10310 2471 10362
rect 2175 10308 2231 10310
rect 2255 10308 2311 10310
rect 2335 10308 2391 10310
rect 2415 10308 2471 10310
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 4613 15802 4669 15804
rect 4693 15802 4749 15804
rect 4773 15802 4829 15804
rect 4853 15802 4909 15804
rect 4613 15750 4659 15802
rect 4659 15750 4669 15802
rect 4693 15750 4723 15802
rect 4723 15750 4735 15802
rect 4735 15750 4749 15802
rect 4773 15750 4787 15802
rect 4787 15750 4799 15802
rect 4799 15750 4829 15802
rect 4853 15750 4863 15802
rect 4863 15750 4909 15802
rect 4613 15748 4669 15750
rect 4693 15748 4749 15750
rect 4773 15748 4829 15750
rect 4853 15748 4909 15750
rect 7051 15802 7107 15804
rect 7131 15802 7187 15804
rect 7211 15802 7267 15804
rect 7291 15802 7347 15804
rect 7051 15750 7097 15802
rect 7097 15750 7107 15802
rect 7131 15750 7161 15802
rect 7161 15750 7173 15802
rect 7173 15750 7187 15802
rect 7211 15750 7225 15802
rect 7225 15750 7237 15802
rect 7237 15750 7267 15802
rect 7291 15750 7301 15802
rect 7301 15750 7347 15802
rect 7051 15748 7107 15750
rect 7131 15748 7187 15750
rect 7211 15748 7267 15750
rect 7291 15748 7347 15750
rect 11058 15952 11114 16008
rect 9489 15802 9545 15804
rect 9569 15802 9625 15804
rect 9649 15802 9705 15804
rect 9729 15802 9785 15804
rect 9489 15750 9535 15802
rect 9535 15750 9545 15802
rect 9569 15750 9599 15802
rect 9599 15750 9611 15802
rect 9611 15750 9625 15802
rect 9649 15750 9663 15802
rect 9663 15750 9675 15802
rect 9675 15750 9705 15802
rect 9729 15750 9739 15802
rect 9739 15750 9785 15802
rect 9489 15748 9545 15750
rect 9569 15748 9625 15750
rect 9649 15748 9705 15750
rect 9729 15748 9785 15750
rect 3394 15258 3450 15260
rect 3474 15258 3530 15260
rect 3554 15258 3610 15260
rect 3634 15258 3690 15260
rect 3394 15206 3440 15258
rect 3440 15206 3450 15258
rect 3474 15206 3504 15258
rect 3504 15206 3516 15258
rect 3516 15206 3530 15258
rect 3554 15206 3568 15258
rect 3568 15206 3580 15258
rect 3580 15206 3610 15258
rect 3634 15206 3644 15258
rect 3644 15206 3690 15258
rect 3394 15204 3450 15206
rect 3474 15204 3530 15206
rect 3554 15204 3610 15206
rect 3634 15204 3690 15206
rect 5832 15258 5888 15260
rect 5912 15258 5968 15260
rect 5992 15258 6048 15260
rect 6072 15258 6128 15260
rect 5832 15206 5878 15258
rect 5878 15206 5888 15258
rect 5912 15206 5942 15258
rect 5942 15206 5954 15258
rect 5954 15206 5968 15258
rect 5992 15206 6006 15258
rect 6006 15206 6018 15258
rect 6018 15206 6048 15258
rect 6072 15206 6082 15258
rect 6082 15206 6128 15258
rect 5832 15204 5888 15206
rect 5912 15204 5968 15206
rect 5992 15204 6048 15206
rect 6072 15204 6128 15206
rect 8270 15258 8326 15260
rect 8350 15258 8406 15260
rect 8430 15258 8486 15260
rect 8510 15258 8566 15260
rect 8270 15206 8316 15258
rect 8316 15206 8326 15258
rect 8350 15206 8380 15258
rect 8380 15206 8392 15258
rect 8392 15206 8406 15258
rect 8430 15206 8444 15258
rect 8444 15206 8456 15258
rect 8456 15206 8486 15258
rect 8510 15206 8520 15258
rect 8520 15206 8566 15258
rect 8270 15204 8326 15206
rect 8350 15204 8406 15206
rect 8430 15204 8486 15206
rect 8510 15204 8566 15206
rect 4613 14714 4669 14716
rect 4693 14714 4749 14716
rect 4773 14714 4829 14716
rect 4853 14714 4909 14716
rect 4613 14662 4659 14714
rect 4659 14662 4669 14714
rect 4693 14662 4723 14714
rect 4723 14662 4735 14714
rect 4735 14662 4749 14714
rect 4773 14662 4787 14714
rect 4787 14662 4799 14714
rect 4799 14662 4829 14714
rect 4853 14662 4863 14714
rect 4863 14662 4909 14714
rect 4613 14660 4669 14662
rect 4693 14660 4749 14662
rect 4773 14660 4829 14662
rect 4853 14660 4909 14662
rect 7051 14714 7107 14716
rect 7131 14714 7187 14716
rect 7211 14714 7267 14716
rect 7291 14714 7347 14716
rect 7051 14662 7097 14714
rect 7097 14662 7107 14714
rect 7131 14662 7161 14714
rect 7161 14662 7173 14714
rect 7173 14662 7187 14714
rect 7211 14662 7225 14714
rect 7225 14662 7237 14714
rect 7237 14662 7267 14714
rect 7291 14662 7301 14714
rect 7301 14662 7347 14714
rect 7051 14660 7107 14662
rect 7131 14660 7187 14662
rect 7211 14660 7267 14662
rect 7291 14660 7347 14662
rect 3394 14170 3450 14172
rect 3474 14170 3530 14172
rect 3554 14170 3610 14172
rect 3634 14170 3690 14172
rect 3394 14118 3440 14170
rect 3440 14118 3450 14170
rect 3474 14118 3504 14170
rect 3504 14118 3516 14170
rect 3516 14118 3530 14170
rect 3554 14118 3568 14170
rect 3568 14118 3580 14170
rect 3580 14118 3610 14170
rect 3634 14118 3644 14170
rect 3644 14118 3690 14170
rect 3394 14116 3450 14118
rect 3474 14116 3530 14118
rect 3554 14116 3610 14118
rect 3634 14116 3690 14118
rect 5832 14170 5888 14172
rect 5912 14170 5968 14172
rect 5992 14170 6048 14172
rect 6072 14170 6128 14172
rect 5832 14118 5878 14170
rect 5878 14118 5888 14170
rect 5912 14118 5942 14170
rect 5942 14118 5954 14170
rect 5954 14118 5968 14170
rect 5992 14118 6006 14170
rect 6006 14118 6018 14170
rect 6018 14118 6048 14170
rect 6072 14118 6082 14170
rect 6082 14118 6128 14170
rect 5832 14116 5888 14118
rect 5912 14116 5968 14118
rect 5992 14116 6048 14118
rect 6072 14116 6128 14118
rect 8270 14170 8326 14172
rect 8350 14170 8406 14172
rect 8430 14170 8486 14172
rect 8510 14170 8566 14172
rect 8270 14118 8316 14170
rect 8316 14118 8326 14170
rect 8350 14118 8380 14170
rect 8380 14118 8392 14170
rect 8392 14118 8406 14170
rect 8430 14118 8444 14170
rect 8444 14118 8456 14170
rect 8456 14118 8486 14170
rect 8510 14118 8520 14170
rect 8520 14118 8566 14170
rect 8270 14116 8326 14118
rect 8350 14116 8406 14118
rect 8430 14116 8486 14118
rect 8510 14116 8566 14118
rect 4613 13626 4669 13628
rect 4693 13626 4749 13628
rect 4773 13626 4829 13628
rect 4853 13626 4909 13628
rect 4613 13574 4659 13626
rect 4659 13574 4669 13626
rect 4693 13574 4723 13626
rect 4723 13574 4735 13626
rect 4735 13574 4749 13626
rect 4773 13574 4787 13626
rect 4787 13574 4799 13626
rect 4799 13574 4829 13626
rect 4853 13574 4863 13626
rect 4863 13574 4909 13626
rect 4613 13572 4669 13574
rect 4693 13572 4749 13574
rect 4773 13572 4829 13574
rect 4853 13572 4909 13574
rect 7051 13626 7107 13628
rect 7131 13626 7187 13628
rect 7211 13626 7267 13628
rect 7291 13626 7347 13628
rect 7051 13574 7097 13626
rect 7097 13574 7107 13626
rect 7131 13574 7161 13626
rect 7161 13574 7173 13626
rect 7173 13574 7187 13626
rect 7211 13574 7225 13626
rect 7225 13574 7237 13626
rect 7237 13574 7267 13626
rect 7291 13574 7301 13626
rect 7301 13574 7347 13626
rect 7051 13572 7107 13574
rect 7131 13572 7187 13574
rect 7211 13572 7267 13574
rect 7291 13572 7347 13574
rect 3394 13082 3450 13084
rect 3474 13082 3530 13084
rect 3554 13082 3610 13084
rect 3634 13082 3690 13084
rect 3394 13030 3440 13082
rect 3440 13030 3450 13082
rect 3474 13030 3504 13082
rect 3504 13030 3516 13082
rect 3516 13030 3530 13082
rect 3554 13030 3568 13082
rect 3568 13030 3580 13082
rect 3580 13030 3610 13082
rect 3634 13030 3644 13082
rect 3644 13030 3690 13082
rect 3394 13028 3450 13030
rect 3474 13028 3530 13030
rect 3554 13028 3610 13030
rect 3634 13028 3690 13030
rect 5832 13082 5888 13084
rect 5912 13082 5968 13084
rect 5992 13082 6048 13084
rect 6072 13082 6128 13084
rect 5832 13030 5878 13082
rect 5878 13030 5888 13082
rect 5912 13030 5942 13082
rect 5942 13030 5954 13082
rect 5954 13030 5968 13082
rect 5992 13030 6006 13082
rect 6006 13030 6018 13082
rect 6018 13030 6048 13082
rect 6072 13030 6082 13082
rect 6082 13030 6128 13082
rect 5832 13028 5888 13030
rect 5912 13028 5968 13030
rect 5992 13028 6048 13030
rect 6072 13028 6128 13030
rect 8270 13082 8326 13084
rect 8350 13082 8406 13084
rect 8430 13082 8486 13084
rect 8510 13082 8566 13084
rect 8270 13030 8316 13082
rect 8316 13030 8326 13082
rect 8350 13030 8380 13082
rect 8380 13030 8392 13082
rect 8392 13030 8406 13082
rect 8430 13030 8444 13082
rect 8444 13030 8456 13082
rect 8456 13030 8486 13082
rect 8510 13030 8520 13082
rect 8520 13030 8566 13082
rect 8270 13028 8326 13030
rect 8350 13028 8406 13030
rect 8430 13028 8486 13030
rect 8510 13028 8566 13030
rect 4613 12538 4669 12540
rect 4693 12538 4749 12540
rect 4773 12538 4829 12540
rect 4853 12538 4909 12540
rect 4613 12486 4659 12538
rect 4659 12486 4669 12538
rect 4693 12486 4723 12538
rect 4723 12486 4735 12538
rect 4735 12486 4749 12538
rect 4773 12486 4787 12538
rect 4787 12486 4799 12538
rect 4799 12486 4829 12538
rect 4853 12486 4863 12538
rect 4863 12486 4909 12538
rect 4613 12484 4669 12486
rect 4693 12484 4749 12486
rect 4773 12484 4829 12486
rect 4853 12484 4909 12486
rect 7051 12538 7107 12540
rect 7131 12538 7187 12540
rect 7211 12538 7267 12540
rect 7291 12538 7347 12540
rect 7051 12486 7097 12538
rect 7097 12486 7107 12538
rect 7131 12486 7161 12538
rect 7161 12486 7173 12538
rect 7173 12486 7187 12538
rect 7211 12486 7225 12538
rect 7225 12486 7237 12538
rect 7237 12486 7267 12538
rect 7291 12486 7301 12538
rect 7301 12486 7347 12538
rect 7051 12484 7107 12486
rect 7131 12484 7187 12486
rect 7211 12484 7267 12486
rect 7291 12484 7347 12486
rect 3394 11994 3450 11996
rect 3474 11994 3530 11996
rect 3554 11994 3610 11996
rect 3634 11994 3690 11996
rect 3394 11942 3440 11994
rect 3440 11942 3450 11994
rect 3474 11942 3504 11994
rect 3504 11942 3516 11994
rect 3516 11942 3530 11994
rect 3554 11942 3568 11994
rect 3568 11942 3580 11994
rect 3580 11942 3610 11994
rect 3634 11942 3644 11994
rect 3644 11942 3690 11994
rect 3394 11940 3450 11942
rect 3474 11940 3530 11942
rect 3554 11940 3610 11942
rect 3634 11940 3690 11942
rect 5832 11994 5888 11996
rect 5912 11994 5968 11996
rect 5992 11994 6048 11996
rect 6072 11994 6128 11996
rect 5832 11942 5878 11994
rect 5878 11942 5888 11994
rect 5912 11942 5942 11994
rect 5942 11942 5954 11994
rect 5954 11942 5968 11994
rect 5992 11942 6006 11994
rect 6006 11942 6018 11994
rect 6018 11942 6048 11994
rect 6072 11942 6082 11994
rect 6082 11942 6128 11994
rect 5832 11940 5888 11942
rect 5912 11940 5968 11942
rect 5992 11940 6048 11942
rect 6072 11940 6128 11942
rect 8270 11994 8326 11996
rect 8350 11994 8406 11996
rect 8430 11994 8486 11996
rect 8510 11994 8566 11996
rect 8270 11942 8316 11994
rect 8316 11942 8326 11994
rect 8350 11942 8380 11994
rect 8380 11942 8392 11994
rect 8392 11942 8406 11994
rect 8430 11942 8444 11994
rect 8444 11942 8456 11994
rect 8456 11942 8486 11994
rect 8510 11942 8520 11994
rect 8520 11942 8566 11994
rect 8270 11940 8326 11942
rect 8350 11940 8406 11942
rect 8430 11940 8486 11942
rect 8510 11940 8566 11942
rect 4613 11450 4669 11452
rect 4693 11450 4749 11452
rect 4773 11450 4829 11452
rect 4853 11450 4909 11452
rect 4613 11398 4659 11450
rect 4659 11398 4669 11450
rect 4693 11398 4723 11450
rect 4723 11398 4735 11450
rect 4735 11398 4749 11450
rect 4773 11398 4787 11450
rect 4787 11398 4799 11450
rect 4799 11398 4829 11450
rect 4853 11398 4863 11450
rect 4863 11398 4909 11450
rect 4613 11396 4669 11398
rect 4693 11396 4749 11398
rect 4773 11396 4829 11398
rect 4853 11396 4909 11398
rect 3394 10906 3450 10908
rect 3474 10906 3530 10908
rect 3554 10906 3610 10908
rect 3634 10906 3690 10908
rect 3394 10854 3440 10906
rect 3440 10854 3450 10906
rect 3474 10854 3504 10906
rect 3504 10854 3516 10906
rect 3516 10854 3530 10906
rect 3554 10854 3568 10906
rect 3568 10854 3580 10906
rect 3580 10854 3610 10906
rect 3634 10854 3644 10906
rect 3644 10854 3690 10906
rect 3394 10852 3450 10854
rect 3474 10852 3530 10854
rect 3554 10852 3610 10854
rect 3634 10852 3690 10854
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 4613 10362 4669 10364
rect 4693 10362 4749 10364
rect 4773 10362 4829 10364
rect 4853 10362 4909 10364
rect 4613 10310 4659 10362
rect 4659 10310 4669 10362
rect 4693 10310 4723 10362
rect 4723 10310 4735 10362
rect 4735 10310 4749 10362
rect 4773 10310 4787 10362
rect 4787 10310 4799 10362
rect 4799 10310 4829 10362
rect 4853 10310 4863 10362
rect 4863 10310 4909 10362
rect 4613 10308 4669 10310
rect 4693 10308 4749 10310
rect 4773 10308 4829 10310
rect 4853 10308 4909 10310
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 5832 10906 5888 10908
rect 5912 10906 5968 10908
rect 5992 10906 6048 10908
rect 6072 10906 6128 10908
rect 5832 10854 5878 10906
rect 5878 10854 5888 10906
rect 5912 10854 5942 10906
rect 5942 10854 5954 10906
rect 5954 10854 5968 10906
rect 5992 10854 6006 10906
rect 6006 10854 6018 10906
rect 6018 10854 6048 10906
rect 6072 10854 6082 10906
rect 6082 10854 6128 10906
rect 5832 10852 5888 10854
rect 5912 10852 5968 10854
rect 5992 10852 6048 10854
rect 6072 10852 6128 10854
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 7051 11450 7107 11452
rect 7131 11450 7187 11452
rect 7211 11450 7267 11452
rect 7291 11450 7347 11452
rect 7051 11398 7097 11450
rect 7097 11398 7107 11450
rect 7131 11398 7161 11450
rect 7161 11398 7173 11450
rect 7173 11398 7187 11450
rect 7211 11398 7225 11450
rect 7225 11398 7237 11450
rect 7237 11398 7267 11450
rect 7291 11398 7301 11450
rect 7301 11398 7347 11450
rect 7051 11396 7107 11398
rect 7131 11396 7187 11398
rect 7211 11396 7267 11398
rect 7291 11396 7347 11398
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 7051 10362 7107 10364
rect 7131 10362 7187 10364
rect 7211 10362 7267 10364
rect 7291 10362 7347 10364
rect 7051 10310 7097 10362
rect 7097 10310 7107 10362
rect 7131 10310 7161 10362
rect 7161 10310 7173 10362
rect 7173 10310 7187 10362
rect 7211 10310 7225 10362
rect 7225 10310 7237 10362
rect 7237 10310 7267 10362
rect 7291 10310 7301 10362
rect 7301 10310 7347 10362
rect 7051 10308 7107 10310
rect 7131 10308 7187 10310
rect 7211 10308 7267 10310
rect 7291 10308 7347 10310
rect 8270 10906 8326 10908
rect 8350 10906 8406 10908
rect 8430 10906 8486 10908
rect 8510 10906 8566 10908
rect 8270 10854 8316 10906
rect 8316 10854 8326 10906
rect 8350 10854 8380 10906
rect 8380 10854 8392 10906
rect 8392 10854 8406 10906
rect 8430 10854 8444 10906
rect 8444 10854 8456 10906
rect 8456 10854 8486 10906
rect 8510 10854 8520 10906
rect 8520 10854 8566 10906
rect 8270 10852 8326 10854
rect 8350 10852 8406 10854
rect 8430 10852 8486 10854
rect 8510 10852 8566 10854
rect 9489 14714 9545 14716
rect 9569 14714 9625 14716
rect 9649 14714 9705 14716
rect 9729 14714 9785 14716
rect 9489 14662 9535 14714
rect 9535 14662 9545 14714
rect 9569 14662 9599 14714
rect 9599 14662 9611 14714
rect 9611 14662 9625 14714
rect 9649 14662 9663 14714
rect 9663 14662 9675 14714
rect 9675 14662 9705 14714
rect 9729 14662 9739 14714
rect 9739 14662 9785 14714
rect 9489 14660 9545 14662
rect 9569 14660 9625 14662
rect 9649 14660 9705 14662
rect 9729 14660 9785 14662
rect 9489 13626 9545 13628
rect 9569 13626 9625 13628
rect 9649 13626 9705 13628
rect 9729 13626 9785 13628
rect 9489 13574 9535 13626
rect 9535 13574 9545 13626
rect 9569 13574 9599 13626
rect 9599 13574 9611 13626
rect 9611 13574 9625 13626
rect 9649 13574 9663 13626
rect 9663 13574 9675 13626
rect 9675 13574 9705 13626
rect 9729 13574 9739 13626
rect 9739 13574 9785 13626
rect 9489 13572 9545 13574
rect 9569 13572 9625 13574
rect 9649 13572 9705 13574
rect 9729 13572 9785 13574
rect 9489 12538 9545 12540
rect 9569 12538 9625 12540
rect 9649 12538 9705 12540
rect 9729 12538 9785 12540
rect 9489 12486 9535 12538
rect 9535 12486 9545 12538
rect 9569 12486 9599 12538
rect 9599 12486 9611 12538
rect 9611 12486 9625 12538
rect 9649 12486 9663 12538
rect 9663 12486 9675 12538
rect 9675 12486 9705 12538
rect 9729 12486 9739 12538
rect 9739 12486 9785 12538
rect 9489 12484 9545 12486
rect 9569 12484 9625 12486
rect 9649 12484 9705 12486
rect 9729 12484 9785 12486
rect 9489 11450 9545 11452
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9489 11398 9535 11450
rect 9535 11398 9545 11450
rect 9569 11398 9599 11450
rect 9599 11398 9611 11450
rect 9611 11398 9625 11450
rect 9649 11398 9663 11450
rect 9663 11398 9675 11450
rect 9675 11398 9705 11450
rect 9729 11398 9739 11450
rect 9739 11398 9785 11450
rect 9489 11396 9545 11398
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 9489 10362 9545 10364
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9489 10310 9535 10362
rect 9535 10310 9545 10362
rect 9569 10310 9599 10362
rect 9599 10310 9611 10362
rect 9611 10310 9625 10362
rect 9649 10310 9663 10362
rect 9663 10310 9675 10362
rect 9675 10310 9705 10362
rect 9729 10310 9739 10362
rect 9739 10310 9785 10362
rect 9489 10308 9545 10310
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 10708 15258 10764 15260
rect 10788 15258 10844 15260
rect 10868 15258 10924 15260
rect 10948 15258 11004 15260
rect 10708 15206 10754 15258
rect 10754 15206 10764 15258
rect 10788 15206 10818 15258
rect 10818 15206 10830 15258
rect 10830 15206 10844 15258
rect 10868 15206 10882 15258
rect 10882 15206 10894 15258
rect 10894 15206 10924 15258
rect 10948 15206 10958 15258
rect 10958 15206 11004 15258
rect 10708 15204 10764 15206
rect 10788 15204 10844 15206
rect 10868 15204 10924 15206
rect 10948 15204 11004 15206
rect 10708 14170 10764 14172
rect 10788 14170 10844 14172
rect 10868 14170 10924 14172
rect 10948 14170 11004 14172
rect 10708 14118 10754 14170
rect 10754 14118 10764 14170
rect 10788 14118 10818 14170
rect 10818 14118 10830 14170
rect 10830 14118 10844 14170
rect 10868 14118 10882 14170
rect 10882 14118 10894 14170
rect 10894 14118 10924 14170
rect 10948 14118 10958 14170
rect 10958 14118 11004 14170
rect 10708 14116 10764 14118
rect 10788 14116 10844 14118
rect 10868 14116 10924 14118
rect 10948 14116 11004 14118
rect 10708 13082 10764 13084
rect 10788 13082 10844 13084
rect 10868 13082 10924 13084
rect 10948 13082 11004 13084
rect 10708 13030 10754 13082
rect 10754 13030 10764 13082
rect 10788 13030 10818 13082
rect 10818 13030 10830 13082
rect 10830 13030 10844 13082
rect 10868 13030 10882 13082
rect 10882 13030 10894 13082
rect 10894 13030 10924 13082
rect 10948 13030 10958 13082
rect 10958 13030 11004 13082
rect 10708 13028 10764 13030
rect 10788 13028 10844 13030
rect 10868 13028 10924 13030
rect 10948 13028 11004 13030
rect 10230 12416 10286 12472
rect 10708 11994 10764 11996
rect 10788 11994 10844 11996
rect 10868 11994 10924 11996
rect 10948 11994 11004 11996
rect 10708 11942 10754 11994
rect 10754 11942 10764 11994
rect 10788 11942 10818 11994
rect 10818 11942 10830 11994
rect 10830 11942 10844 11994
rect 10868 11942 10882 11994
rect 10882 11942 10894 11994
rect 10894 11942 10924 11994
rect 10948 11942 10958 11994
rect 10958 11942 11004 11994
rect 10708 11940 10764 11942
rect 10788 11940 10844 11942
rect 10868 11940 10924 11942
rect 10948 11940 11004 11942
rect 10708 10906 10764 10908
rect 10788 10906 10844 10908
rect 10868 10906 10924 10908
rect 10948 10906 11004 10908
rect 10708 10854 10754 10906
rect 10754 10854 10764 10906
rect 10788 10854 10818 10906
rect 10818 10854 10830 10906
rect 10830 10854 10844 10906
rect 10868 10854 10882 10906
rect 10882 10854 10894 10906
rect 10894 10854 10924 10906
rect 10948 10854 10958 10906
rect 10958 10854 11004 10906
rect 10708 10852 10764 10854
rect 10788 10852 10844 10854
rect 10868 10852 10924 10854
rect 10948 10852 11004 10854
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10230 8900 10286 8936
rect 10230 8880 10232 8900
rect 10232 8880 10284 8900
rect 10284 8880 10286 8900
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 10230 5636 10286 5672
rect 10230 5616 10232 5636
rect 10232 5616 10284 5636
rect 10284 5616 10286 5636
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 10230 1808 10286 1864
<< metal3 >>
rect 11053 16010 11119 16013
rect 11200 16010 12000 16040
rect 11053 16008 12000 16010
rect 11053 15952 11058 16008
rect 11114 15952 12000 16008
rect 11053 15950 12000 15952
rect 11053 15947 11119 15950
rect 11200 15920 12000 15950
rect 2165 15808 2481 15809
rect 2165 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2481 15808
rect 2165 15743 2481 15744
rect 4603 15808 4919 15809
rect 4603 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4919 15808
rect 4603 15743 4919 15744
rect 7041 15808 7357 15809
rect 7041 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7357 15808
rect 7041 15743 7357 15744
rect 9479 15808 9795 15809
rect 9479 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9795 15808
rect 9479 15743 9795 15744
rect 3384 15264 3700 15265
rect 3384 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3700 15264
rect 3384 15199 3700 15200
rect 5822 15264 6138 15265
rect 5822 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6138 15264
rect 5822 15199 6138 15200
rect 8260 15264 8576 15265
rect 8260 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8576 15264
rect 8260 15199 8576 15200
rect 10698 15264 11014 15265
rect 10698 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11014 15264
rect 10698 15199 11014 15200
rect 2165 14720 2481 14721
rect 2165 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2481 14720
rect 2165 14655 2481 14656
rect 4603 14720 4919 14721
rect 4603 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4919 14720
rect 4603 14655 4919 14656
rect 7041 14720 7357 14721
rect 7041 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7357 14720
rect 7041 14655 7357 14656
rect 9479 14720 9795 14721
rect 9479 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9795 14720
rect 9479 14655 9795 14656
rect 3384 14176 3700 14177
rect 3384 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3700 14176
rect 3384 14111 3700 14112
rect 5822 14176 6138 14177
rect 5822 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6138 14176
rect 5822 14111 6138 14112
rect 8260 14176 8576 14177
rect 8260 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8576 14176
rect 8260 14111 8576 14112
rect 10698 14176 11014 14177
rect 10698 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11014 14176
rect 10698 14111 11014 14112
rect 2165 13632 2481 13633
rect 2165 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2481 13632
rect 2165 13567 2481 13568
rect 4603 13632 4919 13633
rect 4603 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4919 13632
rect 4603 13567 4919 13568
rect 7041 13632 7357 13633
rect 7041 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7357 13632
rect 7041 13567 7357 13568
rect 9479 13632 9795 13633
rect 9479 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9795 13632
rect 9479 13567 9795 13568
rect 3384 13088 3700 13089
rect 3384 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3700 13088
rect 3384 13023 3700 13024
rect 5822 13088 6138 13089
rect 5822 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6138 13088
rect 5822 13023 6138 13024
rect 8260 13088 8576 13089
rect 8260 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8576 13088
rect 8260 13023 8576 13024
rect 10698 13088 11014 13089
rect 10698 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11014 13088
rect 10698 13023 11014 13024
rect 2165 12544 2481 12545
rect 2165 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2481 12544
rect 2165 12479 2481 12480
rect 4603 12544 4919 12545
rect 4603 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4919 12544
rect 4603 12479 4919 12480
rect 7041 12544 7357 12545
rect 7041 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7357 12544
rect 7041 12479 7357 12480
rect 9479 12544 9795 12545
rect 9479 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9795 12544
rect 9479 12479 9795 12480
rect 10225 12474 10291 12477
rect 11200 12474 12000 12504
rect 10225 12472 12000 12474
rect 10225 12416 10230 12472
rect 10286 12416 12000 12472
rect 10225 12414 12000 12416
rect 10225 12411 10291 12414
rect 11200 12384 12000 12414
rect 3384 12000 3700 12001
rect 3384 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3700 12000
rect 3384 11935 3700 11936
rect 5822 12000 6138 12001
rect 5822 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6138 12000
rect 5822 11935 6138 11936
rect 8260 12000 8576 12001
rect 8260 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8576 12000
rect 8260 11935 8576 11936
rect 10698 12000 11014 12001
rect 10698 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11014 12000
rect 10698 11935 11014 11936
rect 2165 11456 2481 11457
rect 2165 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2481 11456
rect 2165 11391 2481 11392
rect 4603 11456 4919 11457
rect 4603 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4919 11456
rect 4603 11391 4919 11392
rect 7041 11456 7357 11457
rect 7041 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7357 11456
rect 7041 11391 7357 11392
rect 9479 11456 9795 11457
rect 9479 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9795 11456
rect 9479 11391 9795 11392
rect 3384 10912 3700 10913
rect 3384 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3700 10912
rect 3384 10847 3700 10848
rect 5822 10912 6138 10913
rect 5822 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6138 10912
rect 5822 10847 6138 10848
rect 8260 10912 8576 10913
rect 8260 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8576 10912
rect 8260 10847 8576 10848
rect 10698 10912 11014 10913
rect 10698 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11014 10912
rect 10698 10847 11014 10848
rect 2165 10368 2481 10369
rect 2165 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2481 10368
rect 2165 10303 2481 10304
rect 4603 10368 4919 10369
rect 4603 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4919 10368
rect 4603 10303 4919 10304
rect 7041 10368 7357 10369
rect 7041 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7357 10368
rect 7041 10303 7357 10304
rect 9479 10368 9795 10369
rect 9479 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9795 10368
rect 9479 10303 9795 10304
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 10225 8938 10291 8941
rect 11200 8938 12000 8968
rect 10225 8936 12000 8938
rect 10225 8880 10230 8936
rect 10286 8880 12000 8936
rect 10225 8878 12000 8880
rect 10225 8875 10291 8878
rect 11200 8848 12000 8878
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 10225 5674 10291 5677
rect 10225 5672 11346 5674
rect 10225 5616 10230 5672
rect 10286 5616 11346 5672
rect 10225 5614 11346 5616
rect 10225 5611 10291 5614
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 11286 5432 11346 5614
rect 10698 5407 11014 5408
rect 11200 5312 12000 5432
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 10225 1866 10291 1869
rect 11200 1866 12000 1896
rect 10225 1864 12000 1866
rect 10225 1808 10230 1864
rect 10286 1808 12000 1864
rect 10225 1806 12000 1808
rect 10225 1803 10291 1806
rect 11200 1776 12000 1806
<< via3 >>
rect 2171 15804 2235 15808
rect 2171 15748 2175 15804
rect 2175 15748 2231 15804
rect 2231 15748 2235 15804
rect 2171 15744 2235 15748
rect 2251 15804 2315 15808
rect 2251 15748 2255 15804
rect 2255 15748 2311 15804
rect 2311 15748 2315 15804
rect 2251 15744 2315 15748
rect 2331 15804 2395 15808
rect 2331 15748 2335 15804
rect 2335 15748 2391 15804
rect 2391 15748 2395 15804
rect 2331 15744 2395 15748
rect 2411 15804 2475 15808
rect 2411 15748 2415 15804
rect 2415 15748 2471 15804
rect 2471 15748 2475 15804
rect 2411 15744 2475 15748
rect 4609 15804 4673 15808
rect 4609 15748 4613 15804
rect 4613 15748 4669 15804
rect 4669 15748 4673 15804
rect 4609 15744 4673 15748
rect 4689 15804 4753 15808
rect 4689 15748 4693 15804
rect 4693 15748 4749 15804
rect 4749 15748 4753 15804
rect 4689 15744 4753 15748
rect 4769 15804 4833 15808
rect 4769 15748 4773 15804
rect 4773 15748 4829 15804
rect 4829 15748 4833 15804
rect 4769 15744 4833 15748
rect 4849 15804 4913 15808
rect 4849 15748 4853 15804
rect 4853 15748 4909 15804
rect 4909 15748 4913 15804
rect 4849 15744 4913 15748
rect 7047 15804 7111 15808
rect 7047 15748 7051 15804
rect 7051 15748 7107 15804
rect 7107 15748 7111 15804
rect 7047 15744 7111 15748
rect 7127 15804 7191 15808
rect 7127 15748 7131 15804
rect 7131 15748 7187 15804
rect 7187 15748 7191 15804
rect 7127 15744 7191 15748
rect 7207 15804 7271 15808
rect 7207 15748 7211 15804
rect 7211 15748 7267 15804
rect 7267 15748 7271 15804
rect 7207 15744 7271 15748
rect 7287 15804 7351 15808
rect 7287 15748 7291 15804
rect 7291 15748 7347 15804
rect 7347 15748 7351 15804
rect 7287 15744 7351 15748
rect 9485 15804 9549 15808
rect 9485 15748 9489 15804
rect 9489 15748 9545 15804
rect 9545 15748 9549 15804
rect 9485 15744 9549 15748
rect 9565 15804 9629 15808
rect 9565 15748 9569 15804
rect 9569 15748 9625 15804
rect 9625 15748 9629 15804
rect 9565 15744 9629 15748
rect 9645 15804 9709 15808
rect 9645 15748 9649 15804
rect 9649 15748 9705 15804
rect 9705 15748 9709 15804
rect 9645 15744 9709 15748
rect 9725 15804 9789 15808
rect 9725 15748 9729 15804
rect 9729 15748 9785 15804
rect 9785 15748 9789 15804
rect 9725 15744 9789 15748
rect 3390 15260 3454 15264
rect 3390 15204 3394 15260
rect 3394 15204 3450 15260
rect 3450 15204 3454 15260
rect 3390 15200 3454 15204
rect 3470 15260 3534 15264
rect 3470 15204 3474 15260
rect 3474 15204 3530 15260
rect 3530 15204 3534 15260
rect 3470 15200 3534 15204
rect 3550 15260 3614 15264
rect 3550 15204 3554 15260
rect 3554 15204 3610 15260
rect 3610 15204 3614 15260
rect 3550 15200 3614 15204
rect 3630 15260 3694 15264
rect 3630 15204 3634 15260
rect 3634 15204 3690 15260
rect 3690 15204 3694 15260
rect 3630 15200 3694 15204
rect 5828 15260 5892 15264
rect 5828 15204 5832 15260
rect 5832 15204 5888 15260
rect 5888 15204 5892 15260
rect 5828 15200 5892 15204
rect 5908 15260 5972 15264
rect 5908 15204 5912 15260
rect 5912 15204 5968 15260
rect 5968 15204 5972 15260
rect 5908 15200 5972 15204
rect 5988 15260 6052 15264
rect 5988 15204 5992 15260
rect 5992 15204 6048 15260
rect 6048 15204 6052 15260
rect 5988 15200 6052 15204
rect 6068 15260 6132 15264
rect 6068 15204 6072 15260
rect 6072 15204 6128 15260
rect 6128 15204 6132 15260
rect 6068 15200 6132 15204
rect 8266 15260 8330 15264
rect 8266 15204 8270 15260
rect 8270 15204 8326 15260
rect 8326 15204 8330 15260
rect 8266 15200 8330 15204
rect 8346 15260 8410 15264
rect 8346 15204 8350 15260
rect 8350 15204 8406 15260
rect 8406 15204 8410 15260
rect 8346 15200 8410 15204
rect 8426 15260 8490 15264
rect 8426 15204 8430 15260
rect 8430 15204 8486 15260
rect 8486 15204 8490 15260
rect 8426 15200 8490 15204
rect 8506 15260 8570 15264
rect 8506 15204 8510 15260
rect 8510 15204 8566 15260
rect 8566 15204 8570 15260
rect 8506 15200 8570 15204
rect 10704 15260 10768 15264
rect 10704 15204 10708 15260
rect 10708 15204 10764 15260
rect 10764 15204 10768 15260
rect 10704 15200 10768 15204
rect 10784 15260 10848 15264
rect 10784 15204 10788 15260
rect 10788 15204 10844 15260
rect 10844 15204 10848 15260
rect 10784 15200 10848 15204
rect 10864 15260 10928 15264
rect 10864 15204 10868 15260
rect 10868 15204 10924 15260
rect 10924 15204 10928 15260
rect 10864 15200 10928 15204
rect 10944 15260 11008 15264
rect 10944 15204 10948 15260
rect 10948 15204 11004 15260
rect 11004 15204 11008 15260
rect 10944 15200 11008 15204
rect 2171 14716 2235 14720
rect 2171 14660 2175 14716
rect 2175 14660 2231 14716
rect 2231 14660 2235 14716
rect 2171 14656 2235 14660
rect 2251 14716 2315 14720
rect 2251 14660 2255 14716
rect 2255 14660 2311 14716
rect 2311 14660 2315 14716
rect 2251 14656 2315 14660
rect 2331 14716 2395 14720
rect 2331 14660 2335 14716
rect 2335 14660 2391 14716
rect 2391 14660 2395 14716
rect 2331 14656 2395 14660
rect 2411 14716 2475 14720
rect 2411 14660 2415 14716
rect 2415 14660 2471 14716
rect 2471 14660 2475 14716
rect 2411 14656 2475 14660
rect 4609 14716 4673 14720
rect 4609 14660 4613 14716
rect 4613 14660 4669 14716
rect 4669 14660 4673 14716
rect 4609 14656 4673 14660
rect 4689 14716 4753 14720
rect 4689 14660 4693 14716
rect 4693 14660 4749 14716
rect 4749 14660 4753 14716
rect 4689 14656 4753 14660
rect 4769 14716 4833 14720
rect 4769 14660 4773 14716
rect 4773 14660 4829 14716
rect 4829 14660 4833 14716
rect 4769 14656 4833 14660
rect 4849 14716 4913 14720
rect 4849 14660 4853 14716
rect 4853 14660 4909 14716
rect 4909 14660 4913 14716
rect 4849 14656 4913 14660
rect 7047 14716 7111 14720
rect 7047 14660 7051 14716
rect 7051 14660 7107 14716
rect 7107 14660 7111 14716
rect 7047 14656 7111 14660
rect 7127 14716 7191 14720
rect 7127 14660 7131 14716
rect 7131 14660 7187 14716
rect 7187 14660 7191 14716
rect 7127 14656 7191 14660
rect 7207 14716 7271 14720
rect 7207 14660 7211 14716
rect 7211 14660 7267 14716
rect 7267 14660 7271 14716
rect 7207 14656 7271 14660
rect 7287 14716 7351 14720
rect 7287 14660 7291 14716
rect 7291 14660 7347 14716
rect 7347 14660 7351 14716
rect 7287 14656 7351 14660
rect 9485 14716 9549 14720
rect 9485 14660 9489 14716
rect 9489 14660 9545 14716
rect 9545 14660 9549 14716
rect 9485 14656 9549 14660
rect 9565 14716 9629 14720
rect 9565 14660 9569 14716
rect 9569 14660 9625 14716
rect 9625 14660 9629 14716
rect 9565 14656 9629 14660
rect 9645 14716 9709 14720
rect 9645 14660 9649 14716
rect 9649 14660 9705 14716
rect 9705 14660 9709 14716
rect 9645 14656 9709 14660
rect 9725 14716 9789 14720
rect 9725 14660 9729 14716
rect 9729 14660 9785 14716
rect 9785 14660 9789 14716
rect 9725 14656 9789 14660
rect 3390 14172 3454 14176
rect 3390 14116 3394 14172
rect 3394 14116 3450 14172
rect 3450 14116 3454 14172
rect 3390 14112 3454 14116
rect 3470 14172 3534 14176
rect 3470 14116 3474 14172
rect 3474 14116 3530 14172
rect 3530 14116 3534 14172
rect 3470 14112 3534 14116
rect 3550 14172 3614 14176
rect 3550 14116 3554 14172
rect 3554 14116 3610 14172
rect 3610 14116 3614 14172
rect 3550 14112 3614 14116
rect 3630 14172 3694 14176
rect 3630 14116 3634 14172
rect 3634 14116 3690 14172
rect 3690 14116 3694 14172
rect 3630 14112 3694 14116
rect 5828 14172 5892 14176
rect 5828 14116 5832 14172
rect 5832 14116 5888 14172
rect 5888 14116 5892 14172
rect 5828 14112 5892 14116
rect 5908 14172 5972 14176
rect 5908 14116 5912 14172
rect 5912 14116 5968 14172
rect 5968 14116 5972 14172
rect 5908 14112 5972 14116
rect 5988 14172 6052 14176
rect 5988 14116 5992 14172
rect 5992 14116 6048 14172
rect 6048 14116 6052 14172
rect 5988 14112 6052 14116
rect 6068 14172 6132 14176
rect 6068 14116 6072 14172
rect 6072 14116 6128 14172
rect 6128 14116 6132 14172
rect 6068 14112 6132 14116
rect 8266 14172 8330 14176
rect 8266 14116 8270 14172
rect 8270 14116 8326 14172
rect 8326 14116 8330 14172
rect 8266 14112 8330 14116
rect 8346 14172 8410 14176
rect 8346 14116 8350 14172
rect 8350 14116 8406 14172
rect 8406 14116 8410 14172
rect 8346 14112 8410 14116
rect 8426 14172 8490 14176
rect 8426 14116 8430 14172
rect 8430 14116 8486 14172
rect 8486 14116 8490 14172
rect 8426 14112 8490 14116
rect 8506 14172 8570 14176
rect 8506 14116 8510 14172
rect 8510 14116 8566 14172
rect 8566 14116 8570 14172
rect 8506 14112 8570 14116
rect 10704 14172 10768 14176
rect 10704 14116 10708 14172
rect 10708 14116 10764 14172
rect 10764 14116 10768 14172
rect 10704 14112 10768 14116
rect 10784 14172 10848 14176
rect 10784 14116 10788 14172
rect 10788 14116 10844 14172
rect 10844 14116 10848 14172
rect 10784 14112 10848 14116
rect 10864 14172 10928 14176
rect 10864 14116 10868 14172
rect 10868 14116 10924 14172
rect 10924 14116 10928 14172
rect 10864 14112 10928 14116
rect 10944 14172 11008 14176
rect 10944 14116 10948 14172
rect 10948 14116 11004 14172
rect 11004 14116 11008 14172
rect 10944 14112 11008 14116
rect 2171 13628 2235 13632
rect 2171 13572 2175 13628
rect 2175 13572 2231 13628
rect 2231 13572 2235 13628
rect 2171 13568 2235 13572
rect 2251 13628 2315 13632
rect 2251 13572 2255 13628
rect 2255 13572 2311 13628
rect 2311 13572 2315 13628
rect 2251 13568 2315 13572
rect 2331 13628 2395 13632
rect 2331 13572 2335 13628
rect 2335 13572 2391 13628
rect 2391 13572 2395 13628
rect 2331 13568 2395 13572
rect 2411 13628 2475 13632
rect 2411 13572 2415 13628
rect 2415 13572 2471 13628
rect 2471 13572 2475 13628
rect 2411 13568 2475 13572
rect 4609 13628 4673 13632
rect 4609 13572 4613 13628
rect 4613 13572 4669 13628
rect 4669 13572 4673 13628
rect 4609 13568 4673 13572
rect 4689 13628 4753 13632
rect 4689 13572 4693 13628
rect 4693 13572 4749 13628
rect 4749 13572 4753 13628
rect 4689 13568 4753 13572
rect 4769 13628 4833 13632
rect 4769 13572 4773 13628
rect 4773 13572 4829 13628
rect 4829 13572 4833 13628
rect 4769 13568 4833 13572
rect 4849 13628 4913 13632
rect 4849 13572 4853 13628
rect 4853 13572 4909 13628
rect 4909 13572 4913 13628
rect 4849 13568 4913 13572
rect 7047 13628 7111 13632
rect 7047 13572 7051 13628
rect 7051 13572 7107 13628
rect 7107 13572 7111 13628
rect 7047 13568 7111 13572
rect 7127 13628 7191 13632
rect 7127 13572 7131 13628
rect 7131 13572 7187 13628
rect 7187 13572 7191 13628
rect 7127 13568 7191 13572
rect 7207 13628 7271 13632
rect 7207 13572 7211 13628
rect 7211 13572 7267 13628
rect 7267 13572 7271 13628
rect 7207 13568 7271 13572
rect 7287 13628 7351 13632
rect 7287 13572 7291 13628
rect 7291 13572 7347 13628
rect 7347 13572 7351 13628
rect 7287 13568 7351 13572
rect 9485 13628 9549 13632
rect 9485 13572 9489 13628
rect 9489 13572 9545 13628
rect 9545 13572 9549 13628
rect 9485 13568 9549 13572
rect 9565 13628 9629 13632
rect 9565 13572 9569 13628
rect 9569 13572 9625 13628
rect 9625 13572 9629 13628
rect 9565 13568 9629 13572
rect 9645 13628 9709 13632
rect 9645 13572 9649 13628
rect 9649 13572 9705 13628
rect 9705 13572 9709 13628
rect 9645 13568 9709 13572
rect 9725 13628 9789 13632
rect 9725 13572 9729 13628
rect 9729 13572 9785 13628
rect 9785 13572 9789 13628
rect 9725 13568 9789 13572
rect 3390 13084 3454 13088
rect 3390 13028 3394 13084
rect 3394 13028 3450 13084
rect 3450 13028 3454 13084
rect 3390 13024 3454 13028
rect 3470 13084 3534 13088
rect 3470 13028 3474 13084
rect 3474 13028 3530 13084
rect 3530 13028 3534 13084
rect 3470 13024 3534 13028
rect 3550 13084 3614 13088
rect 3550 13028 3554 13084
rect 3554 13028 3610 13084
rect 3610 13028 3614 13084
rect 3550 13024 3614 13028
rect 3630 13084 3694 13088
rect 3630 13028 3634 13084
rect 3634 13028 3690 13084
rect 3690 13028 3694 13084
rect 3630 13024 3694 13028
rect 5828 13084 5892 13088
rect 5828 13028 5832 13084
rect 5832 13028 5888 13084
rect 5888 13028 5892 13084
rect 5828 13024 5892 13028
rect 5908 13084 5972 13088
rect 5908 13028 5912 13084
rect 5912 13028 5968 13084
rect 5968 13028 5972 13084
rect 5908 13024 5972 13028
rect 5988 13084 6052 13088
rect 5988 13028 5992 13084
rect 5992 13028 6048 13084
rect 6048 13028 6052 13084
rect 5988 13024 6052 13028
rect 6068 13084 6132 13088
rect 6068 13028 6072 13084
rect 6072 13028 6128 13084
rect 6128 13028 6132 13084
rect 6068 13024 6132 13028
rect 8266 13084 8330 13088
rect 8266 13028 8270 13084
rect 8270 13028 8326 13084
rect 8326 13028 8330 13084
rect 8266 13024 8330 13028
rect 8346 13084 8410 13088
rect 8346 13028 8350 13084
rect 8350 13028 8406 13084
rect 8406 13028 8410 13084
rect 8346 13024 8410 13028
rect 8426 13084 8490 13088
rect 8426 13028 8430 13084
rect 8430 13028 8486 13084
rect 8486 13028 8490 13084
rect 8426 13024 8490 13028
rect 8506 13084 8570 13088
rect 8506 13028 8510 13084
rect 8510 13028 8566 13084
rect 8566 13028 8570 13084
rect 8506 13024 8570 13028
rect 10704 13084 10768 13088
rect 10704 13028 10708 13084
rect 10708 13028 10764 13084
rect 10764 13028 10768 13084
rect 10704 13024 10768 13028
rect 10784 13084 10848 13088
rect 10784 13028 10788 13084
rect 10788 13028 10844 13084
rect 10844 13028 10848 13084
rect 10784 13024 10848 13028
rect 10864 13084 10928 13088
rect 10864 13028 10868 13084
rect 10868 13028 10924 13084
rect 10924 13028 10928 13084
rect 10864 13024 10928 13028
rect 10944 13084 11008 13088
rect 10944 13028 10948 13084
rect 10948 13028 11004 13084
rect 11004 13028 11008 13084
rect 10944 13024 11008 13028
rect 2171 12540 2235 12544
rect 2171 12484 2175 12540
rect 2175 12484 2231 12540
rect 2231 12484 2235 12540
rect 2171 12480 2235 12484
rect 2251 12540 2315 12544
rect 2251 12484 2255 12540
rect 2255 12484 2311 12540
rect 2311 12484 2315 12540
rect 2251 12480 2315 12484
rect 2331 12540 2395 12544
rect 2331 12484 2335 12540
rect 2335 12484 2391 12540
rect 2391 12484 2395 12540
rect 2331 12480 2395 12484
rect 2411 12540 2475 12544
rect 2411 12484 2415 12540
rect 2415 12484 2471 12540
rect 2471 12484 2475 12540
rect 2411 12480 2475 12484
rect 4609 12540 4673 12544
rect 4609 12484 4613 12540
rect 4613 12484 4669 12540
rect 4669 12484 4673 12540
rect 4609 12480 4673 12484
rect 4689 12540 4753 12544
rect 4689 12484 4693 12540
rect 4693 12484 4749 12540
rect 4749 12484 4753 12540
rect 4689 12480 4753 12484
rect 4769 12540 4833 12544
rect 4769 12484 4773 12540
rect 4773 12484 4829 12540
rect 4829 12484 4833 12540
rect 4769 12480 4833 12484
rect 4849 12540 4913 12544
rect 4849 12484 4853 12540
rect 4853 12484 4909 12540
rect 4909 12484 4913 12540
rect 4849 12480 4913 12484
rect 7047 12540 7111 12544
rect 7047 12484 7051 12540
rect 7051 12484 7107 12540
rect 7107 12484 7111 12540
rect 7047 12480 7111 12484
rect 7127 12540 7191 12544
rect 7127 12484 7131 12540
rect 7131 12484 7187 12540
rect 7187 12484 7191 12540
rect 7127 12480 7191 12484
rect 7207 12540 7271 12544
rect 7207 12484 7211 12540
rect 7211 12484 7267 12540
rect 7267 12484 7271 12540
rect 7207 12480 7271 12484
rect 7287 12540 7351 12544
rect 7287 12484 7291 12540
rect 7291 12484 7347 12540
rect 7347 12484 7351 12540
rect 7287 12480 7351 12484
rect 9485 12540 9549 12544
rect 9485 12484 9489 12540
rect 9489 12484 9545 12540
rect 9545 12484 9549 12540
rect 9485 12480 9549 12484
rect 9565 12540 9629 12544
rect 9565 12484 9569 12540
rect 9569 12484 9625 12540
rect 9625 12484 9629 12540
rect 9565 12480 9629 12484
rect 9645 12540 9709 12544
rect 9645 12484 9649 12540
rect 9649 12484 9705 12540
rect 9705 12484 9709 12540
rect 9645 12480 9709 12484
rect 9725 12540 9789 12544
rect 9725 12484 9729 12540
rect 9729 12484 9785 12540
rect 9785 12484 9789 12540
rect 9725 12480 9789 12484
rect 3390 11996 3454 12000
rect 3390 11940 3394 11996
rect 3394 11940 3450 11996
rect 3450 11940 3454 11996
rect 3390 11936 3454 11940
rect 3470 11996 3534 12000
rect 3470 11940 3474 11996
rect 3474 11940 3530 11996
rect 3530 11940 3534 11996
rect 3470 11936 3534 11940
rect 3550 11996 3614 12000
rect 3550 11940 3554 11996
rect 3554 11940 3610 11996
rect 3610 11940 3614 11996
rect 3550 11936 3614 11940
rect 3630 11996 3694 12000
rect 3630 11940 3634 11996
rect 3634 11940 3690 11996
rect 3690 11940 3694 11996
rect 3630 11936 3694 11940
rect 5828 11996 5892 12000
rect 5828 11940 5832 11996
rect 5832 11940 5888 11996
rect 5888 11940 5892 11996
rect 5828 11936 5892 11940
rect 5908 11996 5972 12000
rect 5908 11940 5912 11996
rect 5912 11940 5968 11996
rect 5968 11940 5972 11996
rect 5908 11936 5972 11940
rect 5988 11996 6052 12000
rect 5988 11940 5992 11996
rect 5992 11940 6048 11996
rect 6048 11940 6052 11996
rect 5988 11936 6052 11940
rect 6068 11996 6132 12000
rect 6068 11940 6072 11996
rect 6072 11940 6128 11996
rect 6128 11940 6132 11996
rect 6068 11936 6132 11940
rect 8266 11996 8330 12000
rect 8266 11940 8270 11996
rect 8270 11940 8326 11996
rect 8326 11940 8330 11996
rect 8266 11936 8330 11940
rect 8346 11996 8410 12000
rect 8346 11940 8350 11996
rect 8350 11940 8406 11996
rect 8406 11940 8410 11996
rect 8346 11936 8410 11940
rect 8426 11996 8490 12000
rect 8426 11940 8430 11996
rect 8430 11940 8486 11996
rect 8486 11940 8490 11996
rect 8426 11936 8490 11940
rect 8506 11996 8570 12000
rect 8506 11940 8510 11996
rect 8510 11940 8566 11996
rect 8566 11940 8570 11996
rect 8506 11936 8570 11940
rect 10704 11996 10768 12000
rect 10704 11940 10708 11996
rect 10708 11940 10764 11996
rect 10764 11940 10768 11996
rect 10704 11936 10768 11940
rect 10784 11996 10848 12000
rect 10784 11940 10788 11996
rect 10788 11940 10844 11996
rect 10844 11940 10848 11996
rect 10784 11936 10848 11940
rect 10864 11996 10928 12000
rect 10864 11940 10868 11996
rect 10868 11940 10924 11996
rect 10924 11940 10928 11996
rect 10864 11936 10928 11940
rect 10944 11996 11008 12000
rect 10944 11940 10948 11996
rect 10948 11940 11004 11996
rect 11004 11940 11008 11996
rect 10944 11936 11008 11940
rect 2171 11452 2235 11456
rect 2171 11396 2175 11452
rect 2175 11396 2231 11452
rect 2231 11396 2235 11452
rect 2171 11392 2235 11396
rect 2251 11452 2315 11456
rect 2251 11396 2255 11452
rect 2255 11396 2311 11452
rect 2311 11396 2315 11452
rect 2251 11392 2315 11396
rect 2331 11452 2395 11456
rect 2331 11396 2335 11452
rect 2335 11396 2391 11452
rect 2391 11396 2395 11452
rect 2331 11392 2395 11396
rect 2411 11452 2475 11456
rect 2411 11396 2415 11452
rect 2415 11396 2471 11452
rect 2471 11396 2475 11452
rect 2411 11392 2475 11396
rect 4609 11452 4673 11456
rect 4609 11396 4613 11452
rect 4613 11396 4669 11452
rect 4669 11396 4673 11452
rect 4609 11392 4673 11396
rect 4689 11452 4753 11456
rect 4689 11396 4693 11452
rect 4693 11396 4749 11452
rect 4749 11396 4753 11452
rect 4689 11392 4753 11396
rect 4769 11452 4833 11456
rect 4769 11396 4773 11452
rect 4773 11396 4829 11452
rect 4829 11396 4833 11452
rect 4769 11392 4833 11396
rect 4849 11452 4913 11456
rect 4849 11396 4853 11452
rect 4853 11396 4909 11452
rect 4909 11396 4913 11452
rect 4849 11392 4913 11396
rect 7047 11452 7111 11456
rect 7047 11396 7051 11452
rect 7051 11396 7107 11452
rect 7107 11396 7111 11452
rect 7047 11392 7111 11396
rect 7127 11452 7191 11456
rect 7127 11396 7131 11452
rect 7131 11396 7187 11452
rect 7187 11396 7191 11452
rect 7127 11392 7191 11396
rect 7207 11452 7271 11456
rect 7207 11396 7211 11452
rect 7211 11396 7267 11452
rect 7267 11396 7271 11452
rect 7207 11392 7271 11396
rect 7287 11452 7351 11456
rect 7287 11396 7291 11452
rect 7291 11396 7347 11452
rect 7347 11396 7351 11452
rect 7287 11392 7351 11396
rect 9485 11452 9549 11456
rect 9485 11396 9489 11452
rect 9489 11396 9545 11452
rect 9545 11396 9549 11452
rect 9485 11392 9549 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 3390 10908 3454 10912
rect 3390 10852 3394 10908
rect 3394 10852 3450 10908
rect 3450 10852 3454 10908
rect 3390 10848 3454 10852
rect 3470 10908 3534 10912
rect 3470 10852 3474 10908
rect 3474 10852 3530 10908
rect 3530 10852 3534 10908
rect 3470 10848 3534 10852
rect 3550 10908 3614 10912
rect 3550 10852 3554 10908
rect 3554 10852 3610 10908
rect 3610 10852 3614 10908
rect 3550 10848 3614 10852
rect 3630 10908 3694 10912
rect 3630 10852 3634 10908
rect 3634 10852 3690 10908
rect 3690 10852 3694 10908
rect 3630 10848 3694 10852
rect 5828 10908 5892 10912
rect 5828 10852 5832 10908
rect 5832 10852 5888 10908
rect 5888 10852 5892 10908
rect 5828 10848 5892 10852
rect 5908 10908 5972 10912
rect 5908 10852 5912 10908
rect 5912 10852 5968 10908
rect 5968 10852 5972 10908
rect 5908 10848 5972 10852
rect 5988 10908 6052 10912
rect 5988 10852 5992 10908
rect 5992 10852 6048 10908
rect 6048 10852 6052 10908
rect 5988 10848 6052 10852
rect 6068 10908 6132 10912
rect 6068 10852 6072 10908
rect 6072 10852 6128 10908
rect 6128 10852 6132 10908
rect 6068 10848 6132 10852
rect 8266 10908 8330 10912
rect 8266 10852 8270 10908
rect 8270 10852 8326 10908
rect 8326 10852 8330 10908
rect 8266 10848 8330 10852
rect 8346 10908 8410 10912
rect 8346 10852 8350 10908
rect 8350 10852 8406 10908
rect 8406 10852 8410 10908
rect 8346 10848 8410 10852
rect 8426 10908 8490 10912
rect 8426 10852 8430 10908
rect 8430 10852 8486 10908
rect 8486 10852 8490 10908
rect 8426 10848 8490 10852
rect 8506 10908 8570 10912
rect 8506 10852 8510 10908
rect 8510 10852 8566 10908
rect 8566 10852 8570 10908
rect 8506 10848 8570 10852
rect 10704 10908 10768 10912
rect 10704 10852 10708 10908
rect 10708 10852 10764 10908
rect 10764 10852 10768 10908
rect 10704 10848 10768 10852
rect 10784 10908 10848 10912
rect 10784 10852 10788 10908
rect 10788 10852 10844 10908
rect 10844 10852 10848 10908
rect 10784 10848 10848 10852
rect 10864 10908 10928 10912
rect 10864 10852 10868 10908
rect 10868 10852 10924 10908
rect 10924 10852 10928 10908
rect 10864 10848 10928 10852
rect 10944 10908 11008 10912
rect 10944 10852 10948 10908
rect 10948 10852 11004 10908
rect 11004 10852 11008 10908
rect 10944 10848 11008 10852
rect 2171 10364 2235 10368
rect 2171 10308 2175 10364
rect 2175 10308 2231 10364
rect 2231 10308 2235 10364
rect 2171 10304 2235 10308
rect 2251 10364 2315 10368
rect 2251 10308 2255 10364
rect 2255 10308 2311 10364
rect 2311 10308 2315 10364
rect 2251 10304 2315 10308
rect 2331 10364 2395 10368
rect 2331 10308 2335 10364
rect 2335 10308 2391 10364
rect 2391 10308 2395 10364
rect 2331 10304 2395 10308
rect 2411 10364 2475 10368
rect 2411 10308 2415 10364
rect 2415 10308 2471 10364
rect 2471 10308 2475 10364
rect 2411 10304 2475 10308
rect 4609 10364 4673 10368
rect 4609 10308 4613 10364
rect 4613 10308 4669 10364
rect 4669 10308 4673 10364
rect 4609 10304 4673 10308
rect 4689 10364 4753 10368
rect 4689 10308 4693 10364
rect 4693 10308 4749 10364
rect 4749 10308 4753 10364
rect 4689 10304 4753 10308
rect 4769 10364 4833 10368
rect 4769 10308 4773 10364
rect 4773 10308 4829 10364
rect 4829 10308 4833 10364
rect 4769 10304 4833 10308
rect 4849 10364 4913 10368
rect 4849 10308 4853 10364
rect 4853 10308 4909 10364
rect 4909 10308 4913 10364
rect 4849 10304 4913 10308
rect 7047 10364 7111 10368
rect 7047 10308 7051 10364
rect 7051 10308 7107 10364
rect 7107 10308 7111 10364
rect 7047 10304 7111 10308
rect 7127 10364 7191 10368
rect 7127 10308 7131 10364
rect 7131 10308 7187 10364
rect 7187 10308 7191 10364
rect 7127 10304 7191 10308
rect 7207 10364 7271 10368
rect 7207 10308 7211 10364
rect 7211 10308 7267 10364
rect 7267 10308 7271 10364
rect 7207 10304 7271 10308
rect 7287 10364 7351 10368
rect 7287 10308 7291 10364
rect 7291 10308 7347 10364
rect 7347 10308 7351 10364
rect 7287 10304 7351 10308
rect 9485 10364 9549 10368
rect 9485 10308 9489 10364
rect 9489 10308 9545 10364
rect 9545 10308 9549 10364
rect 9485 10304 9549 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 15808 2483 15824
rect 2163 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2483 15808
rect 2163 14720 2483 15744
rect 2163 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2483 14720
rect 2163 13632 2483 14656
rect 2163 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2483 13632
rect 2163 12544 2483 13568
rect 2163 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2483 12544
rect 2163 11456 2483 12480
rect 2163 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2483 11456
rect 2163 10368 2483 11392
rect 2163 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2483 10368
rect 2163 9280 2483 10304
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 15264 3702 15824
rect 3382 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3702 15264
rect 3382 14176 3702 15200
rect 3382 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3702 14176
rect 3382 13088 3702 14112
rect 3382 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3702 13088
rect 3382 12000 3702 13024
rect 3382 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3702 12000
rect 3382 10912 3702 11936
rect 3382 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3702 10912
rect 3382 9824 3702 10848
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 15808 4921 15824
rect 4601 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4921 15808
rect 4601 14720 4921 15744
rect 4601 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4921 14720
rect 4601 13632 4921 14656
rect 4601 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4921 13632
rect 4601 12544 4921 13568
rect 4601 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4921 12544
rect 4601 11456 4921 12480
rect 4601 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4921 11456
rect 4601 10368 4921 11392
rect 4601 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4921 10368
rect 4601 9280 4921 10304
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 15264 6140 15824
rect 5820 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6140 15264
rect 5820 14176 6140 15200
rect 5820 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6140 14176
rect 5820 13088 6140 14112
rect 5820 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6140 13088
rect 5820 12000 6140 13024
rect 5820 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6140 12000
rect 5820 10912 6140 11936
rect 5820 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6140 10912
rect 5820 9824 6140 10848
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 15808 7359 15824
rect 7039 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7359 15808
rect 7039 14720 7359 15744
rect 7039 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7359 14720
rect 7039 13632 7359 14656
rect 7039 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7359 13632
rect 7039 12544 7359 13568
rect 7039 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7359 12544
rect 7039 11456 7359 12480
rect 7039 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7359 11456
rect 7039 10368 7359 11392
rect 7039 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7359 10368
rect 7039 9280 7359 10304
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 15264 8578 15824
rect 8258 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8578 15264
rect 8258 14176 8578 15200
rect 8258 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8578 14176
rect 8258 13088 8578 14112
rect 8258 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8578 13088
rect 8258 12000 8578 13024
rect 8258 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8578 12000
rect 8258 10912 8578 11936
rect 8258 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8578 10912
rect 8258 9824 8578 10848
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 15808 9797 15824
rect 9477 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9797 15808
rect 9477 14720 9797 15744
rect 9477 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9797 14720
rect 9477 13632 9797 14656
rect 9477 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9797 13632
rect 9477 12544 9797 13568
rect 9477 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9797 12544
rect 9477 11456 9797 12480
rect 9477 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9797 11456
rect 9477 10368 9797 11392
rect 9477 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9797 10368
rect 9477 9280 9797 10304
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 15264 11016 15824
rect 10696 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11016 15264
rect 10696 14176 11016 15200
rect 10696 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11016 14176
rect 10696 13088 11016 14112
rect 10696 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11016 13088
rect 10696 12000 11016 13024
rect 10696 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11016 12000
rect 10696 10912 11016 11936
rect 10696 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11016 10912
rect 10696 9824 11016 10848
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform -1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101
timestamp 1676037725
transform 1 0 10396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp 1676037725
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_66
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1676037725
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_86
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1676037725
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_74
timestamp 1676037725
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1676037725
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_83
timestamp 1676037725
transform 1 0 8740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1676037725
transform 1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1676037725
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1676037725
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1676037725
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1676037725
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1676037725
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_60
timestamp 1676037725
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1676037725
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_64
timestamp 1676037725
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_77
timestamp 1676037725
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_89
timestamp 1676037725
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1676037725
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 1676037725
transform 1 0 5520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1676037725
transform 1 0 6900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1676037725
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1676037725
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1676037725
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1676037725
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1676037725
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_74
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_86
timestamp 1676037725
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1676037725
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1676037725
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1676037725
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_60
timestamp 1676037725
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 1676037725
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_62
timestamp 1676037725
transform 1 0 6808 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_74
timestamp 1676037725
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_86
timestamp 1676037725
transform 1 0 9016 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1676037725
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_19
timestamp 1676037725
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 1676037725
transform 1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_66
timestamp 1676037725
transform 1 0 7176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1676037725
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1676037725
transform 1 0 4600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_67
timestamp 1676037725
transform 1 0 7268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_79
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1676037725
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1676037725
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_77
timestamp 1676037725
transform 1 0 8188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_66
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1676037725
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1676037725
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1676037725
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_67
timestamp 1676037725
transform 1 0 7268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_79
timestamp 1676037725
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_91
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1676037725
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_50
timestamp 1676037725
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_57
timestamp 1676037725
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_69
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1676037725
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1676037725
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1676037725
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_72
timestamp 1676037725
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_84
timestamp 1676037725
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_96
timestamp 1676037725
transform 1 0 9936 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_102
timestamp 1676037725
transform 1 0 10488 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1676037725
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _33_
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _34_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _35_
timestamp 1676037725
transform 1 0 6164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _36__1
timestamp 1676037725
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _36__2
timestamp 1676037725
transform -1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp 1676037725
transform 1 0 4876 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _45_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _46_
timestamp 1676037725
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _47_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _48_
timestamp 1676037725
transform -1 0 6072 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _49_
timestamp 1676037725
transform -1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _50_
timestamp 1676037725
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _51_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _53_
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _54_
timestamp 1676037725
transform 1 0 6164 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _55_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6900 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _56_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _57_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _58_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _59_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _60_
timestamp 1676037725
transform -1 0 8556 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _61_
timestamp 1676037725
transform -1 0 7912 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _62_
timestamp 1676037725
transform -1 0 7728 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _63_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _64_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _65_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _66_
timestamp 1676037725
transform -1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _67_
timestamp 1676037725
transform -1 0 6900 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _68__3
timestamp 1676037725
transform -1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _69__4
timestamp 1676037725
transform -1 0 3496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _70__5
timestamp 1676037725
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _71_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _72_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _73_
timestamp 1676037725
transform 1 0 3496 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _74_
timestamp 1676037725
transform 1 0 3680 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _75_
timestamp 1676037725
transform 1 0 3772 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _76_
timestamp 1676037725
transform 1 0 3036 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _77_
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _78_
timestamp 1676037725
transform -1 0 5704 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _80_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform -1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform -1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform -1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1676037725
transform -1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform -1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1676037725
transform -1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1676037725
transform -1 0 3404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 4784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 5980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 6624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_MC14500_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10396 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 2962 17200 3018 18000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 11200 1776 12000 1896 0 FreeSans 480 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 11200 5312 12000 5432 0 FreeSans 480 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 11200 8848 12000 8968 0 FreeSans 480 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 11200 12384 12000 12504 0 FreeSans 480 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 11200 15920 12000 16040 0 FreeSans 480 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 io_oeb
port 6 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 io_out[8]
port 15 nsew signal tristate
flabel metal2 s 8942 17200 8998 18000 0 FreeSans 224 90 0 0 rst
port 16 nsew signal input
flabel metal4 s 2163 2128 2483 15824 0 FreeSans 1920 90 0 0 vccd1
port 17 nsew power bidirectional
flabel metal4 s 4601 2128 4921 15824 0 FreeSans 1920 90 0 0 vccd1
port 17 nsew power bidirectional
flabel metal4 s 7039 2128 7359 15824 0 FreeSans 1920 90 0 0 vccd1
port 17 nsew power bidirectional
flabel metal4 s 9477 2128 9797 15824 0 FreeSans 1920 90 0 0 vccd1
port 17 nsew power bidirectional
flabel metal4 s 3382 2128 3702 15824 0 FreeSans 1920 90 0 0 vssd1
port 18 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 15824 0 FreeSans 1920 90 0 0 vssd1
port 18 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 15824 0 FreeSans 1920 90 0 0 vssd1
port 18 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 15824 0 FreeSans 1920 90 0 0 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 18000
<< end >>
