magic
tech sky130B
magscale 1 2
timestamp 1682095495
<< nwell >>
rect 1066 18757 20922 19323
rect 1066 17669 20922 18235
rect 1066 16581 20922 17147
rect 1066 15493 20922 16059
rect 1066 14405 20922 14971
rect 1066 13317 20922 13883
rect 1066 12229 20922 12795
rect 1066 11141 20922 11707
rect 1066 10053 20922 10619
rect 1066 8965 20922 9531
rect 1066 7877 20922 8443
rect 1066 6789 20922 7355
rect 1066 5701 20922 6267
rect 1066 4613 20922 5179
rect 1066 3525 20922 4091
rect 1066 2437 20922 3003
<< obsli1 >>
rect 1104 2159 20884 19601
<< obsm1 >>
rect 1104 2128 21043 19712
<< metal2 >>
rect 3698 21200 3754 22000
rect 10966 21200 11022 22000
rect 18234 21200 18290 22000
rect 1582 0 1638 800
rect 4250 0 4306 800
rect 6918 0 6974 800
rect 9586 0 9642 800
rect 12254 0 12310 800
rect 14922 0 14978 800
rect 17590 0 17646 800
rect 20258 0 20314 800
<< obsm2 >>
rect 1584 21144 3642 21298
rect 3810 21144 10910 21298
rect 11078 21144 18178 21298
rect 18346 21144 21037 21298
rect 1584 856 21037 21144
rect 1694 800 4194 856
rect 4362 800 6862 856
rect 7030 800 9530 856
rect 9698 800 12198 856
rect 12366 800 14866 856
rect 15034 800 17534 856
rect 17702 800 20202 856
rect 20370 800 21037 856
<< obsm3 >>
rect 3418 2143 21041 19617
<< metal4 >>
rect 3416 2128 3736 19632
rect 5888 2128 6208 19632
rect 8361 2128 8681 19632
rect 10833 2128 11153 19632
rect 13306 2128 13626 19632
rect 15778 2128 16098 19632
rect 18251 2128 18571 19632
rect 20723 2128 21043 19632
<< labels >>
rlabel metal2 s 3698 21200 3754 22000 6 clk
port 1 nsew signal input
rlabel metal2 s 18234 21200 18290 22000 6 io_in
port 2 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 io_out[0]
port 3 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 io_out[1]
port 4 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 io_out[2]
port 5 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 io_out[3]
port 6 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 io_out[4]
port 7 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 io_out[5]
port 8 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 io_out[6]
port 9 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_out[7]
port 10 nsew signal output
rlabel metal2 s 10966 21200 11022 22000 6 rst
port 11 nsew signal input
rlabel metal4 s 3416 2128 3736 19632 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 8361 2128 8681 19632 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 13306 2128 13626 19632 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 18251 2128 18571 19632 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 5888 2128 6208 19632 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 10833 2128 11153 19632 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 15778 2128 16098 19632 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 20723 2128 21043 19632 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1256896
string GDS_FILE /run/media/tholin/Data/Projects/MPW/TMBoC/openlane/Diceroll/runs/23_04_21_18_43/results/signoff/tt2_tholin_diceroll.magic.gds
string GDS_START 488450
<< end >>

