magic
tech sky130B
magscale 1 2
timestamp 1683543228
<< obsli1 >>
rect 1104 2159 73876 72369
<< obsm1 >>
rect 842 2128 74138 74112
<< metal2 >>
rect 3514 74200 3570 75000
rect 9678 74200 9734 75000
rect 15842 74200 15898 75000
rect 22006 74200 22062 75000
rect 28170 74200 28226 75000
rect 34334 74200 34390 75000
rect 40498 74200 40554 75000
rect 46662 74200 46718 75000
rect 52826 74200 52882 75000
rect 58990 74200 59046 75000
rect 65154 74200 65210 75000
rect 71318 74200 71374 75000
<< obsm2 >>
rect 754 74144 3458 74338
rect 3626 74144 9622 74338
rect 9790 74144 15786 74338
rect 15954 74144 21950 74338
rect 22118 74144 28114 74338
rect 28282 74144 34278 74338
rect 34446 74144 40442 74338
rect 40610 74144 46606 74338
rect 46774 74144 52770 74338
rect 52938 74144 58934 74338
rect 59102 74144 65098 74338
rect 65266 74144 71262 74338
rect 71430 74144 74134 74338
rect 754 2139 74134 74144
<< metal3 >>
rect 74200 37408 75000 37528
<< obsm3 >>
rect 749 37608 74200 72385
rect 749 37328 74120 37608
rect 749 2143 74200 37328
<< metal4 >>
rect 4208 2128 4528 72400
rect 19568 2128 19888 72400
rect 34928 2128 35248 72400
rect 50288 2128 50608 72400
rect 65648 2128 65968 72400
<< obsm4 >>
rect 979 3979 4128 60077
rect 4608 3979 19488 60077
rect 19968 3979 34848 60077
rect 35328 3979 50208 60077
rect 50688 3979 65568 60077
rect 66048 3979 70229 60077
<< labels >>
rlabel metal2 s 3514 74200 3570 75000 6 clk
port 1 nsew signal input
rlabel metal3 s 74200 37408 75000 37528 6 io_in
port 2 nsew signal input
rlabel metal2 s 15842 74200 15898 75000 6 io_out[0]
port 3 nsew signal output
rlabel metal2 s 22006 74200 22062 75000 6 io_out[1]
port 4 nsew signal output
rlabel metal2 s 28170 74200 28226 75000 6 io_out[2]
port 5 nsew signal output
rlabel metal2 s 34334 74200 34390 75000 6 io_out[3]
port 6 nsew signal output
rlabel metal2 s 40498 74200 40554 75000 6 io_out[4]
port 7 nsew signal output
rlabel metal2 s 46662 74200 46718 75000 6 io_out[5]
port 8 nsew signal output
rlabel metal2 s 52826 74200 52882 75000 6 io_out[6]
port 9 nsew signal output
rlabel metal2 s 58990 74200 59046 75000 6 io_out[7]
port 10 nsew signal output
rlabel metal2 s 65154 74200 65210 75000 6 io_out[8]
port 11 nsew signal output
rlabel metal2 s 71318 74200 71374 75000 6 io_out[9]
port 12 nsew signal output
rlabel metal2 s 9678 74200 9734 75000 6 rst
port 13 nsew signal input
rlabel metal4 s 4208 2128 4528 72400 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 72400 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 72400 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 72400 6 vssd1
port 15 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 72400 6 vssd1
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 75000 75000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10906666
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/VGATest/runs/23_05_08_12_46/results/signoff/wrapped_vgatest.magic.gds
string GDS_START 1081210
<< end >>

