VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt2_tholin_multiplier
  CLASS BLOCK ;
  FOREIGN tt2_tholin_multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 90.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 79.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.910 10.640 18.510 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.100 10.640 30.700 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.290 10.640 42.890 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.480 10.640 55.080 79.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 78.965 ;
      LAYER met1 ;
        RECT 3.750 10.640 55.590 79.120 ;
      LAYER met2 ;
        RECT 3.780 4.280 55.560 82.805 ;
        RECT 4.330 4.000 10.850 4.280 ;
        RECT 11.690 4.000 18.210 4.280 ;
        RECT 19.050 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.930 4.280 ;
        RECT 33.770 4.000 40.290 4.280 ;
        RECT 41.130 4.000 47.650 4.280 ;
        RECT 48.490 4.000 55.010 4.280 ;
      LAYER met3 ;
        RECT 4.400 81.920 55.070 82.785 ;
        RECT 4.000 72.440 55.070 81.920 ;
        RECT 4.400 71.040 55.070 72.440 ;
        RECT 4.000 61.560 55.070 71.040 ;
        RECT 4.400 60.160 55.070 61.560 ;
        RECT 4.000 50.680 55.070 60.160 ;
        RECT 4.400 49.280 55.070 50.680 ;
        RECT 4.000 39.800 55.070 49.280 ;
        RECT 4.400 38.400 55.070 39.800 ;
        RECT 4.000 28.920 55.070 38.400 ;
        RECT 4.400 27.520 55.070 28.920 ;
        RECT 4.000 18.040 55.070 27.520 ;
        RECT 4.400 16.640 55.070 18.040 ;
        RECT 4.000 7.160 55.070 16.640 ;
        RECT 4.400 6.295 55.070 7.160 ;
  END
END tt2_tholin_multiplier
END LIBRARY

