// This is the unpowered netlist.
module tune_player (OP,
    clk,
    rst);
 output OP;
 input clk;
 input rst;

 wire \LFSR[0] ;
 wire \LFSR[1] ;
 wire \LFSR[2] ;
 wire \LFSR[3] ;
 wire \LFSR[4] ;
 wire \LFSR[5] ;
 wire \LFSR[6] ;
 wire OP_reg;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire \clock_div[0] ;
 wire \clock_div[1] ;
 wire \clock_div[2] ;
 wire \clock_div[3] ;
 wire \clock_div[4] ;
 wire \clock_div[5] ;
 wire \clock_div[6] ;
 wire \clock_div[7] ;
 wire \clock_div[8] ;
 wire just_inc;
 wire just_rst;
 wire prev_clk_div;
 wire \rhythm_LFSR[0] ;
 wire \rhythm_LFSR[1] ;
 wire \rhythm_LFSR[2] ;
 wire \rhythm_LFSR[3] ;
 wire \tempo_LFSR[0] ;
 wire \tempo_LFSR[1] ;
 wire \tempo_LFSR[2] ;
 wire \tempo_LFSR[3] ;
 wire \tune_ROM[0] ;
 wire \tune_ROM[1] ;
 wire \tune_ROM[2] ;
 wire \tune_ROM[3] ;
 wire \tune_ROM[4] ;
 wire \tune_ROM[5] ;
 wire net1;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _220_ (.A(\clock_div[7] ),
    .Y(_202_));
 sky130_fd_sc_hd__and4_1 _221_ (.A(\clock_div[0] ),
    .B(\clock_div[2] ),
    .C(\clock_div[3] ),
    .D(\clock_div[1] ),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_2 _222_ (.A(_203_),
    .X(_204_));
 sky130_fd_sc_hd__and2_1 _223_ (.A(\clock_div[4] ),
    .B(\clock_div[5] ),
    .X(_205_));
 sky130_fd_sc_hd__nand4_1 _224_ (.A(\clock_div[6] ),
    .B(\clock_div[8] ),
    .C(_204_),
    .D(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a41o_1 _225_ (.A1(\clock_div[6] ),
    .A2(\clock_div[7] ),
    .A3(_204_),
    .A4(_205_),
    .B1(\clock_div[8] ),
    .X(_207_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(prev_clk_div),
    .Y(_208_));
 sky130_fd_sc_hd__o211a_1 _227_ (.A1(_202_),
    .A2(_206_),
    .B1(_207_),
    .C1(_208_),
    .X(_209_));
 sky130_fd_sc_hd__clkinv_2 _228_ (.A(just_rst),
    .Y(_210_));
 sky130_fd_sc_hd__or2_1 _229_ (.A(\rhythm_LFSR[1] ),
    .B(\rhythm_LFSR[0] ),
    .X(_211_));
 sky130_fd_sc_hd__or3b_1 _230_ (.A(_211_),
    .B(\rhythm_LFSR[2] ),
    .C_N(\rhythm_LFSR[3] ),
    .X(_212_));
 sky130_fd_sc_hd__nand2_1 _231_ (.A(_210_),
    .B(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__or4b_1 _232_ (.A(\tempo_LFSR[2] ),
    .B(\tempo_LFSR[1] ),
    .C(\tempo_LFSR[0] ),
    .D_N(\tempo_LFSR[3] ),
    .X(_214_));
 sky130_fd_sc_hd__nand2_1 _233_ (.A(_210_),
    .B(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__o2111a_2 _234_ (.A1(just_rst),
    .A2(_209_),
    .B1(_213_),
    .C1(_215_),
    .D1(\PC[0] ),
    .X(_216_));
 sky130_fd_sc_hd__and4_1 _235_ (.A(\PC[3] ),
    .B(\PC[2] ),
    .C(\PC[1] ),
    .D(_216_),
    .X(_217_));
 sky130_fd_sc_hd__a21oi_1 _236_ (.A1(\PC[4] ),
    .A2(_217_),
    .B1(\PC[5] ),
    .Y(_218_));
 sky130_fd_sc_hd__a31o_1 _237_ (.A1(\PC[5] ),
    .A2(\PC[4] ),
    .A3(_217_),
    .B1(net1),
    .X(_219_));
 sky130_fd_sc_hd__or2_1 _238_ (.A(_218_),
    .B(_219_),
    .X(_039_));
 sky130_fd_sc_hd__buf_2 _239_ (.A(_039_),
    .X(_040_));
 sky130_fd_sc_hd__clkbuf_4 _240_ (.A(net1),
    .X(_041_));
 sky130_fd_sc_hd__xnor2_1 _241_ (.A(\PC[4] ),
    .B(_217_),
    .Y(_042_));
 sky130_fd_sc_hd__or2_2 _242_ (.A(_041_),
    .B(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__buf_2 _244_ (.A(_044_),
    .X(_014_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(_212_),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(_214_),
    .Y(_046_));
 sky130_fd_sc_hd__a311o_1 _247_ (.A1(_209_),
    .A2(_045_),
    .A3(_046_),
    .B1(just_rst),
    .C1(\PC[0] ),
    .X(_047_));
 sky130_fd_sc_hd__nor3b_4 _248_ (.A(net1),
    .B(_216_),
    .C_N(_047_),
    .Y(_010_));
 sky130_fd_sc_hd__and2_1 _249_ (.A(\PC[1] ),
    .B(_010_),
    .X(_048_));
 sky130_fd_sc_hd__and3_1 _250_ (.A(\PC[2] ),
    .B(\PC[1] ),
    .C(_216_),
    .X(_049_));
 sky130_fd_sc_hd__a21oi_1 _251_ (.A1(\PC[1] ),
    .A2(_216_),
    .B1(\PC[2] ),
    .Y(_050_));
 sky130_fd_sc_hd__or2_2 _252_ (.A(_049_),
    .B(_050_),
    .X(_051_));
 sky130_fd_sc_hd__a31o_1 _253_ (.A1(\PC[2] ),
    .A2(\PC[1] ),
    .A3(_216_),
    .B1(\PC[3] ),
    .X(_052_));
 sky130_fd_sc_hd__or3b_1 _254_ (.A(net1),
    .B(_217_),
    .C_N(_052_),
    .X(_053_));
 sky130_fd_sc_hd__buf_2 _255_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__a21o_1 _256_ (.A1(_048_),
    .A2(_051_),
    .B1(_054_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _257_ (.A(\PC[1] ),
    .B(_216_),
    .Y(_056_));
 sky130_fd_sc_hd__or2_2 _258_ (.A(net1),
    .B(_056_),
    .X(_057_));
 sky130_fd_sc_hd__or3_1 _259_ (.A(net1),
    .B(_049_),
    .C(_050_),
    .X(_058_));
 sky130_fd_sc_hd__clkbuf_2 _260_ (.A(_058_),
    .X(_059_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(_059_),
    .Y(_012_));
 sky130_fd_sc_hd__and3b_1 _262_ (.A_N(_055_),
    .B(_057_),
    .C(_012_),
    .X(_060_));
 sky130_fd_sc_hd__and2b_1 _263_ (.A_N(_216_),
    .B(_047_),
    .X(_061_));
 sky130_fd_sc_hd__or4_2 _264_ (.A(net1),
    .B(_061_),
    .C(_049_),
    .D(_050_),
    .X(_062_));
 sky130_fd_sc_hd__or2_2 _265_ (.A(_057_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__nand2_1 _266_ (.A(_048_),
    .B(_051_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(_054_),
    .Y(_065_));
 sky130_fd_sc_hd__buf_2 _268_ (.A(_065_),
    .X(_013_));
 sky130_fd_sc_hd__a21oi_1 _269_ (.A1(_063_),
    .A2(_064_),
    .B1(_013_),
    .Y(_066_));
 sky130_fd_sc_hd__or3_1 _270_ (.A(_014_),
    .B(_060_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__clkinv_2 _271_ (.A(_057_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _272_ (.A(_051_),
    .B(_013_),
    .Y(_068_));
 sky130_fd_sc_hd__o31ai_1 _273_ (.A1(_011_),
    .A2(_010_),
    .A3(_068_),
    .B1(_014_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _274_ (.A(\PC[2] ),
    .B(_057_),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _275_ (.A(\PC[1] ),
    .Y(_071_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(_071_),
    .B(_010_),
    .X(_072_));
 sky130_fd_sc_hd__nor2_1 _277_ (.A(_070_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(\PC[1] ),
    .B(_010_),
    .Y(_074_));
 sky130_fd_sc_hd__and3_1 _279_ (.A(_074_),
    .B(_051_),
    .C(_065_),
    .X(_075_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(_040_),
    .Y(_015_));
 sky130_fd_sc_hd__or3_1 _281_ (.A(\PC[2] ),
    .B(_041_),
    .C(_056_),
    .X(_076_));
 sky130_fd_sc_hd__o21ai_1 _282_ (.A1(_048_),
    .A2(_059_),
    .B1(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a221o_1 _283_ (.A1(\PC[2] ),
    .A2(_072_),
    .B1(_013_),
    .B2(_077_),
    .C1(_043_),
    .X(_078_));
 sky130_fd_sc_hd__o311a_1 _284_ (.A1(_073_),
    .A2(_014_),
    .A3(_075_),
    .B1(_015_),
    .C1(_078_),
    .X(_079_));
 sky130_fd_sc_hd__a31o_1 _285_ (.A1(_040_),
    .A2(_067_),
    .A3(_069_),
    .B1(_079_),
    .X(_000_));
 sky130_fd_sc_hd__nor3_1 _286_ (.A(\PC[4] ),
    .B(_054_),
    .C(_064_),
    .Y(_080_));
 sky130_fd_sc_hd__o2111a_1 _287_ (.A1(\PC[2] ),
    .A2(_013_),
    .B1(_071_),
    .C1(\PC[4] ),
    .D1(_010_),
    .X(_081_));
 sky130_fd_sc_hd__nand2_1 _288_ (.A(_051_),
    .B(_065_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(_048_),
    .A1(_072_),
    .S(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_1 _290_ (.A(_011_),
    .B(_062_),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(\PC[2] ),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _292_ (.A(_085_),
    .B(_074_),
    .Y(_086_));
 sky130_fd_sc_hd__or2b_1 _293_ (.A(_217_),
    .B_N(_052_),
    .X(_087_));
 sky130_fd_sc_hd__o221a_1 _294_ (.A1(_013_),
    .A2(_084_),
    .B1(_086_),
    .B2(_087_),
    .C1(_044_),
    .X(_088_));
 sky130_fd_sc_hd__a211o_1 _295_ (.A1(_043_),
    .A2(_083_),
    .B1(_088_),
    .C1(_040_),
    .X(_089_));
 sky130_fd_sc_hd__o31a_1 _296_ (.A1(_015_),
    .A2(_080_),
    .A3(_081_),
    .B1(_089_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_1 _297_ (.A(\PC[2] ),
    .B(_011_),
    .Y(_090_));
 sky130_fd_sc_hd__a21oi_1 _298_ (.A1(_010_),
    .A2(_090_),
    .B1(_075_),
    .Y(_091_));
 sky130_fd_sc_hd__and3_1 _299_ (.A(_072_),
    .B(_051_),
    .C(_065_),
    .X(_092_));
 sky130_fd_sc_hd__a211o_1 _300_ (.A1(_063_),
    .A2(_091_),
    .B1(_092_),
    .C1(_040_),
    .X(_093_));
 sky130_fd_sc_hd__nor2_1 _301_ (.A(_013_),
    .B(_084_),
    .Y(_094_));
 sky130_fd_sc_hd__or3_1 _302_ (.A(_041_),
    .B(_056_),
    .C(_061_),
    .X(_095_));
 sky130_fd_sc_hd__nand2_1 _303_ (.A(_059_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__nand2_1 _304_ (.A(_063_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__a221o_1 _305_ (.A1(_074_),
    .A2(_094_),
    .B1(_097_),
    .B2(_013_),
    .C1(_015_),
    .X(_098_));
 sky130_fd_sc_hd__o2bb2a_1 _306_ (.A1_N(_059_),
    .A2_N(_095_),
    .B1(_085_),
    .B2(_057_),
    .X(_099_));
 sky130_fd_sc_hd__a21oi_1 _307_ (.A1(_076_),
    .A2(_062_),
    .B1(_054_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_1 _308_ (.A1(_054_),
    .A2(_099_),
    .B1(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__a2111o_1 _309_ (.A1(_057_),
    .A2(_059_),
    .B1(_015_),
    .C1(_054_),
    .D1(_048_),
    .X(_102_));
 sky130_fd_sc_hd__o211a_1 _310_ (.A1(_040_),
    .A2(_101_),
    .B1(_102_),
    .C1(_043_),
    .X(_103_));
 sky130_fd_sc_hd__a31o_1 _311_ (.A1(_014_),
    .A2(_093_),
    .A3(_098_),
    .B1(_103_),
    .X(_002_));
 sky130_fd_sc_hd__a31o_1 _312_ (.A1(_076_),
    .A2(_065_),
    .A3(_063_),
    .B1(_015_),
    .X(_104_));
 sky130_fd_sc_hd__o211a_1 _313_ (.A1(_011_),
    .A2(_010_),
    .B1(_054_),
    .C1(_062_),
    .X(_105_));
 sky130_fd_sc_hd__and2b_1 _314_ (.A_N(_072_),
    .B(_059_),
    .X(_106_));
 sky130_fd_sc_hd__o31a_1 _315_ (.A1(_054_),
    .A2(_099_),
    .A3(_106_),
    .B1(_015_),
    .X(_107_));
 sky130_fd_sc_hd__o21ai_1 _316_ (.A1(_054_),
    .A2(_099_),
    .B1(_106_),
    .Y(_108_));
 sky130_fd_sc_hd__a2bb2o_1 _317_ (.A1_N(_104_),
    .A2_N(_105_),
    .B1(_107_),
    .B2(_108_),
    .X(_109_));
 sky130_fd_sc_hd__or3b_1 _318_ (.A(_092_),
    .B(_040_),
    .C_N(_095_),
    .X(_110_));
 sky130_fd_sc_hd__nor2_1 _319_ (.A(_013_),
    .B(_106_),
    .Y(_111_));
 sky130_fd_sc_hd__o41a_1 _320_ (.A1(_070_),
    .A2(_015_),
    .A3(_086_),
    .A4(_111_),
    .B1(_043_),
    .X(_112_));
 sky130_fd_sc_hd__a22o_1 _321_ (.A1(_014_),
    .A2(_109_),
    .B1(_110_),
    .B2(_112_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(\PC[3] ),
    .A1(_055_),
    .S(_063_),
    .X(_113_));
 sky130_fd_sc_hd__o21ai_1 _323_ (.A1(_074_),
    .A2(_082_),
    .B1(_014_),
    .Y(_114_));
 sky130_fd_sc_hd__o22a_1 _324_ (.A1(_014_),
    .A2(_113_),
    .B1(_114_),
    .B2(_084_),
    .X(_115_));
 sky130_fd_sc_hd__o22a_1 _325_ (.A1(_011_),
    .A2(_010_),
    .B1(_048_),
    .B2(_059_),
    .X(_116_));
 sky130_fd_sc_hd__a21oi_1 _326_ (.A1(_014_),
    .A2(_116_),
    .B1(_015_),
    .Y(_117_));
 sky130_fd_sc_hd__a211o_1 _327_ (.A1(_014_),
    .A2(_082_),
    .B1(_111_),
    .C1(_116_),
    .X(_118_));
 sky130_fd_sc_hd__a2bb2o_1 _328_ (.A1_N(_040_),
    .A2_N(_115_),
    .B1(_117_),
    .B2(_118_),
    .X(_004_));
 sky130_fd_sc_hd__a2bb2o_1 _329_ (.A1_N(\PC[4] ),
    .A2_N(_116_),
    .B1(_044_),
    .B2(_056_),
    .X(_119_));
 sky130_fd_sc_hd__nand2_1 _330_ (.A(_013_),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__o211a_1 _331_ (.A1(\PC[3] ),
    .A2(_063_),
    .B1(_055_),
    .C1(_042_),
    .X(_121_));
 sky130_fd_sc_hd__o2bb2a_1 _332_ (.A1_N(_117_),
    .A2_N(_120_),
    .B1(_121_),
    .B2(_040_),
    .X(_005_));
 sky130_fd_sc_hd__and2_1 _333_ (.A(OP_reg),
    .B(just_inc),
    .X(_122_));
 sky130_fd_sc_hd__buf_2 _334_ (.A(_122_),
    .X(OP));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(\tune_ROM[1] ),
    .B(_213_),
    .Y(_123_));
 sky130_fd_sc_hd__o21a_1 _336_ (.A1(\rhythm_LFSR[1] ),
    .A2(_213_),
    .B1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__nor2_1 _337_ (.A(just_rst),
    .B(_209_),
    .Y(_125_));
 sky130_fd_sc_hd__nor2_2 _338_ (.A(_041_),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__mux2_1 _339_ (.A0(\rhythm_LFSR[0] ),
    .A1(_124_),
    .S(_126_),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _340_ (.A(_127_),
    .X(_006_));
 sky130_fd_sc_hd__nand2_1 _341_ (.A(\tune_ROM[0] ),
    .B(\tune_ROM[1] ),
    .Y(_128_));
 sky130_fd_sc_hd__or2_1 _342_ (.A(\tune_ROM[0] ),
    .B(\tune_ROM[1] ),
    .X(_129_));
 sky130_fd_sc_hd__a32o_1 _343_ (.A1(_213_),
    .A2(_128_),
    .A3(_129_),
    .B1(\rhythm_LFSR[2] ),
    .B2(_210_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _344_ (.A0(\rhythm_LFSR[1] ),
    .A1(_130_),
    .S(_126_),
    .X(_131_));
 sky130_fd_sc_hd__clkbuf_1 _345_ (.A(_131_),
    .X(_007_));
 sky130_fd_sc_hd__nor2_1 _346_ (.A(just_rst),
    .B(_045_),
    .Y(_132_));
 sky130_fd_sc_hd__o22a_1 _347_ (.A1(just_rst),
    .A2(\rhythm_LFSR[3] ),
    .B1(\tune_ROM[0] ),
    .B2(_132_),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _348_ (.A0(\rhythm_LFSR[2] ),
    .A1(_133_),
    .S(_126_),
    .X(_134_));
 sky130_fd_sc_hd__clkbuf_1 _349_ (.A(_134_),
    .X(_008_));
 sky130_fd_sc_hd__a21oi_1 _350_ (.A1(\rhythm_LFSR[1] ),
    .A2(\rhythm_LFSR[0] ),
    .B1(just_rst),
    .Y(_135_));
 sky130_fd_sc_hd__a2bb2o_1 _351_ (.A1_N(\tune_ROM[0] ),
    .A2_N(_123_),
    .B1(_135_),
    .B2(_211_),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\rhythm_LFSR[3] ),
    .A1(_136_),
    .S(_126_),
    .X(_137_));
 sky130_fd_sc_hd__clkbuf_1 _353_ (.A(_137_),
    .X(_009_));
 sky130_fd_sc_hd__clkbuf_4 _354_ (.A(_041_),
    .X(_138_));
 sky130_fd_sc_hd__a31o_1 _355_ (.A1(_209_),
    .A2(_045_),
    .A3(_046_),
    .B1(just_rst),
    .X(_139_));
 sky130_fd_sc_hd__o21ba_1 _356_ (.A1(_125_),
    .A2(_132_),
    .B1_N(just_inc),
    .X(_140_));
 sky130_fd_sc_hd__nor3_1 _357_ (.A(_138_),
    .B(_139_),
    .C(_140_),
    .Y(_016_));
 sky130_fd_sc_hd__or2_1 _358_ (.A(\LFSR[1] ),
    .B(\LFSR[0] ),
    .X(_141_));
 sky130_fd_sc_hd__or4b_1 _359_ (.A(\LFSR[3] ),
    .B(_141_),
    .C(\LFSR[2] ),
    .D_N(\LFSR[6] ),
    .X(_142_));
 sky130_fd_sc_hd__o31ai_4 _360_ (.A1(\LFSR[5] ),
    .A2(\LFSR[4] ),
    .A3(_142_),
    .B1(_210_),
    .Y(_143_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(_041_),
    .Y(_144_));
 sky130_fd_sc_hd__o21ai_1 _362_ (.A1(OP_reg),
    .A2(_143_),
    .B1(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _363_ (.A1(OP_reg),
    .A2(_143_),
    .B1(_145_),
    .Y(_017_));
 sky130_fd_sc_hd__clkbuf_2 _364_ (.A(\tune_ROM[5] ),
    .X(_146_));
 sky130_fd_sc_hd__nor2_1 _365_ (.A(\tune_ROM[2] ),
    .B(\tune_ROM[3] ),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_1 _366_ (.A1(_146_),
    .A2(_147_),
    .B1(\tune_ROM[4] ),
    .Y(_148_));
 sky130_fd_sc_hd__nand2_1 _367_ (.A(\tune_ROM[2] ),
    .B(\tune_ROM[3] ),
    .Y(_149_));
 sky130_fd_sc_hd__or2_1 _368_ (.A(\tune_ROM[4] ),
    .B(\tune_ROM[3] ),
    .X(_150_));
 sky130_fd_sc_hd__nand3_1 _369_ (.A(_148_),
    .B(_149_),
    .C(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(\LFSR[1] ),
    .A1(_151_),
    .S(_143_),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(\LFSR[0] ),
    .A1(_152_),
    .S(_144_),
    .X(_153_));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(_153_),
    .X(_018_));
 sky130_fd_sc_hd__nor2_1 _373_ (.A(\tune_ROM[4] ),
    .B(_147_),
    .Y(_154_));
 sky130_fd_sc_hd__and2_1 _374_ (.A(\tune_ROM[4] ),
    .B(_147_),
    .X(_155_));
 sky130_fd_sc_hd__o21ai_1 _375_ (.A1(_154_),
    .A2(_155_),
    .B1(_146_),
    .Y(_156_));
 sky130_fd_sc_hd__or2_1 _376_ (.A(_146_),
    .B(_149_),
    .X(_157_));
 sky130_fd_sc_hd__a32o_1 _377_ (.A1(_143_),
    .A2(_156_),
    .A3(_157_),
    .B1(\LFSR[2] ),
    .B2(_210_),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\LFSR[1] ),
    .A1(_158_),
    .S(_144_),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_159_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(\tune_ROM[4] ),
    .B(\tune_ROM[3] ),
    .Y(_160_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(\tune_ROM[4] ),
    .Y(_161_));
 sky130_fd_sc_hd__o21ai_1 _382_ (.A1(_161_),
    .A2(_146_),
    .B1(\tune_ROM[2] ),
    .Y(_162_));
 sky130_fd_sc_hd__o211ai_1 _383_ (.A1(_146_),
    .A2(_150_),
    .B1(_160_),
    .C1(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(\LFSR[3] ),
    .A1(_163_),
    .S(_143_),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(\LFSR[2] ),
    .A1(_164_),
    .S(_144_),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_1 _386_ (.A(_165_),
    .X(_020_));
 sky130_fd_sc_hd__or2_1 _387_ (.A(\tune_ROM[4] ),
    .B(_149_),
    .X(_166_));
 sky130_fd_sc_hd__nand2_1 _388_ (.A(\tune_ROM[4] ),
    .B(_149_),
    .Y(_167_));
 sky130_fd_sc_hd__a22o_1 _389_ (.A1(_146_),
    .A2(_149_),
    .B1(_166_),
    .B2(_167_),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(\LFSR[4] ),
    .A1(_168_),
    .S(_143_),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\LFSR[3] ),
    .A1(_169_),
    .S(_144_),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_1 _392_ (.A(_170_),
    .X(_021_));
 sky130_fd_sc_hd__a21bo_1 _393_ (.A1(_161_),
    .A2(\tune_ROM[2] ),
    .B1_N(\tune_ROM[5] ),
    .X(_171_));
 sky130_fd_sc_hd__a211o_1 _394_ (.A1(_150_),
    .A2(_167_),
    .B1(_155_),
    .C1(_146_),
    .X(_172_));
 sky130_fd_sc_hd__o21ai_1 _395_ (.A1(_155_),
    .A2(_171_),
    .B1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(\LFSR[5] ),
    .A1(_173_),
    .S(_143_),
    .X(_174_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(\LFSR[4] ),
    .A1(_174_),
    .S(_144_),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _398_ (.A(_175_),
    .X(_022_));
 sky130_fd_sc_hd__and4bb_1 _399_ (.A_N(_146_),
    .B_N(_147_),
    .C(_150_),
    .D(_160_),
    .X(_176_));
 sky130_fd_sc_hd__a31o_1 _400_ (.A1(_146_),
    .A2(_149_),
    .A3(_154_),
    .B1(_176_),
    .X(_177_));
 sky130_fd_sc_hd__nand2_1 _401_ (.A(_143_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__o21a_1 _402_ (.A1(just_rst),
    .A2(\LFSR[6] ),
    .B1(_144_),
    .X(_179_));
 sky130_fd_sc_hd__a22o_1 _403_ (.A1(_138_),
    .A2(\LFSR[5] ),
    .B1(_178_),
    .B2(_179_),
    .X(_023_));
 sky130_fd_sc_hd__nand3b_1 _404_ (.A_N(_146_),
    .B(_166_),
    .C(_167_),
    .Y(_180_));
 sky130_fd_sc_hd__nand2_1 _405_ (.A(\LFSR[1] ),
    .B(\LFSR[0] ),
    .Y(_181_));
 sky130_fd_sc_hd__a21oi_1 _406_ (.A1(_141_),
    .A2(_181_),
    .B1(_143_),
    .Y(_182_));
 sky130_fd_sc_hd__a311o_1 _407_ (.A1(_143_),
    .A2(_171_),
    .A3(_180_),
    .B1(_182_),
    .C1(_041_),
    .X(_183_));
 sky130_fd_sc_hd__a21bo_1 _408_ (.A1(_138_),
    .A2(\LFSR[6] ),
    .B1_N(_183_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(\clock_div[8] ),
    .A1(prev_clk_div),
    .S(_041_),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _410_ (.A(_184_),
    .X(_025_));
 sky130_fd_sc_hd__nor2_1 _411_ (.A(\clock_div[0] ),
    .B(_138_),
    .Y(_026_));
 sky130_fd_sc_hd__a21oi_1 _412_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(_138_),
    .Y(_185_));
 sky130_fd_sc_hd__o21a_1 _413_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(_185_),
    .X(_027_));
 sky130_fd_sc_hd__and3_1 _414_ (.A(\clock_div[0] ),
    .B(\clock_div[2] ),
    .C(\clock_div[1] ),
    .X(_186_));
 sky130_fd_sc_hd__a21oi_1 _415_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(\clock_div[2] ),
    .Y(_187_));
 sky130_fd_sc_hd__nor3_1 _416_ (.A(_138_),
    .B(_186_),
    .C(_187_),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_1 _417_ (.A(_138_),
    .B(_204_),
    .Y(_188_));
 sky130_fd_sc_hd__o21a_1 _418_ (.A1(\clock_div[3] ),
    .A2(_186_),
    .B1(_188_),
    .X(_029_));
 sky130_fd_sc_hd__a21oi_1 _419_ (.A1(\clock_div[4] ),
    .A2(_204_),
    .B1(_138_),
    .Y(_189_));
 sky130_fd_sc_hd__o21a_1 _420_ (.A1(\clock_div[4] ),
    .A2(_204_),
    .B1(_189_),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _421_ (.A(_204_),
    .B(_205_),
    .X(_190_));
 sky130_fd_sc_hd__a21oi_1 _422_ (.A1(\clock_div[4] ),
    .A2(_204_),
    .B1(\clock_div[5] ),
    .Y(_191_));
 sky130_fd_sc_hd__nor3_1 _423_ (.A(_138_),
    .B(_190_),
    .C(_191_),
    .Y(_031_));
 sky130_fd_sc_hd__and3_1 _424_ (.A(\clock_div[6] ),
    .B(_204_),
    .C(_205_),
    .X(_192_));
 sky130_fd_sc_hd__nor2_1 _425_ (.A(_138_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__o21a_1 _426_ (.A1(\clock_div[6] ),
    .A2(_190_),
    .B1(_193_),
    .X(_032_));
 sky130_fd_sc_hd__a21o_1 _427_ (.A1(\clock_div[7] ),
    .A2(_192_),
    .B1(_041_),
    .X(_194_));
 sky130_fd_sc_hd__o21ba_1 _428_ (.A1(\clock_div[7] ),
    .A2(_192_),
    .B1_N(_194_),
    .X(_033_));
 sky130_fd_sc_hd__o211a_1 _429_ (.A1(_202_),
    .A2(_206_),
    .B1(_207_),
    .C1(_144_),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _430_ (.A(_213_),
    .B(_126_),
    .X(_195_));
 sky130_fd_sc_hd__or4_2 _431_ (.A(_041_),
    .B(_125_),
    .C(_132_),
    .D(_215_),
    .X(_196_));
 sky130_fd_sc_hd__o22a_1 _432_ (.A1(\tempo_LFSR[0] ),
    .A2(_195_),
    .B1(_196_),
    .B2(\tempo_LFSR[1] ),
    .X(_035_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(\tempo_LFSR[2] ),
    .Y(_197_));
 sky130_fd_sc_hd__nor2_1 _434_ (.A(_197_),
    .B(just_rst),
    .Y(_198_));
 sky130_fd_sc_hd__mux2_1 _435_ (.A0(\tempo_LFSR[1] ),
    .A1(_198_),
    .S(_195_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _436_ (.A(_199_),
    .X(_036_));
 sky130_fd_sc_hd__clkinv_2 _437_ (.A(_196_),
    .Y(_200_));
 sky130_fd_sc_hd__a2bb2o_1 _438_ (.A1_N(_197_),
    .A2_N(_195_),
    .B1(_200_),
    .B2(\tempo_LFSR[3] ),
    .X(_037_));
 sky130_fd_sc_hd__xor2_1 _439_ (.A(\tempo_LFSR[1] ),
    .B(\tempo_LFSR[0] ),
    .X(_201_));
 sky130_fd_sc_hd__o22a_1 _440_ (.A1(\tempo_LFSR[3] ),
    .A2(_195_),
    .B1(_196_),
    .B2(_201_),
    .X(_038_));
 sky130_fd_sc_hd__dfxtp_1 _441_ (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .Q(\tune_ROM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _442_ (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .Q(\tune_ROM[1] ));
 sky130_fd_sc_hd__dfxtp_1 _443_ (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .Q(\tune_ROM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _444_ (.CLK(clknet_2_2__leaf_clk),
    .D(_003_),
    .Q(\tune_ROM[3] ));
 sky130_fd_sc_hd__dfxtp_2 _445_ (.CLK(clknet_2_2__leaf_clk),
    .D(_004_),
    .Q(\tune_ROM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _446_ (.CLK(clknet_2_2__leaf_clk),
    .D(_005_),
    .Q(\tune_ROM[5] ));
 sky130_fd_sc_hd__dfxtp_1 _447_ (.CLK(clknet_2_3__leaf_clk),
    .D(_006_),
    .Q(\rhythm_LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _448_ (.CLK(clknet_2_3__leaf_clk),
    .D(_007_),
    .Q(\rhythm_LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _449_ (.CLK(clknet_2_3__leaf_clk),
    .D(_008_),
    .Q(\rhythm_LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _450_ (.CLK(clknet_2_3__leaf_clk),
    .D(_009_),
    .Q(\rhythm_LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _451_ (.CLK(clknet_2_3__leaf_clk),
    .D(_010_),
    .Q(\PC[0] ));
 sky130_fd_sc_hd__dfxtp_2 _452_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .Q(\PC[1] ));
 sky130_fd_sc_hd__dfxtp_2 _453_ (.CLK(clknet_2_2__leaf_clk),
    .D(_012_),
    .Q(\PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _454_ (.CLK(clknet_2_2__leaf_clk),
    .D(_013_),
    .Q(\PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _455_ (.CLK(clknet_2_2__leaf_clk),
    .D(_014_),
    .Q(\PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _456_ (.CLK(clknet_2_2__leaf_clk),
    .D(_015_),
    .Q(\PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _457_ (.CLK(clknet_2_3__leaf_clk),
    .D(_016_),
    .Q(just_inc));
 sky130_fd_sc_hd__dfxtp_1 _458_ (.CLK(clknet_2_1__leaf_clk),
    .D(_017_),
    .Q(OP_reg));
 sky130_fd_sc_hd__dfxtp_1 _459_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .Q(\LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _460_ (.CLK(clknet_2_1__leaf_clk),
    .D(_019_),
    .Q(\LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _461_ (.CLK(clknet_2_1__leaf_clk),
    .D(_020_),
    .Q(\LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _462_ (.CLK(clknet_2_1__leaf_clk),
    .D(_021_),
    .Q(\LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _463_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .Q(\LFSR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _464_ (.CLK(clknet_2_1__leaf_clk),
    .D(_023_),
    .Q(\LFSR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _465_ (.CLK(clknet_2_1__leaf_clk),
    .D(_024_),
    .Q(\LFSR[6] ));
 sky130_fd_sc_hd__dfxtp_1 _466_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .Q(prev_clk_div));
 sky130_fd_sc_hd__dfxtp_1 _467_ (.CLK(clknet_2_2__leaf_clk),
    .D(_026_),
    .Q(\clock_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _468_ (.CLK(clknet_2_2__leaf_clk),
    .D(_027_),
    .Q(\clock_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _469_ (.CLK(clknet_2_2__leaf_clk),
    .D(_028_),
    .Q(\clock_div[2] ));
 sky130_fd_sc_hd__dfxtp_1 _470_ (.CLK(clknet_2_0__leaf_clk),
    .D(_029_),
    .Q(\clock_div[3] ));
 sky130_fd_sc_hd__dfxtp_1 _471_ (.CLK(clknet_2_0__leaf_clk),
    .D(_030_),
    .Q(\clock_div[4] ));
 sky130_fd_sc_hd__dfxtp_1 _472_ (.CLK(clknet_2_0__leaf_clk),
    .D(_031_),
    .Q(\clock_div[5] ));
 sky130_fd_sc_hd__dfxtp_1 _473_ (.CLK(clknet_2_0__leaf_clk),
    .D(_032_),
    .Q(\clock_div[6] ));
 sky130_fd_sc_hd__dfxtp_1 _474_ (.CLK(clknet_2_0__leaf_clk),
    .D(_033_),
    .Q(\clock_div[7] ));
 sky130_fd_sc_hd__dfxtp_1 _475_ (.CLK(clknet_2_0__leaf_clk),
    .D(_034_),
    .Q(\clock_div[8] ));
 sky130_fd_sc_hd__dfxtp_1 _476_ (.CLK(clknet_2_3__leaf_clk),
    .D(_035_),
    .Q(\tempo_LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _477_ (.CLK(clknet_2_3__leaf_clk),
    .D(_036_),
    .Q(\tempo_LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _478_ (.CLK(clknet_2_3__leaf_clk),
    .D(_037_),
    .Q(\tempo_LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _479_ (.CLK(clknet_2_3__leaf_clk),
    .D(_038_),
    .Q(\tempo_LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_2 _480_ (.CLK(clknet_2_0__leaf_clk),
    .D(net1),
    .Q(just_rst));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__427__B1 (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__409__S (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__C1 (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__361__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__354__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__302__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__B (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__242__A (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__254__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B1 (.DIODE(net1));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_225 ();
endmodule

