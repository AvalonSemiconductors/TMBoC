magic
tech sky130B
magscale 1 2
timestamp 1683540519
<< viali >>
rect 4905 33541 4939 33575
rect 7849 33541 7883 33575
rect 10793 33541 10827 33575
rect 14473 33541 14507 33575
rect 17049 33541 17083 33575
rect 19717 33541 19751 33575
rect 22661 33541 22695 33575
rect 25605 33541 25639 33575
rect 28549 33541 28583 33575
rect 31493 33541 31527 33575
rect 34253 33541 34287 33575
rect 10977 33337 11011 33371
rect 14289 33337 14323 33371
rect 16865 33337 16899 33371
rect 19533 33337 19567 33371
rect 22477 33337 22511 33371
rect 25421 33337 25455 33371
rect 28365 33337 28399 33371
rect 31309 33337 31343 33371
rect 34069 33337 34103 33371
rect 4997 33269 5031 33303
rect 7941 33269 7975 33303
rect 20637 32929 20671 32963
rect 10241 32861 10275 32895
rect 16313 32861 16347 32895
rect 16497 32861 16531 32895
rect 16589 32861 16623 32895
rect 20545 32861 20579 32895
rect 22385 32861 22419 32895
rect 15853 32793 15887 32827
rect 10149 32725 10183 32759
rect 20913 32725 20947 32759
rect 22293 32725 22327 32759
rect 12265 32521 12299 32555
rect 13461 32521 13495 32555
rect 17325 32521 17359 32555
rect 18061 32521 18095 32555
rect 12357 32453 12391 32487
rect 13277 32453 13311 32487
rect 13553 32453 13587 32487
rect 21189 32453 21223 32487
rect 22109 32453 22143 32487
rect 9873 32385 9907 32419
rect 10425 32385 10459 32419
rect 10517 32385 10551 32419
rect 12081 32385 12115 32419
rect 16129 32385 16163 32419
rect 16313 32385 16347 32419
rect 17233 32385 17267 32419
rect 18061 32385 18095 32419
rect 18245 32385 18279 32419
rect 21097 32385 21131 32419
rect 22017 32385 22051 32419
rect 22201 32385 22235 32419
rect 23029 32385 23063 32419
rect 23213 32385 23247 32419
rect 24501 32385 24535 32419
rect 24685 32385 24719 32419
rect 27721 32385 27755 32419
rect 28089 32385 28123 32419
rect 30481 32385 30515 32419
rect 33333 32385 33367 32419
rect 10701 32317 10735 32351
rect 16221 32317 16255 32351
rect 17417 32317 17451 32351
rect 21281 32317 21315 32351
rect 27169 32317 27203 32351
rect 16865 32249 16899 32283
rect 20729 32249 20763 32283
rect 22937 32249 22971 32283
rect 9873 32181 9907 32215
rect 10609 32181 10643 32215
rect 11805 32181 11839 32215
rect 13001 32181 13035 32215
rect 24593 32181 24627 32215
rect 30297 32181 30331 32215
rect 33149 32181 33183 32215
rect 15761 31977 15795 32011
rect 15945 31977 15979 32011
rect 18061 31977 18095 32011
rect 21281 31977 21315 32011
rect 23673 31977 23707 32011
rect 9321 31909 9355 31943
rect 11161 31909 11195 31943
rect 18337 31909 18371 31943
rect 24593 31909 24627 31943
rect 8493 31841 8527 31875
rect 9781 31841 9815 31875
rect 9873 31841 9907 31875
rect 11621 31841 11655 31875
rect 13553 31841 13587 31875
rect 14381 31841 14415 31875
rect 17141 31841 17175 31875
rect 19441 31841 19475 31875
rect 22017 31841 22051 31875
rect 22569 31841 22603 31875
rect 23029 31841 23063 31875
rect 25053 31841 25087 31875
rect 25145 31841 25179 31875
rect 8401 31773 8435 31807
rect 8585 31773 8619 31807
rect 9689 31773 9723 31807
rect 12633 31773 12667 31807
rect 13461 31773 13495 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 16405 31773 16439 31807
rect 17233 31773 17267 31807
rect 17325 31773 17359 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 20269 31773 20303 31807
rect 20453 31773 20487 31807
rect 21005 31773 21039 31807
rect 21281 31773 21315 31807
rect 22845 31773 22879 31807
rect 23765 31773 23799 31807
rect 23857 31773 23891 31807
rect 26433 31773 26467 31807
rect 26617 31773 26651 31807
rect 11621 31705 11655 31739
rect 11713 31705 11747 31739
rect 15577 31705 15611 31739
rect 16865 31705 16899 31739
rect 21097 31705 21131 31739
rect 15777 31637 15811 31671
rect 23489 31637 23523 31671
rect 24961 31637 24995 31671
rect 9505 31433 9539 31467
rect 13553 31433 13587 31467
rect 16129 31433 16163 31467
rect 17049 31433 17083 31467
rect 17601 31433 17635 31467
rect 20846 31433 20880 31467
rect 24777 31433 24811 31467
rect 25881 31433 25915 31467
rect 28641 31433 28675 31467
rect 10333 31365 10367 31399
rect 10701 31365 10735 31399
rect 16865 31365 16899 31399
rect 22201 31365 22235 31399
rect 9137 31297 9171 31331
rect 10241 31297 10275 31331
rect 13185 31297 13219 31331
rect 14105 31297 14139 31331
rect 14841 31297 14875 31331
rect 14933 31297 14967 31331
rect 16129 31297 16163 31331
rect 16313 31297 16347 31331
rect 17141 31297 17175 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 20637 31297 20671 31331
rect 21097 31297 21131 31331
rect 22661 31297 22695 31331
rect 22937 31297 22971 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 23489 31297 23523 31331
rect 24225 31297 24259 31331
rect 25237 31297 25271 31331
rect 25421 31297 25455 31331
rect 25697 31297 25731 31331
rect 27353 31297 27387 31331
rect 27629 31297 27663 31331
rect 28579 31297 28613 31331
rect 9229 31229 9263 31263
rect 10425 31229 10459 31263
rect 13277 31229 13311 31263
rect 20545 31229 20579 31263
rect 24501 31229 24535 31263
rect 25605 31229 25639 31263
rect 27169 31229 27203 31263
rect 29101 31229 29135 31263
rect 10885 31161 10919 31195
rect 16865 31161 16899 31195
rect 25513 31161 25547 31195
rect 14289 31093 14323 31127
rect 24593 31093 24627 31127
rect 28457 31093 28491 31127
rect 29009 31093 29043 31127
rect 9413 30889 9447 30923
rect 10057 30889 10091 30923
rect 10701 30889 10735 30923
rect 13553 30889 13587 30923
rect 21005 30889 21039 30923
rect 22753 30889 22787 30923
rect 23121 30821 23155 30855
rect 27537 30821 27571 30855
rect 13461 30753 13495 30787
rect 13645 30753 13679 30787
rect 15761 30753 15795 30787
rect 20637 30753 20671 30787
rect 9321 30685 9355 30719
rect 9505 30685 9539 30719
rect 9965 30685 9999 30719
rect 10149 30685 10183 30719
rect 10609 30685 10643 30719
rect 10793 30685 10827 30719
rect 13737 30685 13771 30719
rect 14657 30685 14691 30719
rect 15025 30685 15059 30719
rect 15577 30685 15611 30719
rect 16037 30685 16071 30719
rect 16221 30685 16255 30719
rect 20821 30685 20855 30719
rect 22937 30685 22971 30719
rect 23213 30685 23247 30719
rect 25053 30685 25087 30719
rect 25605 30685 25639 30719
rect 25789 30685 25823 30719
rect 26249 30685 26283 30719
rect 27721 30685 27755 30719
rect 28089 30685 28123 30719
rect 28457 30685 28491 30719
rect 28917 30685 28951 30719
rect 26157 30617 26191 30651
rect 29745 30345 29779 30379
rect 28089 30277 28123 30311
rect 28549 30277 28583 30311
rect 14289 30209 14323 30243
rect 14933 30209 14967 30243
rect 19717 30209 19751 30243
rect 20269 30209 20303 30243
rect 21005 30209 21039 30243
rect 24685 30209 24719 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25789 30209 25823 30243
rect 25881 30209 25915 30243
rect 26065 30209 26099 30243
rect 27353 30209 27387 30243
rect 27629 30209 27663 30243
rect 28733 30209 28767 30243
rect 29009 30209 29043 30243
rect 29193 30209 29227 30243
rect 29653 30209 29687 30243
rect 29837 30209 29871 30243
rect 27445 30141 27479 30175
rect 13461 30005 13495 30039
rect 20913 30005 20947 30039
rect 14841 29801 14875 29835
rect 25053 29801 25087 29835
rect 10425 29733 10459 29767
rect 27353 29733 27387 29767
rect 27721 29733 27755 29767
rect 30021 29733 30055 29767
rect 20453 29665 20487 29699
rect 21557 29665 21591 29699
rect 28825 29665 28859 29699
rect 9689 29597 9723 29631
rect 9965 29597 9999 29631
rect 10425 29597 10459 29631
rect 10517 29597 10551 29631
rect 13001 29597 13035 29631
rect 13185 29597 13219 29631
rect 14933 29597 14967 29631
rect 19625 29597 19659 29631
rect 20177 29597 20211 29631
rect 21005 29597 21039 29631
rect 21373 29597 21407 29631
rect 24777 29597 24811 29631
rect 24869 29597 24903 29631
rect 27537 29597 27571 29631
rect 27629 29597 27663 29631
rect 27813 29597 27847 29631
rect 28365 29597 28399 29631
rect 28549 29597 28583 29631
rect 28917 29597 28951 29631
rect 29745 29597 29779 29631
rect 29929 29597 29963 29631
rect 10701 29529 10735 29563
rect 15117 29529 15151 29563
rect 9505 29461 9539 29495
rect 9873 29461 9907 29495
rect 12817 29461 12851 29495
rect 19533 29461 19567 29495
rect 21373 29461 21407 29495
rect 14565 29257 14599 29291
rect 20177 29257 20211 29291
rect 22109 29257 22143 29291
rect 27905 29257 27939 29291
rect 28933 29257 28967 29291
rect 29101 29257 29135 29291
rect 15393 29189 15427 29223
rect 17693 29189 17727 29223
rect 25237 29189 25271 29223
rect 27261 29189 27295 29223
rect 28733 29189 28767 29223
rect 9045 29121 9079 29155
rect 9321 29121 9355 29155
rect 9505 29121 9539 29155
rect 11897 29121 11931 29155
rect 12541 29121 12575 29155
rect 12633 29121 12667 29155
rect 12909 29121 12943 29155
rect 13185 29121 13219 29155
rect 14749 29121 14783 29155
rect 15577 29121 15611 29155
rect 15761 29121 15795 29155
rect 19165 29121 19199 29155
rect 19533 29121 19567 29155
rect 20361 29121 20395 29155
rect 20453 29121 20487 29155
rect 20637 29121 20671 29155
rect 20729 29121 20763 29155
rect 21189 29121 21223 29155
rect 21373 29121 21407 29155
rect 22293 29121 22327 29155
rect 22569 29121 22603 29155
rect 22753 29121 22787 29155
rect 25329 29121 25363 29155
rect 25605 29121 25639 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 28089 29121 28123 29155
rect 12449 29053 12483 29087
rect 14933 29053 14967 29087
rect 28273 29053 28307 29087
rect 21281 28985 21315 29019
rect 22385 28985 22419 29019
rect 22477 28985 22511 29019
rect 9413 28917 9447 28951
rect 28917 28917 28951 28951
rect 21189 28713 21223 28747
rect 28825 28713 28859 28747
rect 15209 28645 15243 28679
rect 10977 28577 11011 28611
rect 11621 28577 11655 28611
rect 13185 28577 13219 28611
rect 13369 28577 13403 28611
rect 26249 28577 26283 28611
rect 9321 28509 9355 28543
rect 9597 28509 9631 28543
rect 11253 28509 11287 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 13093 28509 13127 28543
rect 13277 28509 13311 28543
rect 14565 28509 14599 28543
rect 14933 28509 14967 28543
rect 15393 28509 15427 28543
rect 16313 28509 16347 28543
rect 16681 28509 16715 28543
rect 19901 28509 19935 28543
rect 19993 28509 20027 28543
rect 20637 28509 20671 28543
rect 20729 28509 20763 28543
rect 20913 28509 20947 28543
rect 21005 28509 21039 28543
rect 23305 28509 23339 28543
rect 23949 28509 23983 28543
rect 28733 28509 28767 28543
rect 20177 28441 20211 28475
rect 9137 28373 9171 28407
rect 9505 28373 9539 28407
rect 12909 28373 12943 28407
rect 27261 28373 27295 28407
rect 8125 28169 8159 28203
rect 15393 28169 15427 28203
rect 22293 28169 22327 28203
rect 23213 28169 23247 28203
rect 15945 28101 15979 28135
rect 20637 28101 20671 28135
rect 30205 28101 30239 28135
rect 7941 28033 7975 28067
rect 8217 28033 8251 28067
rect 9045 28033 9079 28067
rect 9689 28033 9723 28067
rect 9873 28033 9907 28067
rect 11897 28033 11931 28067
rect 12541 28033 12575 28067
rect 12909 28033 12943 28067
rect 13369 28033 13403 28067
rect 13829 28033 13863 28067
rect 14013 28033 14047 28067
rect 14197 28033 14231 28067
rect 15393 28033 15427 28067
rect 19257 28033 19291 28067
rect 19441 28033 19475 28067
rect 20269 28033 20303 28067
rect 20545 28033 20579 28067
rect 23673 28033 23707 28067
rect 25053 28033 25087 28067
rect 25697 28033 25731 28067
rect 27261 28033 27295 28067
rect 27537 28033 27571 28067
rect 30021 28033 30055 28067
rect 30297 28033 30331 28067
rect 8769 27965 8803 27999
rect 8861 27965 8895 27999
rect 8953 27965 8987 27999
rect 12449 27965 12483 27999
rect 15301 27965 15335 27999
rect 19349 27965 19383 27999
rect 22753 27965 22787 27999
rect 26065 27965 26099 27999
rect 27169 27965 27203 27999
rect 22477 27897 22511 27931
rect 23397 27897 23431 27931
rect 24869 27897 24903 27931
rect 7757 27829 7791 27863
rect 9229 27829 9263 27863
rect 9781 27829 9815 27863
rect 29837 27829 29871 27863
rect 16865 27557 16899 27591
rect 25237 27557 25271 27591
rect 27905 27557 27939 27591
rect 9229 27489 9263 27523
rect 12817 27489 12851 27523
rect 28457 27489 28491 27523
rect 9321 27421 9355 27455
rect 9689 27421 9723 27455
rect 13185 27421 13219 27455
rect 13369 27421 13403 27455
rect 14933 27421 14967 27455
rect 15945 27421 15979 27455
rect 16037 27421 16071 27455
rect 16221 27421 16255 27455
rect 18245 27421 18279 27455
rect 22017 27421 22051 27455
rect 22293 27421 22327 27455
rect 25421 27421 25455 27455
rect 25697 27421 25731 27455
rect 25973 27421 26007 27455
rect 26617 27421 26651 27455
rect 26893 27421 26927 27455
rect 27445 27421 27479 27455
rect 27721 27421 27755 27455
rect 28365 27421 28399 27455
rect 28549 27421 28583 27455
rect 29837 27421 29871 27455
rect 10149 27353 10183 27387
rect 14381 27353 14415 27387
rect 16405 27353 16439 27387
rect 17978 27353 18012 27387
rect 30104 27353 30138 27387
rect 22109 27285 22143 27319
rect 22477 27285 22511 27319
rect 27537 27285 27571 27319
rect 31217 27285 31251 27319
rect 19533 27081 19567 27115
rect 31125 27081 31159 27115
rect 8309 27013 8343 27047
rect 15485 27013 15519 27047
rect 22661 27013 22695 27047
rect 27537 27013 27571 27047
rect 8217 26945 8251 26979
rect 8493 26945 8527 26979
rect 9229 26945 9263 26979
rect 11897 26945 11931 26979
rect 12081 26945 12115 26979
rect 12173 26945 12207 26979
rect 13645 26945 13679 26979
rect 15669 26945 15703 26979
rect 15853 26945 15887 26979
rect 18245 26945 18279 26979
rect 21005 26945 21039 26979
rect 21189 26945 21223 26979
rect 21281 26945 21315 26979
rect 22109 26945 22143 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25605 26945 25639 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 27261 26945 27295 26979
rect 27445 26945 27479 26979
rect 30021 26945 30055 26979
rect 9045 26877 9079 26911
rect 9137 26877 9171 26911
rect 9321 26877 9355 26911
rect 26433 26877 26467 26911
rect 29745 26877 29779 26911
rect 8493 26809 8527 26843
rect 9505 26741 9539 26775
rect 11713 26741 11747 26775
rect 13645 26741 13679 26775
rect 20821 26741 20855 26775
rect 12357 26537 12391 26571
rect 13461 26537 13495 26571
rect 16681 26537 16715 26571
rect 25237 26537 25271 26571
rect 27077 26537 27111 26571
rect 32229 26537 32263 26571
rect 9413 26469 9447 26503
rect 13277 26469 13311 26503
rect 31309 26469 31343 26503
rect 11161 26401 11195 26435
rect 11713 26401 11747 26435
rect 12725 26401 12759 26435
rect 18061 26401 18095 26435
rect 27721 26401 27755 26435
rect 11345 26333 11379 26367
rect 12633 26333 12667 26367
rect 19625 26333 19659 26367
rect 19809 26333 19843 26367
rect 19901 26333 19935 26367
rect 25421 26333 25455 26367
rect 25513 26333 25547 26367
rect 25605 26333 25639 26367
rect 25697 26333 25731 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 26617 26333 26651 26367
rect 26801 26333 26835 26367
rect 26893 26333 26927 26367
rect 27537 26333 27571 26367
rect 32413 26333 32447 26367
rect 32597 26333 32631 26367
rect 32689 26333 32723 26367
rect 9137 26265 9171 26299
rect 11621 26265 11655 26299
rect 13429 26265 13463 26299
rect 13645 26265 13679 26299
rect 17794 26265 17828 26299
rect 19441 26265 19475 26299
rect 22569 26265 22603 26299
rect 30021 26265 30055 26299
rect 9597 26197 9631 26231
rect 21097 26197 21131 26231
rect 12357 25993 12391 26027
rect 12449 25993 12483 26027
rect 16865 25993 16899 26027
rect 17233 25993 17267 26027
rect 25605 25993 25639 26027
rect 27169 25993 27203 26027
rect 29929 25993 29963 26027
rect 10517 25925 10551 25959
rect 12081 25925 12115 25959
rect 12265 25925 12299 25959
rect 13093 25925 13127 25959
rect 13369 25925 13403 25959
rect 21373 25925 21407 25959
rect 24593 25925 24627 25959
rect 25145 25925 25179 25959
rect 9505 25857 9539 25891
rect 9721 25857 9755 25891
rect 10425 25857 10459 25891
rect 10701 25857 10735 25891
rect 13277 25857 13311 25891
rect 13466 25857 13500 25891
rect 17049 25857 17083 25891
rect 17325 25857 17359 25891
rect 19625 25857 19659 25891
rect 20821 25857 20855 25891
rect 22017 25857 22051 25891
rect 22293 25857 22327 25891
rect 24501 25857 24535 25891
rect 24685 25857 24719 25891
rect 26525 25857 26559 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 28641 25857 28675 25891
rect 32505 25857 32539 25891
rect 32689 25857 32723 25891
rect 32781 25857 32815 25891
rect 9597 25789 9631 25823
rect 9965 25789 9999 25823
rect 23489 25789 23523 25823
rect 27353 25789 27387 25823
rect 27629 25789 27663 25823
rect 10701 25721 10735 25755
rect 25421 25721 25455 25755
rect 12633 25653 12667 25687
rect 13093 25653 13127 25687
rect 18337 25653 18371 25687
rect 26341 25653 26375 25687
rect 32321 25653 32355 25687
rect 15393 25449 15427 25483
rect 19809 25449 19843 25483
rect 26065 25449 26099 25483
rect 26249 25449 26283 25483
rect 28273 25449 28307 25483
rect 16313 25381 16347 25415
rect 26617 25381 26651 25415
rect 21189 25313 21223 25347
rect 3433 25245 3467 25279
rect 4077 25245 4111 25279
rect 4353 25245 4387 25279
rect 6745 25245 6779 25279
rect 6929 25245 6963 25279
rect 12265 25245 12299 25279
rect 12541 25245 12575 25279
rect 12725 25245 12759 25279
rect 16037 25245 16071 25279
rect 16313 25245 16347 25279
rect 20922 25245 20956 25279
rect 24593 25245 24627 25279
rect 27352 25245 27386 25279
rect 27445 25245 27479 25279
rect 28365 25245 28399 25279
rect 30113 25245 30147 25279
rect 3985 25177 4019 25211
rect 15577 25177 15611 25211
rect 21649 25177 21683 25211
rect 24869 25177 24903 25211
rect 26249 25177 26283 25211
rect 30380 25177 30414 25211
rect 3341 25109 3375 25143
rect 6745 25109 6779 25143
rect 12081 25109 12115 25143
rect 15209 25109 15243 25143
rect 15377 25109 15411 25143
rect 16129 25109 16163 25143
rect 22937 25109 22971 25143
rect 27077 25109 27111 25143
rect 31493 25109 31527 25143
rect 25145 24905 25179 24939
rect 5273 24837 5307 24871
rect 28641 24837 28675 24871
rect 28825 24837 28859 24871
rect 2329 24769 2363 24803
rect 6929 24769 6963 24803
rect 14749 24769 14783 24803
rect 15025 24769 15059 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 15853 24769 15887 24803
rect 16037 24769 16071 24803
rect 18153 24769 18187 24803
rect 21005 24769 21039 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 21465 24769 21499 24803
rect 22273 24769 22307 24803
rect 25237 24769 25271 24803
rect 25329 24769 25363 24803
rect 26157 24769 26191 24803
rect 29101 24769 29135 24803
rect 30380 24769 30414 24803
rect 2605 24701 2639 24735
rect 4721 24701 4755 24735
rect 7941 24701 7975 24735
rect 17877 24701 17911 24735
rect 19349 24701 19383 24735
rect 22017 24701 22051 24735
rect 26433 24701 26467 24735
rect 30113 24701 30147 24735
rect 15209 24633 15243 24667
rect 26341 24633 26375 24667
rect 31493 24633 31527 24667
rect 3893 24565 3927 24599
rect 16037 24565 16071 24599
rect 23397 24565 23431 24599
rect 25973 24565 26007 24599
rect 28825 24565 28859 24599
rect 2789 24361 2823 24395
rect 6837 24361 6871 24395
rect 22845 24361 22879 24395
rect 30573 24361 30607 24395
rect 2329 24293 2363 24327
rect 5273 24293 5307 24327
rect 2973 24225 3007 24259
rect 4169 24225 4203 24259
rect 4353 24225 4387 24259
rect 5181 24225 5215 24259
rect 15853 24225 15887 24259
rect 21005 24225 21039 24259
rect 2053 24157 2087 24191
rect 3065 24157 3099 24191
rect 4445 24157 4479 24191
rect 4537 24157 4571 24191
rect 4629 24157 4663 24191
rect 5549 24157 5583 24191
rect 5733 24157 5767 24191
rect 7573 24157 7607 24191
rect 8493 24157 8527 24191
rect 11897 24157 11931 24191
rect 12081 24157 12115 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15669 24157 15703 24191
rect 17049 24157 17083 24191
rect 17233 24157 17267 24191
rect 17877 24157 17911 24191
rect 18153 24157 18187 24191
rect 20637 24157 20671 24191
rect 20821 24157 20855 24191
rect 21465 24157 21499 24191
rect 23489 24157 23523 24191
rect 23765 24157 23799 24191
rect 25237 24157 25271 24191
rect 25421 24157 25455 24191
rect 30757 24157 30791 24191
rect 30941 24157 30975 24191
rect 31033 24157 31067 24191
rect 2329 24089 2363 24123
rect 3341 24089 3375 24123
rect 3433 24089 3467 24123
rect 18061 24089 18095 24123
rect 21732 24089 21766 24123
rect 23305 24089 23339 24123
rect 2145 24021 2179 24055
rect 12081 24021 12115 24055
rect 14289 24021 14323 24055
rect 15485 24021 15519 24055
rect 17141 24021 17175 24055
rect 17693 24021 17727 24055
rect 23673 24021 23707 24055
rect 25329 24021 25363 24055
rect 5089 23817 5123 23851
rect 14933 23817 14967 23851
rect 15117 23817 15151 23851
rect 15945 23817 15979 23851
rect 30113 23817 30147 23851
rect 4629 23749 4663 23783
rect 16129 23749 16163 23783
rect 19993 23749 20027 23783
rect 22109 23749 22143 23783
rect 28641 23749 28675 23783
rect 2789 23681 2823 23715
rect 3709 23681 3743 23715
rect 5457 23681 5491 23715
rect 5549 23681 5583 23715
rect 9229 23681 9263 23715
rect 9873 23681 9907 23715
rect 10057 23681 10091 23715
rect 12909 23681 12943 23715
rect 13277 23681 13311 23715
rect 14381 23681 14415 23715
rect 16313 23681 16347 23715
rect 20453 23681 20487 23715
rect 20729 23681 20763 23715
rect 22661 23681 22695 23715
rect 25513 23681 25547 23715
rect 5273 23613 5307 23647
rect 5365 23613 5399 23647
rect 6837 23613 6871 23647
rect 7113 23613 7147 23647
rect 8493 23613 8527 23647
rect 9413 23613 9447 23647
rect 12265 23613 12299 23647
rect 13001 23613 13035 23647
rect 13185 23613 13219 23647
rect 14841 23613 14875 23647
rect 15209 23613 15243 23647
rect 15301 23613 15335 23647
rect 20821 23613 20855 23647
rect 9965 23545 9999 23579
rect 14289 23545 14323 23579
rect 18705 23545 18739 23579
rect 9045 23477 9079 23511
rect 15485 23477 15519 23511
rect 25421 23477 25455 23511
rect 3249 23273 3283 23307
rect 3341 23273 3375 23307
rect 4169 23273 4203 23307
rect 6929 23273 6963 23307
rect 10333 23273 10367 23307
rect 18705 23273 18739 23307
rect 21925 23273 21959 23307
rect 9137 23205 9171 23239
rect 15577 23205 15611 23239
rect 16129 23205 16163 23239
rect 19717 23205 19751 23239
rect 3433 23137 3467 23171
rect 8125 23137 8159 23171
rect 8217 23137 8251 23171
rect 8309 23137 8343 23171
rect 8401 23137 8435 23171
rect 8585 23137 8619 23171
rect 11805 23137 11839 23171
rect 15117 23137 15151 23171
rect 15209 23137 15243 23171
rect 15301 23137 15335 23171
rect 16497 23137 16531 23171
rect 17325 23137 17359 23171
rect 24961 23137 24995 23171
rect 25329 23137 25363 23171
rect 32689 23137 32723 23171
rect 33149 23137 33183 23171
rect 3157 23069 3191 23103
rect 7113 23069 7147 23103
rect 7205 23069 7239 23103
rect 7573 23069 7607 23103
rect 9413 23069 9447 23103
rect 12081 23069 12115 23103
rect 12541 23069 12575 23103
rect 15393 23069 15427 23103
rect 17592 23069 17626 23103
rect 19441 23069 19475 23103
rect 19717 23069 19751 23103
rect 20637 23069 20671 23103
rect 24869 23069 24903 23103
rect 27537 23069 27571 23103
rect 28089 23069 28123 23103
rect 28273 23069 28307 23103
rect 31769 23069 31803 23103
rect 32045 23069 32079 23103
rect 32781 23069 32815 23103
rect 33609 23069 33643 23103
rect 33793 23069 33827 23103
rect 4353 23001 4387 23035
rect 7297 23001 7331 23035
rect 7435 23001 7469 23035
rect 9137 23001 9171 23035
rect 13277 23001 13311 23035
rect 24685 23001 24719 23035
rect 27813 23001 27847 23035
rect 3985 22933 4019 22967
rect 4153 22933 4187 22967
rect 9321 22933 9355 22967
rect 16037 22933 16071 22967
rect 25145 22933 25179 22967
rect 25237 22933 25271 22967
rect 31033 22933 31067 22967
rect 33701 22933 33735 22967
rect 7205 22729 7239 22763
rect 32413 22729 32447 22763
rect 8125 22661 8159 22695
rect 8309 22661 8343 22695
rect 8493 22661 8527 22695
rect 9689 22661 9723 22695
rect 12541 22661 12575 22695
rect 14381 22661 14415 22695
rect 18613 22661 18647 22695
rect 23765 22661 23799 22695
rect 25237 22661 25271 22695
rect 33057 22661 33091 22695
rect 33517 22661 33551 22695
rect 4445 22593 4479 22627
rect 7389 22593 7423 22627
rect 7573 22593 7607 22627
rect 7665 22593 7699 22627
rect 9413 22593 9447 22627
rect 9505 22593 9539 22627
rect 10333 22593 10367 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 12909 22593 12943 22627
rect 13277 22593 13311 22627
rect 13369 22593 13403 22627
rect 13645 22593 13679 22627
rect 13921 22593 13955 22627
rect 14657 22593 14691 22627
rect 15301 22593 15335 22627
rect 15485 22593 15519 22627
rect 15577 22593 15611 22627
rect 17325 22593 17359 22627
rect 17509 22593 17543 22627
rect 19993 22593 20027 22627
rect 20085 22593 20119 22627
rect 20269 22593 20303 22627
rect 20361 22593 20395 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 23673 22593 23707 22627
rect 24869 22593 24903 22627
rect 28181 22593 28215 22627
rect 28825 22593 28859 22627
rect 29929 22593 29963 22627
rect 30113 22593 30147 22627
rect 31309 22593 31343 22627
rect 32689 22593 32723 22627
rect 33701 22593 33735 22627
rect 10977 22525 11011 22559
rect 14381 22525 14415 22559
rect 18153 22525 18187 22559
rect 18245 22525 18279 22559
rect 24777 22525 24811 22559
rect 25145 22525 25179 22559
rect 29745 22525 29779 22559
rect 31033 22525 31067 22559
rect 31125 22525 31159 22559
rect 31217 22525 31251 22559
rect 32551 22525 32585 22559
rect 32965 22525 32999 22559
rect 4537 22457 4571 22491
rect 17417 22457 17451 22491
rect 22017 22457 22051 22491
rect 11805 22389 11839 22423
rect 14565 22389 14599 22423
rect 15117 22389 15151 22423
rect 17969 22389 18003 22423
rect 19809 22389 19843 22423
rect 24593 22389 24627 22423
rect 27353 22389 27387 22423
rect 30849 22389 30883 22423
rect 33793 22389 33827 22423
rect 11725 22185 11759 22219
rect 23213 22185 23247 22219
rect 33517 22185 33551 22219
rect 12821 22117 12855 22151
rect 23029 22117 23063 22151
rect 10241 22049 10275 22083
rect 11989 22049 12023 22083
rect 17785 22049 17819 22083
rect 25053 22049 25087 22083
rect 26985 22049 27019 22083
rect 30021 22049 30055 22083
rect 33149 22049 33183 22083
rect 7205 21981 7239 22015
rect 8585 21981 8619 22015
rect 12725 21981 12759 22015
rect 12909 21981 12943 22015
rect 13001 21981 13035 22015
rect 17969 21981 18003 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 20821 21981 20855 22015
rect 23213 21981 23247 22015
rect 23397 21981 23431 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 24961 21981 24995 22015
rect 26065 21981 26099 22015
rect 26249 21981 26283 22015
rect 27261 21981 27295 22015
rect 27813 21981 27847 22015
rect 28641 21981 28675 22015
rect 30113 21981 30147 22015
rect 31033 21981 31067 22015
rect 31401 21981 31435 22015
rect 31585 21981 31619 22015
rect 32045 21981 32079 22015
rect 32413 21981 32447 22015
rect 32597 21981 32631 22015
rect 33333 21981 33367 22015
rect 19809 21913 19843 21947
rect 20177 21913 20211 21947
rect 26157 21913 26191 21947
rect 28273 21913 28307 21947
rect 28457 21913 28491 21947
rect 31125 21913 31159 21947
rect 32137 21913 32171 21947
rect 7205 21845 7239 21879
rect 8493 21845 8527 21879
rect 12541 21845 12575 21879
rect 22293 21845 22327 21879
rect 25237 21845 25271 21879
rect 27721 21845 27755 21879
rect 29745 21845 29779 21879
rect 27169 21641 27203 21675
rect 30297 21641 30331 21675
rect 31677 21641 31711 21675
rect 11713 21573 11747 21607
rect 30481 21573 30515 21607
rect 2881 21505 2915 21539
rect 3801 21505 3835 21539
rect 4077 21505 4111 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 14473 21505 14507 21539
rect 14565 21505 14599 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 19533 21505 19567 21539
rect 19809 21505 19843 21539
rect 20545 21505 20579 21539
rect 20637 21505 20671 21539
rect 22017 21505 22051 21539
rect 22293 21505 22327 21539
rect 27537 21505 27571 21539
rect 28181 21505 28215 21539
rect 28365 21505 28399 21539
rect 30205 21505 30239 21539
rect 31493 21505 31527 21539
rect 31677 21505 31711 21539
rect 2973 21437 3007 21471
rect 3157 21437 3191 21471
rect 22385 21437 22419 21471
rect 23213 21437 23247 21471
rect 23489 21437 23523 21471
rect 24593 21437 24627 21471
rect 27445 21437 27479 21471
rect 3893 21369 3927 21403
rect 3985 21369 4019 21403
rect 3065 21301 3099 21335
rect 3617 21301 3651 21335
rect 15485 21301 15519 21335
rect 19441 21301 19475 21335
rect 28365 21301 28399 21335
rect 30481 21301 30515 21335
rect 13461 21097 13495 21131
rect 14749 21097 14783 21131
rect 16129 21097 16163 21131
rect 21281 21097 21315 21131
rect 23581 21097 23615 21131
rect 32413 21097 32447 21131
rect 31309 21029 31343 21063
rect 7389 20961 7423 20995
rect 20085 20961 20119 20995
rect 20177 20961 20211 20995
rect 33057 20961 33091 20995
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 7573 20893 7607 20927
rect 7665 20893 7699 20927
rect 10425 20893 10459 20927
rect 10609 20893 10643 20927
rect 10701 20893 10735 20927
rect 13553 20893 13587 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 17417 20893 17451 20927
rect 19717 20893 19751 20927
rect 19809 20893 19843 20927
rect 22569 20893 22603 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24777 20893 24811 20927
rect 25053 20893 25087 20927
rect 31584 20893 31618 20927
rect 31677 20893 31711 20927
rect 32229 20893 32263 20927
rect 32413 20893 32447 20927
rect 32965 20893 32999 20927
rect 33149 20893 33183 20927
rect 24593 20825 24627 20859
rect 3341 20757 3375 20791
rect 7389 20757 7423 20791
rect 10241 20757 10275 20791
rect 14381 20757 14415 20791
rect 19533 20757 19567 20791
rect 24961 20757 24995 20791
rect 7849 20553 7883 20587
rect 8401 20553 8435 20587
rect 19533 20553 19567 20587
rect 21097 20553 21131 20587
rect 31585 20553 31619 20587
rect 32597 20553 32631 20587
rect 3525 20485 3559 20519
rect 3617 20485 3651 20519
rect 7481 20485 7515 20519
rect 23213 20485 23247 20519
rect 3157 20417 3191 20451
rect 3249 20417 3283 20451
rect 4445 20417 4479 20451
rect 7389 20417 7423 20451
rect 7665 20417 7699 20451
rect 8309 20417 8343 20451
rect 8493 20417 8527 20451
rect 8585 20417 8619 20451
rect 11069 20417 11103 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 15117 20417 15151 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 19349 20417 19383 20451
rect 19625 20417 19659 20451
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 20821 20417 20855 20451
rect 20913 20417 20947 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 32781 20417 32815 20451
rect 33057 20417 33091 20451
rect 4077 20349 4111 20383
rect 4353 20349 4387 20383
rect 10425 20349 10459 20383
rect 14841 20349 14875 20383
rect 27629 20281 27663 20315
rect 32965 20281 32999 20315
rect 2973 20213 3007 20247
rect 13093 20213 13127 20247
rect 15853 20213 15887 20247
rect 19165 20213 19199 20247
rect 24501 20213 24535 20247
rect 27997 20213 28031 20247
rect 3985 20009 4019 20043
rect 7573 20009 7607 20043
rect 14473 20009 14507 20043
rect 18797 20009 18831 20043
rect 20085 20009 20119 20043
rect 5089 19941 5123 19975
rect 7113 19941 7147 19975
rect 7757 19941 7791 19975
rect 9137 19941 9171 19975
rect 32321 19941 32355 19975
rect 2421 19873 2455 19907
rect 3249 19873 3283 19907
rect 10517 19873 10551 19907
rect 11897 19873 11931 19907
rect 13737 19873 13771 19907
rect 22569 19873 22603 19907
rect 1685 19805 1719 19839
rect 1869 19805 1903 19839
rect 3157 19805 3191 19839
rect 4169 19805 4203 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 5365 19805 5399 19839
rect 6837 19805 6871 19839
rect 6929 19805 6963 19839
rect 7113 19805 7147 19839
rect 8033 19805 8067 19839
rect 9413 19805 9447 19839
rect 10425 19805 10459 19839
rect 10793 19805 10827 19839
rect 11069 19805 11103 19839
rect 11713 19805 11747 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14381 19805 14415 19839
rect 15117 19805 15151 19839
rect 16865 19805 16899 19839
rect 18521 19805 18555 19839
rect 19441 19805 19475 19839
rect 19534 19805 19568 19839
rect 19717 19805 19751 19839
rect 19809 19805 19843 19839
rect 19906 19805 19940 19839
rect 31953 19805 31987 19839
rect 32229 19805 32263 19839
rect 32413 19805 32447 19839
rect 32597 19805 32631 19839
rect 1777 19737 1811 19771
rect 4261 19737 4295 19771
rect 4353 19737 4387 19771
rect 5089 19737 5123 19771
rect 9137 19737 9171 19771
rect 9321 19737 9355 19771
rect 15669 19737 15703 19771
rect 16313 19737 16347 19771
rect 20821 19737 20855 19771
rect 5273 19669 5307 19703
rect 11529 19669 11563 19703
rect 4445 19465 4479 19499
rect 16313 19465 16347 19499
rect 17233 19465 17267 19499
rect 20361 19465 20395 19499
rect 21189 19465 21223 19499
rect 32597 19465 32631 19499
rect 32873 19465 32907 19499
rect 2780 19397 2814 19431
rect 12449 19397 12483 19431
rect 24777 19397 24811 19431
rect 28365 19397 28399 19431
rect 32689 19397 32723 19431
rect 2513 19329 2547 19363
rect 4629 19329 4663 19363
rect 7113 19329 7147 19363
rect 7380 19329 7414 19363
rect 9045 19329 9079 19363
rect 9229 19329 9263 19363
rect 10701 19329 10735 19363
rect 12725 19329 12759 19363
rect 15200 19329 15234 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17325 19329 17359 19363
rect 18981 19329 19015 19363
rect 19248 19329 19282 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 23121 19329 23155 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 29009 19329 29043 19363
rect 29377 19329 29411 19363
rect 31217 19329 31251 19363
rect 31401 19329 31435 19363
rect 32321 19329 32355 19363
rect 32505 19329 32539 19363
rect 4813 19261 4847 19295
rect 10425 19261 10459 19295
rect 14933 19261 14967 19295
rect 20821 19261 20855 19295
rect 23397 19261 23431 19295
rect 28825 19261 28859 19295
rect 29285 19261 29319 19295
rect 3893 19193 3927 19227
rect 31401 19193 31435 19227
rect 8493 19125 8527 19159
rect 9137 19125 9171 19159
rect 10149 19125 10183 19159
rect 10609 19125 10643 19159
rect 27261 19125 27295 19159
rect 7665 18921 7699 18955
rect 14565 18921 14599 18955
rect 16681 18921 16715 18955
rect 18705 18921 18739 18955
rect 20821 18921 20855 18955
rect 25881 18921 25915 18955
rect 33149 18921 33183 18955
rect 3157 18853 3191 18887
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 8217 18785 8251 18819
rect 12357 18785 12391 18819
rect 26157 18785 26191 18819
rect 31861 18785 31895 18819
rect 32781 18785 32815 18819
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 8309 18717 8343 18751
rect 10425 18717 10459 18751
rect 10517 18717 10551 18751
rect 11989 18717 12023 18751
rect 12265 18717 12299 18751
rect 15301 18717 15335 18751
rect 19441 18717 19475 18751
rect 23765 18717 23799 18751
rect 24041 18717 24075 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 26065 18717 26099 18751
rect 26249 18717 26283 18751
rect 26341 18717 26375 18751
rect 27721 18717 27755 18751
rect 27905 18717 27939 18751
rect 28549 18717 28583 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29837 18717 29871 18751
rect 30021 18717 30055 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 32689 18717 32723 18751
rect 32965 18717 32999 18751
rect 3157 18649 3191 18683
rect 14381 18649 14415 18683
rect 14565 18649 14599 18683
rect 15568 18649 15602 18683
rect 18889 18649 18923 18683
rect 19708 18649 19742 18683
rect 27353 18649 27387 18683
rect 29745 18649 29779 18683
rect 8033 18581 8067 18615
rect 14749 18581 14783 18615
rect 18521 18581 18555 18615
rect 18705 18581 18739 18615
rect 23581 18581 23615 18615
rect 23949 18581 23983 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 28365 18581 28399 18615
rect 8217 18377 8251 18411
rect 15761 18377 15795 18411
rect 16129 18377 16163 18411
rect 25697 18377 25731 18411
rect 32781 18377 32815 18411
rect 6837 18309 6871 18343
rect 14749 18309 14783 18343
rect 19257 18309 19291 18343
rect 24869 18309 24903 18343
rect 8033 18241 8067 18275
rect 8217 18241 8251 18275
rect 10333 18241 10367 18275
rect 12265 18241 12299 18275
rect 12449 18241 12483 18275
rect 13001 18241 13035 18275
rect 15945 18241 15979 18275
rect 16221 18241 16255 18275
rect 23489 18241 23523 18275
rect 25329 18241 25363 18275
rect 27905 18241 27939 18275
rect 28733 18241 28767 18275
rect 29101 18241 29135 18275
rect 29377 18241 29411 18275
rect 29745 18241 29779 18275
rect 32505 18241 32539 18275
rect 6745 18173 6779 18207
rect 6929 18173 6963 18207
rect 12173 18173 12207 18207
rect 23213 18173 23247 18207
rect 25421 18173 25455 18207
rect 27537 18173 27571 18207
rect 27997 18173 28031 18207
rect 32321 18173 32355 18207
rect 32873 18173 32907 18207
rect 34345 18173 34379 18207
rect 7297 18105 7331 18139
rect 28641 18105 28675 18139
rect 10241 18037 10275 18071
rect 20545 18037 20579 18071
rect 25329 18037 25363 18071
rect 6469 17833 6503 17867
rect 21649 17833 21683 17867
rect 27997 17833 28031 17867
rect 32689 17833 32723 17867
rect 3433 17765 3467 17799
rect 13093 17697 13127 17731
rect 27629 17697 27663 17731
rect 28457 17697 28491 17731
rect 33609 17697 33643 17731
rect 3249 17629 3283 17663
rect 6377 17629 6411 17663
rect 6561 17629 6595 17663
rect 15209 17629 15243 17663
rect 17601 17629 17635 17663
rect 17877 17629 17911 17663
rect 18429 17629 18463 17663
rect 18705 17629 18739 17663
rect 19441 17629 19475 17663
rect 21373 17629 21407 17663
rect 24777 17629 24811 17663
rect 25053 17629 25087 17663
rect 27537 17629 27571 17663
rect 27721 17629 27755 17663
rect 27813 17629 27847 17663
rect 28641 17629 28675 17663
rect 28917 17629 28951 17663
rect 30757 17629 30791 17663
rect 30941 17629 30975 17663
rect 31769 17629 31803 17663
rect 31953 17629 31987 17663
rect 32597 17629 32631 17663
rect 33241 17629 33275 17663
rect 33425 17629 33459 17663
rect 2881 17561 2915 17595
rect 12817 17561 12851 17595
rect 18889 17561 18923 17595
rect 19686 17561 19720 17595
rect 31125 17561 31159 17595
rect 31861 17561 31895 17595
rect 32413 17561 32447 17595
rect 3065 17493 3099 17527
rect 3157 17493 3191 17527
rect 11345 17493 11379 17527
rect 16497 17493 16531 17527
rect 17417 17493 17451 17527
rect 17785 17493 17819 17527
rect 18521 17493 18555 17527
rect 20821 17493 20855 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 28825 17493 28859 17527
rect 4445 17289 4479 17323
rect 25697 17289 25731 17323
rect 28549 17289 28583 17323
rect 30757 17289 30791 17323
rect 30941 17289 30975 17323
rect 32521 17289 32555 17323
rect 32689 17289 32723 17323
rect 33241 17289 33275 17323
rect 2973 17221 3007 17255
rect 9597 17221 9631 17255
rect 13277 17221 13311 17255
rect 18245 17221 18279 17255
rect 19809 17221 19843 17255
rect 20821 17221 20855 17255
rect 23388 17221 23422 17255
rect 25421 17221 25455 17255
rect 28641 17221 28675 17255
rect 29837 17221 29871 17255
rect 30849 17221 30883 17255
rect 31493 17221 31527 17255
rect 32321 17221 32355 17255
rect 6653 17153 6687 17187
rect 6745 17153 6779 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 9873 17153 9907 17187
rect 16221 17153 16255 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 20637 17153 20671 17187
rect 20913 17153 20947 17187
rect 25053 17153 25087 17187
rect 25146 17153 25180 17187
rect 25329 17153 25363 17187
rect 25518 17153 25552 17187
rect 26157 17153 26191 17187
rect 28549 17153 28583 17187
rect 28825 17153 28859 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30481 17153 30515 17187
rect 30625 17153 30659 17187
rect 31677 17153 31711 17187
rect 31769 17153 31803 17187
rect 33149 17153 33183 17187
rect 33333 17153 33367 17187
rect 2697 17085 2731 17119
rect 9781 17085 9815 17119
rect 13553 17085 13587 17119
rect 15945 17085 15979 17119
rect 23121 17085 23155 17119
rect 26433 17085 26467 17119
rect 31493 17017 31527 17051
rect 8217 16949 8251 16983
rect 9781 16949 9815 16983
rect 10057 16949 10091 16983
rect 11805 16949 11839 16983
rect 20453 16949 20487 16983
rect 24501 16949 24535 16983
rect 32505 16949 32539 16983
rect 3065 16745 3099 16779
rect 3249 16745 3283 16779
rect 4261 16745 4295 16779
rect 6837 16745 6871 16779
rect 9781 16745 9815 16779
rect 12265 16745 12299 16779
rect 21373 16745 21407 16779
rect 25973 16745 26007 16779
rect 31217 16745 31251 16779
rect 32229 16745 32263 16779
rect 5917 16677 5951 16711
rect 7205 16677 7239 16711
rect 14841 16677 14875 16711
rect 16681 16677 16715 16711
rect 7113 16609 7147 16643
rect 7334 16609 7368 16643
rect 15301 16609 15335 16643
rect 29745 16609 29779 16643
rect 32597 16609 32631 16643
rect 4077 16541 4111 16575
rect 4261 16541 4295 16575
rect 9689 16541 9723 16575
rect 9965 16541 9999 16575
rect 10055 16541 10089 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15568 16541 15602 16575
rect 17233 16541 17267 16575
rect 18337 16541 18371 16575
rect 18521 16541 18555 16575
rect 19441 16541 19475 16575
rect 19708 16541 19742 16575
rect 21557 16541 21591 16575
rect 24593 16541 24627 16575
rect 24860 16541 24894 16575
rect 26433 16541 26467 16575
rect 26709 16541 26743 16575
rect 29929 16541 29963 16575
rect 31217 16541 31251 16575
rect 31493 16541 31527 16575
rect 31621 16541 31655 16575
rect 32413 16541 32447 16575
rect 3433 16473 3467 16507
rect 5549 16473 5583 16507
rect 7481 16473 7515 16507
rect 14473 16473 14507 16507
rect 17601 16473 17635 16507
rect 18705 16473 18739 16507
rect 31401 16473 31435 16507
rect 3233 16405 3267 16439
rect 6009 16405 6043 16439
rect 10241 16405 10275 16439
rect 20821 16405 20855 16439
rect 30021 16405 30055 16439
rect 30113 16405 30147 16439
rect 30297 16405 30331 16439
rect 6745 16201 6779 16235
rect 13461 16201 13495 16235
rect 19533 16201 19567 16235
rect 20453 16201 20487 16235
rect 22661 16201 22695 16235
rect 33701 16201 33735 16235
rect 5733 16133 5767 16167
rect 15200 16133 15234 16167
rect 18245 16133 18279 16167
rect 20821 16133 20855 16167
rect 22293 16133 22327 16167
rect 26525 16133 26559 16167
rect 28641 16133 28675 16167
rect 5549 16065 5583 16099
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 9597 16065 9631 16099
rect 13277 16065 13311 16099
rect 14013 16065 14047 16099
rect 14289 16065 14323 16099
rect 16865 16065 16899 16099
rect 17049 16065 17083 16099
rect 20591 16065 20625 16099
rect 20729 16065 20763 16099
rect 20949 16065 20983 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 22110 16065 22144 16099
rect 22385 16065 22419 16099
rect 22523 16065 22557 16099
rect 25145 16065 25179 16099
rect 26341 16065 26375 16099
rect 26617 16065 26651 16099
rect 28549 16065 28583 16099
rect 28733 16065 28767 16099
rect 28917 16065 28951 16099
rect 29561 16065 29595 16099
rect 32588 16065 32622 16099
rect 5365 15997 5399 16031
rect 14933 15997 14967 16031
rect 17417 15997 17451 16031
rect 32321 15997 32355 16031
rect 8309 15861 8343 15895
rect 16313 15861 16347 15895
rect 23857 15861 23891 15895
rect 26157 15861 26191 15895
rect 28365 15861 28399 15895
rect 29469 15861 29503 15895
rect 5273 15657 5307 15691
rect 7757 15657 7791 15691
rect 9229 15657 9263 15691
rect 23765 15657 23799 15691
rect 26525 15657 26559 15691
rect 27997 15657 28031 15691
rect 31677 15657 31711 15691
rect 33885 15657 33919 15691
rect 7941 15589 7975 15623
rect 13645 15589 13679 15623
rect 7665 15521 7699 15555
rect 14933 15521 14967 15555
rect 18245 15521 18279 15555
rect 22569 15521 22603 15555
rect 28181 15521 28215 15555
rect 28365 15521 28399 15555
rect 2605 15453 2639 15487
rect 2881 15453 2915 15487
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 6745 15453 6779 15487
rect 7389 15453 7423 15487
rect 9137 15453 9171 15487
rect 10425 15453 10459 15487
rect 10977 15453 11011 15487
rect 11161 15453 11195 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 13369 15453 13403 15487
rect 13645 15453 13679 15487
rect 15025 15453 15059 15487
rect 15301 15453 15335 15487
rect 16129 15453 16163 15487
rect 16313 15453 16347 15487
rect 17693 15453 17727 15487
rect 17877 15453 17911 15487
rect 20821 15453 20855 15487
rect 24041 15453 24075 15487
rect 25237 15453 25271 15487
rect 28273 15453 28307 15487
rect 28457 15453 28491 15487
rect 33425 15453 33459 15487
rect 33701 15453 33735 15487
rect 2973 15385 3007 15419
rect 5457 15385 5491 15419
rect 23581 15385 23615 15419
rect 32965 15385 32999 15419
rect 5089 15317 5123 15351
rect 5257 15317 5291 15351
rect 6193 15317 6227 15351
rect 6837 15317 6871 15351
rect 10977 15317 11011 15351
rect 16313 15317 16347 15351
rect 23765 15317 23799 15351
rect 33517 15317 33551 15351
rect 5448 15113 5482 15147
rect 9137 15113 9171 15147
rect 16037 15113 16071 15147
rect 22385 15113 22419 15147
rect 33609 15113 33643 15147
rect 5825 15045 5859 15079
rect 9045 15045 9079 15079
rect 4169 14977 4203 15011
rect 9321 14977 9355 15011
rect 10425 14977 10459 15011
rect 10517 14977 10551 15011
rect 10701 14977 10735 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 17325 14977 17359 15011
rect 17509 14977 17543 15011
rect 18245 14977 18279 15011
rect 20637 14977 20671 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 22201 14977 22235 15011
rect 22477 14977 22511 15011
rect 25154 14977 25188 15011
rect 29837 14977 29871 15011
rect 32321 14977 32355 15011
rect 1685 14909 1719 14943
rect 1961 14909 1995 14943
rect 4077 14909 4111 14943
rect 11161 14909 11195 14943
rect 17785 14909 17819 14943
rect 25421 14909 25455 14943
rect 3433 14841 3467 14875
rect 29653 14841 29687 14875
rect 5273 14773 5307 14807
rect 5457 14773 5491 14807
rect 9597 14773 9631 14807
rect 19717 14773 19751 14807
rect 20453 14773 20487 14807
rect 22017 14773 22051 14807
rect 24041 14773 24075 14807
rect 6193 14569 6227 14603
rect 7205 14569 7239 14603
rect 7389 14569 7423 14603
rect 19625 14569 19659 14603
rect 22109 14569 22143 14603
rect 25973 14569 26007 14603
rect 8493 14501 8527 14535
rect 9229 14501 9263 14535
rect 18061 14501 18095 14535
rect 17325 14433 17359 14467
rect 24593 14433 24627 14467
rect 31401 14433 31435 14467
rect 31861 14433 31895 14467
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 6101 14365 6135 14399
rect 6377 14365 6411 14399
rect 12817 14365 12851 14399
rect 12909 14365 12943 14399
rect 15577 14365 15611 14399
rect 17785 14365 17819 14399
rect 18061 14365 18095 14399
rect 20729 14365 20763 14399
rect 20996 14365 21030 14399
rect 24860 14365 24894 14399
rect 26433 14365 26467 14399
rect 28273 14365 28307 14399
rect 28549 14365 28583 14399
rect 31125 14365 31159 14399
rect 32137 14365 32171 14399
rect 2973 14297 3007 14331
rect 7021 14297 7055 14331
rect 7237 14297 7271 14331
rect 7941 14297 7975 14331
rect 8217 14297 8251 14331
rect 9505 14297 9539 14331
rect 9781 14297 9815 14331
rect 13093 14297 13127 14331
rect 19441 14297 19475 14331
rect 19625 14297 19659 14331
rect 26700 14297 26734 14331
rect 28733 14297 28767 14331
rect 29745 14297 29779 14331
rect 6561 14229 6595 14263
rect 8033 14229 8067 14263
rect 9689 14229 9723 14263
rect 19809 14229 19843 14263
rect 27813 14229 27847 14263
rect 28365 14229 28399 14263
rect 33241 14229 33275 14263
rect 2605 14025 2639 14059
rect 5917 14025 5951 14059
rect 16957 14025 16991 14059
rect 21097 14025 21131 14059
rect 22017 14025 22051 14059
rect 24685 14025 24719 14059
rect 25053 14025 25087 14059
rect 28917 14025 28951 14059
rect 29101 14025 29135 14059
rect 30113 14025 30147 14059
rect 31401 14025 31435 14059
rect 33701 14025 33735 14059
rect 4445 13957 4479 13991
rect 6561 13957 6595 13991
rect 6745 13957 6779 13991
rect 12081 13957 12115 13991
rect 19073 13957 19107 13991
rect 19984 13957 20018 13991
rect 27721 13957 27755 13991
rect 28733 13957 28767 13991
rect 2697 13889 2731 13923
rect 9505 13889 9539 13923
rect 9781 13889 9815 13923
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 15393 13889 15427 13923
rect 16313 13889 16347 13923
rect 16865 13889 16899 13923
rect 17417 13889 17451 13923
rect 18797 13889 18831 13923
rect 19717 13889 19751 13923
rect 22201 13889 22235 13923
rect 22293 13889 22327 13923
rect 22385 13889 22419 13923
rect 22569 13889 22603 13923
rect 23305 13889 23339 13923
rect 24593 13889 24627 13923
rect 24869 13889 24903 13923
rect 27491 13889 27525 13923
rect 27629 13889 27663 13923
rect 27813 13895 27847 13929
rect 29653 13889 29687 13923
rect 29745 13889 29779 13923
rect 29929 13889 29963 13923
rect 31309 13889 31343 13923
rect 31585 13889 31619 13923
rect 31769 13889 31803 13923
rect 32597 13889 32631 13923
rect 4169 13821 4203 13855
rect 9873 13821 9907 13855
rect 11805 13821 11839 13855
rect 14105 13821 14139 13855
rect 27353 13821 27387 13855
rect 27997 13821 28031 13855
rect 32321 13821 32355 13855
rect 6929 13753 6963 13787
rect 16037 13753 16071 13787
rect 6745 13685 6779 13719
rect 13553 13685 13587 13719
rect 23121 13685 23155 13719
rect 28917 13685 28951 13719
rect 3433 13481 3467 13515
rect 5549 13481 5583 13515
rect 15669 13481 15703 13515
rect 27353 13481 27387 13515
rect 31677 13481 31711 13515
rect 9413 13345 9447 13379
rect 16773 13345 16807 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 2973 13277 3007 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 4629 13277 4663 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 9137 13277 9171 13311
rect 11805 13277 11839 13311
rect 15025 13277 15059 13311
rect 15485 13277 15519 13311
rect 16405 13277 16439 13311
rect 17693 13277 17727 13311
rect 18245 13277 18279 13311
rect 20269 13277 20303 13311
rect 26065 13277 26099 13311
rect 32965 13277 32999 13311
rect 4261 13209 4295 13243
rect 8585 13209 8619 13243
rect 12081 13209 12115 13243
rect 16221 13209 16255 13243
rect 18429 13209 18463 13243
rect 2421 13141 2455 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 21557 13141 21591 13175
rect 3893 12937 3927 12971
rect 4353 12937 4387 12971
rect 22937 12937 22971 12971
rect 27905 12937 27939 12971
rect 32321 12937 32355 12971
rect 32689 12937 32723 12971
rect 13001 12869 13035 12903
rect 14749 12869 14783 12903
rect 19165 12869 19199 12903
rect 22569 12869 22603 12903
rect 22661 12869 22695 12903
rect 27629 12869 27663 12903
rect 2145 12801 2179 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 9597 12801 9631 12835
rect 15393 12801 15427 12835
rect 16037 12801 16071 12835
rect 17601 12801 17635 12835
rect 18061 12801 18095 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19973 12801 20007 12835
rect 22293 12801 22327 12835
rect 22386 12801 22420 12835
rect 22758 12801 22792 12835
rect 27261 12801 27295 12835
rect 27409 12801 27443 12835
rect 27537 12801 27571 12835
rect 27726 12801 27760 12835
rect 28549 12801 28583 12835
rect 28733 12801 28767 12835
rect 28825 12801 28859 12835
rect 29745 12801 29779 12835
rect 32505 12801 32539 12835
rect 32781 12801 32815 12835
rect 2421 12733 2455 12767
rect 9321 12733 9355 12767
rect 16129 12733 16163 12767
rect 18337 12733 18371 12767
rect 19717 12733 19751 12767
rect 29561 12733 29595 12767
rect 7849 12597 7883 12631
rect 21097 12597 21131 12631
rect 28365 12597 28399 12631
rect 3065 12393 3099 12427
rect 19901 12393 19935 12427
rect 22109 12393 22143 12427
rect 23029 12325 23063 12359
rect 27997 12325 28031 12359
rect 16681 12257 16715 12291
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 14565 12189 14599 12223
rect 15209 12189 15243 12223
rect 15945 12189 15979 12223
rect 16773 12189 16807 12223
rect 17509 12189 17543 12223
rect 17969 12189 18003 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 19717 12189 19751 12223
rect 23213 12189 23247 12223
rect 23305 12189 23339 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 28176 12189 28210 12223
rect 28548 12189 28582 12223
rect 28641 12189 28675 12223
rect 15025 12121 15059 12155
rect 18245 12121 18279 12155
rect 20821 12121 20855 12155
rect 28273 12121 28307 12155
rect 28365 12121 28399 12155
rect 24593 12053 24627 12087
rect 24961 12053 24995 12087
rect 22385 11849 22419 11883
rect 25237 11849 25271 11883
rect 25881 11849 25915 11883
rect 28733 11849 28767 11883
rect 31217 11849 31251 11883
rect 32689 11849 32723 11883
rect 15761 11781 15795 11815
rect 16313 11781 16347 11815
rect 22753 11781 22787 11815
rect 24124 11781 24158 11815
rect 25697 11781 25731 11815
rect 27620 11781 27654 11815
rect 14197 11713 14231 11747
rect 14565 11713 14599 11747
rect 14749 11713 14783 11747
rect 15945 11713 15979 11747
rect 17509 11713 17543 11747
rect 18061 11713 18095 11747
rect 20352 11713 20386 11747
rect 22569 11713 22603 11747
rect 22661 11713 22695 11747
rect 22937 11713 22971 11747
rect 31125 11713 31159 11747
rect 31401 11713 31435 11747
rect 32505 11713 32539 11747
rect 32781 11713 32815 11747
rect 18245 11645 18279 11679
rect 20085 11645 20119 11679
rect 23857 11645 23891 11679
rect 27353 11645 27387 11679
rect 21465 11577 21499 11611
rect 31585 11577 31619 11611
rect 25881 11509 25915 11543
rect 26065 11509 26099 11543
rect 32321 11509 32355 11543
rect 4169 11305 4203 11339
rect 20545 11305 20579 11339
rect 21005 11305 21039 11339
rect 31401 11305 31435 11339
rect 17877 11237 17911 11271
rect 5549 11101 5583 11135
rect 10333 11101 10367 11135
rect 12725 11101 12759 11135
rect 13093 11101 13127 11135
rect 13475 11101 13509 11135
rect 16957 11101 16991 11135
rect 17141 11101 17175 11135
rect 17601 11101 17635 11135
rect 17877 11101 17911 11135
rect 19901 11101 19935 11135
rect 19994 11101 20028 11135
rect 20177 11101 20211 11135
rect 20269 11101 20303 11135
rect 20366 11101 20400 11135
rect 21189 11101 21223 11135
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 23765 11101 23799 11135
rect 23949 11101 23983 11135
rect 24041 11101 24075 11135
rect 26065 11101 26099 11135
rect 29929 11101 29963 11135
rect 30205 11101 30239 11135
rect 32781 11101 32815 11135
rect 3985 11033 4019 11067
rect 4201 11033 4235 11067
rect 5816 11033 5850 11067
rect 10600 11033 10634 11067
rect 12633 11033 12667 11067
rect 16773 11033 16807 11067
rect 23581 11033 23615 11067
rect 32514 11033 32548 11067
rect 4353 10965 4387 10999
rect 6929 10965 6963 10999
rect 11713 10965 11747 10999
rect 12357 10965 12391 10999
rect 13645 10965 13679 10999
rect 27353 10965 27387 10999
rect 29745 10965 29779 10999
rect 30113 10965 30147 10999
rect 7941 10761 7975 10795
rect 9965 10761 9999 10795
rect 13645 10761 13679 10795
rect 25973 10761 26007 10795
rect 28733 10761 28767 10795
rect 33701 10761 33735 10795
rect 6837 10693 6871 10727
rect 7113 10693 7147 10727
rect 7205 10693 7239 10727
rect 7573 10693 7607 10727
rect 8861 10693 8895 10727
rect 9597 10693 9631 10727
rect 12541 10693 12575 10727
rect 12909 10693 12943 10727
rect 13277 10693 13311 10727
rect 18245 10693 18279 10727
rect 19993 10693 20027 10727
rect 24860 10693 24894 10727
rect 27620 10693 27654 10727
rect 29377 10693 29411 10727
rect 29561 10693 29595 10727
rect 3249 10625 3283 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 12817 10625 12851 10659
rect 32577 10625 32611 10659
rect 3065 10557 3099 10591
rect 3157 10557 3191 10591
rect 3341 10557 3375 10591
rect 4077 10557 4111 10591
rect 24593 10557 24627 10591
rect 27353 10557 27387 10591
rect 32321 10557 32355 10591
rect 3525 10489 3559 10523
rect 8125 10421 8159 10455
rect 10149 10421 10183 10455
rect 13829 10421 13863 10455
rect 29561 10421 29595 10455
rect 29745 10421 29779 10455
rect 4169 10217 4203 10251
rect 6745 10217 6779 10251
rect 8585 10217 8619 10251
rect 12633 10217 12667 10251
rect 21281 10217 21315 10251
rect 24961 10217 24995 10251
rect 27353 10217 27387 10251
rect 28273 10217 28307 10251
rect 32505 10217 32539 10251
rect 2145 10149 2179 10183
rect 29745 10149 29779 10183
rect 2881 10081 2915 10115
rect 7205 10081 7239 10115
rect 11253 10081 11287 10115
rect 2237 10013 2271 10047
rect 2697 10013 2731 10047
rect 2973 10013 3007 10047
rect 3341 10013 3375 10047
rect 5365 10013 5399 10047
rect 11520 10013 11554 10047
rect 22569 10013 22603 10047
rect 25140 10013 25174 10047
rect 25329 10013 25363 10047
rect 25512 10013 25546 10047
rect 25605 10013 25639 10047
rect 26065 10013 26099 10047
rect 28411 10013 28445 10047
rect 28641 10013 28675 10047
rect 28824 10013 28858 10047
rect 28917 10013 28951 10047
rect 29929 10013 29963 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 33425 10013 33459 10047
rect 33701 10013 33735 10047
rect 3985 9945 4019 9979
rect 4201 9945 4235 9979
rect 5632 9945 5666 9979
rect 7472 9945 7506 9979
rect 25237 9945 25271 9979
rect 28549 9945 28583 9979
rect 30021 9945 30055 9979
rect 31217 9945 31251 9979
rect 3065 9877 3099 9911
rect 3249 9877 3283 9911
rect 4353 9877 4387 9911
rect 33517 9877 33551 9911
rect 33885 9877 33919 9911
rect 5197 9673 5231 9707
rect 8585 9673 8619 9707
rect 27721 9673 27755 9707
rect 1961 9605 1995 9639
rect 4169 9605 4203 9639
rect 4997 9605 5031 9639
rect 11980 9605 12014 9639
rect 17233 9605 17267 9639
rect 21005 9605 21039 9639
rect 22385 9605 22419 9639
rect 27353 9605 27387 9639
rect 32413 9605 32447 9639
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 2421 9537 2455 9571
rect 3249 9537 3283 9571
rect 4077 9537 4111 9571
rect 4353 9537 4387 9571
rect 4537 9537 4571 9571
rect 7205 9537 7239 9571
rect 7472 9537 7506 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 19441 9537 19475 9571
rect 19625 9537 19659 9571
rect 19717 9537 19751 9571
rect 19809 9537 19843 9571
rect 20637 9537 20671 9571
rect 20730 9537 20764 9571
rect 20913 9537 20947 9571
rect 21102 9537 21136 9571
rect 22201 9537 22235 9571
rect 22477 9537 22511 9571
rect 27169 9537 27203 9571
rect 27445 9537 27479 9571
rect 27537 9537 27571 9571
rect 31312 9537 31346 9571
rect 31401 9537 31435 9571
rect 31539 9537 31573 9571
rect 3341 9469 3375 9503
rect 3433 9469 3467 9503
rect 11713 9469 11747 9503
rect 5365 9401 5399 9435
rect 13093 9401 13127 9435
rect 19993 9401 20027 9435
rect 33701 9401 33735 9435
rect 2881 9333 2915 9367
rect 5181 9333 5215 9367
rect 16865 9333 16899 9367
rect 21281 9333 21315 9367
rect 22017 9333 22051 9367
rect 31769 9333 31803 9367
rect 2789 9129 2823 9163
rect 2973 9129 3007 9163
rect 12173 9129 12207 9163
rect 15577 9129 15611 9163
rect 18889 9129 18923 9163
rect 21281 9129 21315 9163
rect 33701 9129 33735 9163
rect 3985 8993 4019 9027
rect 10793 8993 10827 9027
rect 3341 8925 3375 8959
rect 4169 8925 4203 8959
rect 16701 8925 16735 8959
rect 16957 8925 16991 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 17877 8925 17911 8959
rect 18337 8925 18371 8959
rect 18705 8925 18739 8959
rect 19901 8925 19935 8959
rect 20168 8925 20202 8959
rect 24593 8925 24627 8959
rect 24869 8925 24903 8959
rect 28917 8925 28951 8959
rect 29193 8925 29227 8959
rect 32321 8925 32355 8959
rect 32588 8925 32622 8959
rect 2927 8857 2961 8891
rect 11060 8857 11094 8891
rect 18521 8857 18555 8891
rect 18613 8857 18647 8891
rect 4353 8789 4387 8823
rect 24685 8789 24719 8823
rect 25053 8789 25087 8823
rect 28733 8789 28767 8823
rect 29101 8789 29135 8823
rect 3433 8585 3467 8619
rect 4077 8585 4111 8619
rect 16221 8585 16255 8619
rect 21005 8585 21039 8619
rect 23673 8585 23707 8619
rect 25881 8585 25915 8619
rect 33701 8585 33735 8619
rect 9597 8517 9631 8551
rect 15209 8517 15243 8551
rect 15393 8517 15427 8551
rect 18245 8517 18279 8551
rect 19993 8517 20027 8551
rect 20637 8517 20671 8551
rect 22753 8517 22787 8551
rect 22937 8517 22971 8551
rect 30573 8517 30607 8551
rect 32566 8517 32600 8551
rect 3525 8449 3559 8483
rect 3985 8449 4019 8483
rect 16037 8449 16071 8483
rect 16313 8449 16347 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 20453 8449 20487 8483
rect 20729 8449 20763 8483
rect 20821 8449 20855 8483
rect 24797 8449 24831 8483
rect 25053 8449 25087 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 28621 8449 28655 8483
rect 30205 8449 30239 8483
rect 30389 8449 30423 8483
rect 30665 8449 30699 8483
rect 28365 8381 28399 8415
rect 32321 8381 32355 8415
rect 15025 8313 15059 8347
rect 15853 8313 15887 8347
rect 17325 8313 17359 8347
rect 23121 8313 23155 8347
rect 25513 8313 25547 8347
rect 29745 8313 29779 8347
rect 8125 8245 8159 8279
rect 15209 8245 15243 8279
rect 22937 8245 22971 8279
rect 16957 8041 16991 8075
rect 23765 8041 23799 8075
rect 29929 8041 29963 8075
rect 32505 8041 32539 8075
rect 25881 7973 25915 8007
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 18613 7837 18647 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 22385 7837 22419 7871
rect 24593 7837 24627 7871
rect 31217 7837 31251 7871
rect 7389 7769 7423 7803
rect 10149 7769 10183 7803
rect 15669 7769 15703 7803
rect 18429 7769 18463 7803
rect 20177 7769 20211 7803
rect 22652 7769 22686 7803
rect 28549 7769 28583 7803
rect 29745 7769 29779 7803
rect 29929 7769 29963 7803
rect 21465 7701 21499 7735
rect 27261 7701 27295 7735
rect 30113 7701 30147 7735
rect 14933 7497 14967 7531
rect 20545 7497 20579 7531
rect 20729 7497 20763 7531
rect 22569 7497 22603 7531
rect 22937 7497 22971 7531
rect 24685 7497 24719 7531
rect 25973 7497 26007 7531
rect 27813 7497 27847 7531
rect 28181 7497 28215 7531
rect 6837 7429 6871 7463
rect 11958 7429 11992 7463
rect 16068 7429 16102 7463
rect 18245 7429 18279 7463
rect 19993 7429 20027 7463
rect 20913 7429 20947 7463
rect 23397 7429 23431 7463
rect 30573 7429 30607 7463
rect 2513 7361 2547 7395
rect 13553 7361 13587 7395
rect 13737 7361 13771 7395
rect 16313 7361 16347 7395
rect 22477 7361 22511 7395
rect 22753 7361 22787 7395
rect 25789 7361 25823 7395
rect 26065 7361 26099 7395
rect 27721 7361 27755 7395
rect 27997 7361 28031 7395
rect 6561 7293 6595 7327
rect 8953 7293 8987 7327
rect 9229 7293 9263 7327
rect 11713 7293 11747 7327
rect 28825 7293 28859 7327
rect 13553 7225 13587 7259
rect 2605 7157 2639 7191
rect 8309 7157 8343 7191
rect 10701 7157 10735 7191
rect 13093 7157 13127 7191
rect 20729 7157 20763 7191
rect 25605 7157 25639 7191
rect 1685 6953 1719 6987
rect 3169 6953 3203 6987
rect 27813 6885 27847 6919
rect 3433 6817 3467 6851
rect 7849 6817 7883 6851
rect 10149 6817 10183 6851
rect 10701 6817 10735 6851
rect 12265 6817 12299 6851
rect 5457 6749 5491 6783
rect 5724 6749 5758 6783
rect 7665 6749 7699 6783
rect 10241 6749 10275 6783
rect 10563 6749 10597 6783
rect 12357 6749 12391 6783
rect 15301 6749 15335 6783
rect 19441 6749 19475 6783
rect 19708 6749 19742 6783
rect 21465 6749 21499 6783
rect 21741 6749 21775 6783
rect 23765 6749 23799 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 24593 6749 24627 6783
rect 24860 6749 24894 6783
rect 29193 6749 29227 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 30205 6749 30239 6783
rect 7757 6681 7791 6715
rect 12449 6681 12483 6715
rect 21649 6681 21683 6715
rect 28948 6681 28982 6715
rect 29745 6681 29779 6715
rect 6837 6613 6871 6647
rect 7297 6613 7331 6647
rect 10977 6613 11011 6647
rect 12817 6613 12851 6647
rect 16589 6613 16623 6647
rect 20821 6613 20855 6647
rect 21281 6613 21315 6647
rect 23581 6613 23615 6647
rect 25973 6613 26007 6647
rect 6929 6409 6963 6443
rect 12909 6409 12943 6443
rect 13001 6409 13035 6443
rect 16313 6409 16347 6443
rect 20913 6409 20947 6443
rect 30021 6409 30055 6443
rect 2789 6341 2823 6375
rect 3709 6341 3743 6375
rect 6837 6341 6871 6375
rect 15200 6341 15234 6375
rect 19800 6341 19834 6375
rect 24694 6341 24728 6375
rect 28908 6341 28942 6375
rect 2973 6273 3007 6307
rect 3157 6273 3191 6307
rect 28641 6273 28675 6307
rect 6653 6205 6687 6239
rect 12725 6205 12759 6239
rect 14933 6205 14967 6239
rect 19533 6205 19567 6239
rect 24961 6205 24995 6239
rect 7297 6137 7331 6171
rect 23581 6137 23615 6171
rect 3801 6069 3835 6103
rect 13369 6069 13403 6103
rect 25973 5865 26007 5899
rect 16957 5797 16991 5831
rect 3985 5729 4019 5763
rect 4353 5729 4387 5763
rect 5825 5729 5859 5763
rect 14565 5729 14599 5763
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 15577 5661 15611 5695
rect 24593 5661 24627 5695
rect 24860 5661 24894 5695
rect 15844 5593 15878 5627
rect 14565 5525 14599 5559
rect 9597 5321 9631 5355
rect 10517 5321 10551 5355
rect 13461 5321 13495 5355
rect 19533 5321 19567 5355
rect 24685 5321 24719 5355
rect 29745 5321 29779 5355
rect 4353 5253 4387 5287
rect 9505 5253 9539 5287
rect 14749 5253 14783 5287
rect 18245 5253 18279 5287
rect 23397 5253 23431 5287
rect 28632 5253 28666 5287
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 5825 5185 5859 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 15209 5185 15243 5219
rect 25789 5185 25823 5219
rect 25973 5185 26007 5219
rect 5917 5117 5951 5151
rect 9321 5117 9355 5151
rect 28365 5117 28399 5151
rect 9965 4981 9999 5015
rect 15301 4981 15335 5015
rect 25605 4981 25639 5015
rect 13093 4709 13127 4743
rect 14565 4709 14599 4743
rect 24685 4709 24719 4743
rect 7205 4641 7239 4675
rect 9137 4641 9171 4675
rect 9413 4641 9447 4675
rect 16221 4641 16255 4675
rect 18705 4641 18739 4675
rect 20453 4641 20487 4675
rect 25053 4641 25087 4675
rect 7472 4573 7506 4607
rect 11713 4573 11747 4607
rect 11980 4573 12014 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 17417 4573 17451 4607
rect 18429 4573 18463 4607
rect 20177 4573 20211 4607
rect 21649 4573 21683 4607
rect 22293 4573 22327 4607
rect 26065 4573 26099 4607
rect 15945 4505 15979 4539
rect 26332 4505 26366 4539
rect 8585 4437 8619 4471
rect 10885 4437 10919 4471
rect 14381 4437 14415 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 17509 4437 17543 4471
rect 18061 4437 18095 4471
rect 18521 4437 18555 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 21557 4437 21591 4471
rect 22201 4437 22235 4471
rect 24593 4437 24627 4471
rect 27445 4437 27479 4471
rect 9321 4233 9355 4267
rect 9689 4233 9723 4267
rect 26157 4233 26191 4267
rect 7389 4165 7423 4199
rect 13369 4165 13403 4199
rect 17960 4165 17994 4199
rect 9781 4097 9815 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 11897 4097 11931 4131
rect 12265 4097 12299 4131
rect 13461 4097 13495 4131
rect 14933 4097 14967 4131
rect 15200 4097 15234 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 21198 4097 21232 4131
rect 21465 4097 21499 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 24584 4097 24618 4131
rect 27169 4097 27203 4131
rect 27436 4097 27470 4131
rect 7113 4029 7147 4063
rect 8861 4029 8895 4063
rect 9873 4029 9907 4063
rect 13645 4029 13679 4063
rect 24317 4029 24351 4063
rect 26617 4029 26651 4063
rect 12449 3961 12483 3995
rect 26249 3961 26283 3995
rect 11989 3893 12023 3927
rect 13001 3893 13035 3927
rect 16313 3893 16347 3927
rect 16957 3893 16991 3927
rect 19073 3893 19107 3927
rect 20085 3893 20119 3927
rect 23397 3893 23431 3927
rect 25697 3893 25731 3927
rect 28549 3893 28583 3927
rect 7941 3689 7975 3723
rect 20821 3689 20855 3723
rect 22109 3689 22143 3723
rect 24593 3689 24627 3723
rect 26801 3689 26835 3723
rect 26893 3621 26927 3655
rect 16681 3553 16715 3587
rect 22753 3553 22787 3587
rect 25973 3553 26007 3587
rect 26985 3553 27019 3587
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 12357 3485 12391 3519
rect 12624 3485 12658 3519
rect 15669 3485 15703 3519
rect 19441 3485 19475 3519
rect 19708 3485 19742 3519
rect 22477 3485 22511 3519
rect 22569 3485 22603 3519
rect 25706 3485 25740 3519
rect 26433 3485 26467 3519
rect 15402 3417 15436 3451
rect 16948 3417 16982 3451
rect 27353 3417 27387 3451
rect 13737 3349 13771 3383
rect 14289 3349 14323 3383
rect 18061 3349 18095 3383
rect 12541 3145 12575 3179
rect 14749 3145 14783 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 17417 3145 17451 3179
rect 19625 3145 19659 3179
rect 20729 3145 20763 3179
rect 21097 3145 21131 3179
rect 27629 3145 27663 3179
rect 29929 3145 29963 3179
rect 27169 3077 27203 3111
rect 28641 3077 28675 3111
rect 12633 3009 12667 3043
rect 14381 3009 14415 3043
rect 15209 3009 15243 3043
rect 17325 3009 17359 3043
rect 19717 3009 19751 3043
rect 20913 3009 20947 3043
rect 21189 3009 21223 3043
rect 25145 3009 25179 3043
rect 14197 2941 14231 2975
rect 14289 2941 14323 2975
rect 17601 2941 17635 2975
rect 25513 2941 25547 2975
rect 25605 2873 25639 2907
rect 26065 2873 26099 2907
rect 27445 2873 27479 2907
rect 25697 2805 25731 2839
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4445 2397 4479 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 11713 2397 11747 2431
rect 12909 2397 12943 2431
rect 14289 2397 14323 2431
rect 15485 2397 15519 2431
rect 16865 2397 16899 2431
rect 18061 2397 18095 2431
rect 19441 2397 19475 2431
rect 20637 2397 20671 2431
rect 22017 2397 22051 2431
rect 23213 2397 23247 2431
rect 25053 2397 25087 2431
rect 26249 2397 26283 2431
rect 27169 2397 27203 2431
rect 28365 2397 28399 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33517 2397 33551 2431
rect 1777 2329 1811 2363
rect 2789 2329 2823 2363
rect 4169 2329 4203 2363
rect 5365 2329 5399 2363
rect 14565 2329 14599 2363
rect 15761 2329 15795 2363
rect 17141 2329 17175 2363
rect 18337 2329 18371 2363
rect 19717 2329 19751 2363
rect 20913 2329 20947 2363
rect 22293 2329 22327 2363
rect 23489 2329 23523 2363
rect 24777 2329 24811 2363
rect 25973 2329 26007 2363
rect 27445 2329 27479 2363
rect 28641 2329 28675 2363
rect 34345 2261 34379 2295
<< metal1 >>
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 4890 33532 4896 33584
rect 4948 33532 4954 33584
rect 7834 33532 7840 33584
rect 7892 33532 7898 33584
rect 10594 33532 10600 33584
rect 10652 33572 10658 33584
rect 10781 33575 10839 33581
rect 10781 33572 10793 33575
rect 10652 33544 10793 33572
rect 10652 33532 10658 33544
rect 10781 33541 10793 33544
rect 10827 33541 10839 33575
rect 10781 33535 10839 33541
rect 13814 33532 13820 33584
rect 13872 33572 13878 33584
rect 14461 33575 14519 33581
rect 14461 33572 14473 33575
rect 13872 33544 14473 33572
rect 13872 33532 13878 33544
rect 14461 33541 14473 33544
rect 14507 33541 14519 33575
rect 14461 33535 14519 33541
rect 16574 33532 16580 33584
rect 16632 33572 16638 33584
rect 17037 33575 17095 33581
rect 17037 33572 17049 33575
rect 16632 33544 17049 33572
rect 16632 33532 16638 33544
rect 17037 33541 17049 33544
rect 17083 33541 17095 33575
rect 17037 33535 17095 33541
rect 19426 33532 19432 33584
rect 19484 33572 19490 33584
rect 19705 33575 19763 33581
rect 19705 33572 19717 33575
rect 19484 33544 19717 33572
rect 19484 33532 19490 33544
rect 19705 33541 19717 33544
rect 19751 33541 19763 33575
rect 19705 33535 19763 33541
rect 22370 33532 22376 33584
rect 22428 33572 22434 33584
rect 22649 33575 22707 33581
rect 22649 33572 22661 33575
rect 22428 33544 22661 33572
rect 22428 33532 22434 33544
rect 22649 33541 22661 33544
rect 22695 33541 22707 33575
rect 22649 33535 22707 33541
rect 25590 33532 25596 33584
rect 25648 33532 25654 33584
rect 28534 33532 28540 33584
rect 28592 33532 28598 33584
rect 31478 33532 31484 33584
rect 31536 33532 31542 33584
rect 34238 33532 34244 33584
rect 34296 33532 34302 33584
rect 10965 33371 11023 33377
rect 10965 33337 10977 33371
rect 11011 33368 11023 33371
rect 12250 33368 12256 33380
rect 11011 33340 12256 33368
rect 11011 33337 11023 33340
rect 10965 33331 11023 33337
rect 12250 33328 12256 33340
rect 12308 33328 12314 33380
rect 14274 33328 14280 33380
rect 14332 33328 14338 33380
rect 16850 33328 16856 33380
rect 16908 33328 16914 33380
rect 19518 33328 19524 33380
rect 19576 33328 19582 33380
rect 22462 33328 22468 33380
rect 22520 33328 22526 33380
rect 25406 33328 25412 33380
rect 25464 33328 25470 33380
rect 28350 33328 28356 33380
rect 28408 33328 28414 33380
rect 31294 33328 31300 33380
rect 31352 33328 31358 33380
rect 33318 33328 33324 33380
rect 33376 33368 33382 33380
rect 34057 33371 34115 33377
rect 34057 33368 34069 33371
rect 33376 33340 34069 33368
rect 33376 33328 33382 33340
rect 34057 33337 34069 33340
rect 34103 33337 34115 33371
rect 34057 33331 34115 33337
rect 4982 33260 4988 33312
rect 5040 33260 5046 33312
rect 7929 33303 7987 33309
rect 7929 33269 7941 33303
rect 7975 33300 7987 33303
rect 11606 33300 11612 33312
rect 7975 33272 11612 33300
rect 7975 33269 7987 33272
rect 7929 33263 7987 33269
rect 11606 33260 11612 33272
rect 11664 33260 11670 33312
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 28350 33096 28356 33108
rect 20364 33068 28356 33096
rect 16850 32960 16856 32972
rect 16500 32932 16856 32960
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32892 10287 32895
rect 10502 32892 10508 32904
rect 10275 32864 10508 32892
rect 10275 32861 10287 32864
rect 10229 32855 10287 32861
rect 10502 32852 10508 32864
rect 10560 32852 10566 32904
rect 16500 32901 16528 32932
rect 16850 32920 16856 32932
rect 16908 32920 16914 32972
rect 16301 32895 16359 32901
rect 16301 32861 16313 32895
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32892 16635 32895
rect 20364 32892 20392 33068
rect 28350 33056 28356 33068
rect 28408 33056 28414 33108
rect 20622 32920 20628 32972
rect 20680 32920 20686 32972
rect 24762 32960 24768 32972
rect 21928 32932 24768 32960
rect 16623 32864 20392 32892
rect 20533 32895 20591 32901
rect 16623 32861 16635 32864
rect 16577 32855 16635 32861
rect 20533 32861 20545 32895
rect 20579 32892 20591 32895
rect 21928 32892 21956 32932
rect 24762 32920 24768 32932
rect 24820 32920 24826 32972
rect 20579 32864 21956 32892
rect 22373 32895 22431 32901
rect 20579 32861 20591 32864
rect 20533 32855 20591 32861
rect 22373 32861 22385 32895
rect 22419 32892 22431 32895
rect 22830 32892 22836 32904
rect 22419 32864 22836 32892
rect 22419 32861 22431 32864
rect 22373 32855 22431 32861
rect 15470 32784 15476 32836
rect 15528 32824 15534 32836
rect 15841 32827 15899 32833
rect 15841 32824 15853 32827
rect 15528 32796 15853 32824
rect 15528 32784 15534 32796
rect 15841 32793 15853 32796
rect 15887 32793 15899 32827
rect 16316 32824 16344 32855
rect 16758 32824 16764 32836
rect 16316 32796 16764 32824
rect 15841 32787 15899 32793
rect 16758 32784 16764 32796
rect 16816 32784 16822 32836
rect 18322 32784 18328 32836
rect 18380 32824 18386 32836
rect 20548 32824 20576 32855
rect 22830 32852 22836 32864
rect 22888 32852 22894 32904
rect 25406 32824 25412 32836
rect 18380 32796 20576 32824
rect 20824 32796 25412 32824
rect 18380 32784 18386 32796
rect 10134 32716 10140 32768
rect 10192 32716 10198 32768
rect 13262 32716 13268 32768
rect 13320 32756 13326 32768
rect 20824 32756 20852 32796
rect 25406 32784 25412 32796
rect 25464 32784 25470 32836
rect 13320 32728 20852 32756
rect 20901 32759 20959 32765
rect 13320 32716 13326 32728
rect 20901 32725 20913 32759
rect 20947 32756 20959 32759
rect 21266 32756 21272 32768
rect 20947 32728 21272 32756
rect 20947 32725 20959 32728
rect 20901 32719 20959 32725
rect 21266 32716 21272 32728
rect 21324 32716 21330 32768
rect 22002 32716 22008 32768
rect 22060 32756 22066 32768
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 22060 32728 22293 32756
rect 22060 32716 22066 32728
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 22281 32719 22339 32725
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 12250 32512 12256 32564
rect 12308 32512 12314 32564
rect 13449 32555 13507 32561
rect 12360 32524 13400 32552
rect 11790 32444 11796 32496
rect 11848 32484 11854 32496
rect 12360 32493 12388 32524
rect 12345 32487 12403 32493
rect 12345 32484 12357 32487
rect 11848 32456 12357 32484
rect 11848 32444 11854 32456
rect 12345 32453 12357 32456
rect 12391 32453 12403 32487
rect 12345 32447 12403 32453
rect 13262 32444 13268 32496
rect 13320 32444 13326 32496
rect 13372 32484 13400 32524
rect 13449 32521 13461 32555
rect 13495 32552 13507 32555
rect 14274 32552 14280 32564
rect 13495 32524 14280 32552
rect 13495 32521 13507 32524
rect 13449 32515 13507 32521
rect 14274 32512 14280 32524
rect 14332 32512 14338 32564
rect 16758 32552 16764 32564
rect 14384 32524 16764 32552
rect 13541 32487 13599 32493
rect 13541 32484 13553 32487
rect 13372 32456 13553 32484
rect 13541 32453 13553 32456
rect 13587 32484 13599 32487
rect 14384 32484 14412 32524
rect 16758 32512 16764 32524
rect 16816 32512 16822 32564
rect 17313 32555 17371 32561
rect 17313 32521 17325 32555
rect 17359 32552 17371 32555
rect 18049 32555 18107 32561
rect 18049 32552 18061 32555
rect 17359 32524 18061 32552
rect 17359 32521 17371 32524
rect 17313 32515 17371 32521
rect 18049 32521 18061 32524
rect 18095 32521 18107 32555
rect 22462 32552 22468 32564
rect 18049 32515 18107 32521
rect 19536 32524 22468 32552
rect 19536 32484 19564 32524
rect 22462 32512 22468 32524
rect 22520 32512 22526 32564
rect 13587 32456 14412 32484
rect 14476 32456 19564 32484
rect 21177 32487 21235 32493
rect 13587 32453 13599 32456
rect 13541 32447 13599 32453
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32416 9919 32419
rect 10410 32416 10416 32428
rect 9907 32388 10416 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 10410 32376 10416 32388
rect 10468 32376 10474 32428
rect 10502 32376 10508 32428
rect 10560 32376 10566 32428
rect 12069 32419 12127 32425
rect 12069 32385 12081 32419
rect 12115 32416 12127 32419
rect 14476 32416 14504 32456
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 21223 32456 22109 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 23382 32484 23388 32496
rect 22097 32447 22155 32453
rect 23032 32456 23388 32484
rect 12115 32388 14504 32416
rect 12115 32385 12127 32388
rect 12069 32379 12127 32385
rect 15930 32376 15936 32428
rect 15988 32416 15994 32428
rect 16117 32419 16175 32425
rect 16117 32416 16129 32419
rect 15988 32388 16129 32416
rect 15988 32376 15994 32388
rect 16117 32385 16129 32388
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 16301 32419 16359 32425
rect 16301 32385 16313 32419
rect 16347 32416 16359 32419
rect 16850 32416 16856 32428
rect 16347 32388 16856 32416
rect 16347 32385 16359 32388
rect 16301 32379 16359 32385
rect 16850 32376 16856 32388
rect 16908 32376 16914 32428
rect 17221 32419 17279 32425
rect 17221 32385 17233 32419
rect 17267 32416 17279 32419
rect 17862 32416 17868 32428
rect 17267 32388 17868 32416
rect 17267 32385 17279 32388
rect 17221 32379 17279 32385
rect 17862 32376 17868 32388
rect 17920 32416 17926 32428
rect 18049 32419 18107 32425
rect 18049 32416 18061 32419
rect 17920 32388 18061 32416
rect 17920 32376 17926 32388
rect 18049 32385 18061 32388
rect 18095 32385 18107 32419
rect 18049 32379 18107 32385
rect 18230 32376 18236 32428
rect 18288 32416 18294 32428
rect 21085 32419 21143 32425
rect 18288 32388 20760 32416
rect 18288 32376 18294 32388
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32317 10747 32351
rect 10689 32311 10747 32317
rect 16209 32351 16267 32357
rect 16209 32317 16221 32351
rect 16255 32348 16267 32351
rect 17405 32351 17463 32357
rect 16255 32320 16988 32348
rect 16255 32317 16267 32320
rect 16209 32311 16267 32317
rect 8570 32240 8576 32292
rect 8628 32280 8634 32292
rect 10704 32280 10732 32311
rect 16853 32283 16911 32289
rect 16853 32280 16865 32283
rect 8628 32252 16865 32280
rect 8628 32240 8634 32252
rect 16853 32249 16865 32252
rect 16899 32249 16911 32283
rect 16960 32280 16988 32320
rect 17405 32317 17417 32351
rect 17451 32317 17463 32351
rect 17405 32311 17463 32317
rect 17420 32280 17448 32311
rect 20732 32289 20760 32388
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 22002 32416 22008 32428
rect 21131 32388 22008 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 22646 32416 22652 32428
rect 22235 32388 22652 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22646 32376 22652 32388
rect 22704 32376 22710 32428
rect 23032 32425 23060 32456
rect 23382 32444 23388 32456
rect 23440 32444 23446 32496
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 23198 32376 23204 32428
rect 23256 32376 23262 32428
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32416 24547 32419
rect 24578 32416 24584 32428
rect 24535 32388 24584 32416
rect 24535 32385 24547 32388
rect 24489 32379 24547 32385
rect 24578 32376 24584 32388
rect 24636 32376 24642 32428
rect 24673 32419 24731 32425
rect 24673 32385 24685 32419
rect 24719 32416 24731 32419
rect 24762 32416 24768 32428
rect 24719 32388 24768 32416
rect 24719 32385 24731 32388
rect 24673 32379 24731 32385
rect 24762 32376 24768 32388
rect 24820 32376 24826 32428
rect 27706 32376 27712 32428
rect 27764 32376 27770 32428
rect 28074 32376 28080 32428
rect 28132 32376 28138 32428
rect 30469 32419 30527 32425
rect 30469 32385 30481 32419
rect 30515 32416 30527 32419
rect 31294 32416 31300 32428
rect 30515 32388 31300 32416
rect 30515 32385 30527 32388
rect 30469 32379 30527 32385
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 33318 32376 33324 32428
rect 33376 32376 33382 32428
rect 21266 32308 21272 32360
rect 21324 32308 21330 32360
rect 22830 32308 22836 32360
rect 22888 32348 22894 32360
rect 27157 32351 27215 32357
rect 27157 32348 27169 32351
rect 22888 32320 27169 32348
rect 22888 32308 22894 32320
rect 27157 32317 27169 32320
rect 27203 32317 27215 32351
rect 27157 32311 27215 32317
rect 16960 32252 17448 32280
rect 20717 32283 20775 32289
rect 16853 32243 16911 32249
rect 20717 32249 20729 32283
rect 20763 32249 20775 32283
rect 20717 32243 20775 32249
rect 21082 32240 21088 32292
rect 21140 32280 21146 32292
rect 22925 32283 22983 32289
rect 22925 32280 22937 32283
rect 21140 32252 22937 32280
rect 21140 32240 21146 32252
rect 22925 32249 22937 32252
rect 22971 32249 22983 32283
rect 22925 32243 22983 32249
rect 9861 32215 9919 32221
rect 9861 32181 9873 32215
rect 9907 32212 9919 32215
rect 10042 32212 10048 32224
rect 9907 32184 10048 32212
rect 9907 32181 9919 32184
rect 9861 32175 9919 32181
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 10594 32172 10600 32224
rect 10652 32172 10658 32224
rect 11793 32215 11851 32221
rect 11793 32181 11805 32215
rect 11839 32212 11851 32215
rect 11882 32212 11888 32224
rect 11839 32184 11888 32212
rect 11839 32181 11851 32184
rect 11793 32175 11851 32181
rect 11882 32172 11888 32184
rect 11940 32172 11946 32224
rect 12989 32215 13047 32221
rect 12989 32181 13001 32215
rect 13035 32212 13047 32215
rect 13170 32212 13176 32224
rect 13035 32184 13176 32212
rect 13035 32181 13047 32184
rect 12989 32175 13047 32181
rect 13170 32172 13176 32184
rect 13228 32172 13234 32224
rect 13354 32172 13360 32224
rect 13412 32212 13418 32224
rect 19518 32212 19524 32224
rect 13412 32184 19524 32212
rect 13412 32172 13418 32184
rect 19518 32172 19524 32184
rect 19576 32172 19582 32224
rect 24581 32215 24639 32221
rect 24581 32181 24593 32215
rect 24627 32212 24639 32215
rect 25038 32212 25044 32224
rect 24627 32184 25044 32212
rect 24627 32181 24639 32184
rect 24581 32175 24639 32181
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 30190 32172 30196 32224
rect 30248 32212 30254 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 30248 32184 30297 32212
rect 30248 32172 30254 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 30285 32175 30343 32181
rect 33134 32172 33140 32224
rect 33192 32172 33198 32224
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 15749 32011 15807 32017
rect 15749 31977 15761 32011
rect 15795 32008 15807 32011
rect 15838 32008 15844 32020
rect 15795 31980 15844 32008
rect 15795 31977 15807 31980
rect 15749 31971 15807 31977
rect 15838 31968 15844 31980
rect 15896 31968 15902 32020
rect 15930 31968 15936 32020
rect 15988 31968 15994 32020
rect 18049 32011 18107 32017
rect 18049 31977 18061 32011
rect 18095 32008 18107 32011
rect 18230 32008 18236 32020
rect 18095 31980 18236 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 20622 31968 20628 32020
rect 20680 32008 20686 32020
rect 21269 32011 21327 32017
rect 21269 32008 21281 32011
rect 20680 31980 21281 32008
rect 20680 31968 20686 31980
rect 21269 31977 21281 31980
rect 21315 31977 21327 32011
rect 21269 31971 21327 31977
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 23661 32011 23719 32017
rect 23661 32008 23673 32011
rect 23256 31980 23673 32008
rect 23256 31968 23262 31980
rect 23661 31977 23673 31980
rect 23707 31977 23719 32011
rect 23661 31971 23719 31977
rect 8754 31900 8760 31952
rect 8812 31940 8818 31952
rect 9309 31943 9367 31949
rect 9309 31940 9321 31943
rect 8812 31912 9321 31940
rect 8812 31900 8818 31912
rect 9309 31909 9321 31912
rect 9355 31909 9367 31943
rect 9309 31903 9367 31909
rect 11149 31943 11207 31949
rect 11149 31909 11161 31943
rect 11195 31940 11207 31943
rect 11698 31940 11704 31952
rect 11195 31912 11704 31940
rect 11195 31909 11207 31912
rect 11149 31903 11207 31909
rect 11698 31900 11704 31912
rect 11756 31900 11762 31952
rect 15654 31940 15660 31952
rect 13464 31912 15660 31940
rect 8481 31875 8539 31881
rect 8481 31841 8493 31875
rect 8527 31872 8539 31875
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 8527 31844 9781 31872
rect 8527 31841 8539 31844
rect 8481 31835 8539 31841
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 9769 31835 9827 31841
rect 9858 31832 9864 31884
rect 9916 31832 9922 31884
rect 11609 31875 11667 31881
rect 11609 31841 11621 31875
rect 11655 31872 11667 31875
rect 13354 31872 13360 31884
rect 11655 31844 13360 31872
rect 11655 31841 11667 31844
rect 11609 31835 11667 31841
rect 13354 31832 13360 31844
rect 13412 31832 13418 31884
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31804 8447 31807
rect 8435 31776 8524 31804
rect 8435 31773 8447 31776
rect 8389 31767 8447 31773
rect 8496 31736 8524 31776
rect 8570 31764 8576 31816
rect 8628 31764 8634 31816
rect 9677 31807 9735 31813
rect 9677 31804 9689 31807
rect 8680 31776 9689 31804
rect 8680 31736 8708 31776
rect 9677 31773 9689 31776
rect 9723 31804 9735 31807
rect 10134 31804 10140 31816
rect 9723 31776 10140 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 10502 31764 10508 31816
rect 10560 31804 10566 31816
rect 13464 31813 13492 31912
rect 15654 31900 15660 31912
rect 15712 31900 15718 31952
rect 18325 31943 18383 31949
rect 18325 31909 18337 31943
rect 18371 31909 18383 31943
rect 18325 31903 18383 31909
rect 13541 31875 13599 31881
rect 13541 31841 13553 31875
rect 13587 31872 13599 31875
rect 14369 31875 14427 31881
rect 14369 31872 14381 31875
rect 13587 31844 14381 31872
rect 13587 31841 13599 31844
rect 13541 31835 13599 31841
rect 14369 31841 14381 31844
rect 14415 31841 14427 31875
rect 14369 31835 14427 31841
rect 17126 31832 17132 31884
rect 17184 31832 17190 31884
rect 18340 31872 18368 31903
rect 20530 31900 20536 31952
rect 20588 31940 20594 31952
rect 20588 31912 22048 31940
rect 20588 31900 20594 31912
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 17420 31844 18368 31872
rect 18432 31844 19441 31872
rect 12621 31807 12679 31813
rect 12621 31804 12633 31807
rect 10560 31776 12633 31804
rect 10560 31764 10566 31776
rect 12621 31773 12633 31776
rect 12667 31773 12679 31807
rect 12621 31767 12679 31773
rect 13449 31807 13507 31813
rect 13449 31773 13461 31807
rect 13495 31773 13507 31807
rect 13449 31767 13507 31773
rect 14274 31764 14280 31816
rect 14332 31764 14338 31816
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14642 31804 14648 31816
rect 14507 31776 14648 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 14642 31764 14648 31776
rect 14700 31804 14706 31816
rect 16393 31807 16451 31813
rect 16393 31804 16405 31807
rect 14700 31776 16405 31804
rect 14700 31764 14706 31776
rect 16393 31773 16405 31776
rect 16439 31773 16451 31807
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 16393 31767 16451 31773
rect 16776 31776 17233 31804
rect 8496 31708 8708 31736
rect 11606 31696 11612 31748
rect 11664 31696 11670 31748
rect 11701 31739 11759 31745
rect 11701 31705 11713 31739
rect 11747 31736 11759 31739
rect 11790 31736 11796 31748
rect 11747 31708 11796 31736
rect 11747 31705 11759 31708
rect 11701 31699 11759 31705
rect 11790 31696 11796 31708
rect 11848 31696 11854 31748
rect 15565 31739 15623 31745
rect 15565 31705 15577 31739
rect 15611 31736 15623 31739
rect 15611 31708 15884 31736
rect 15611 31705 15623 31708
rect 15565 31699 15623 31705
rect 10042 31628 10048 31680
rect 10100 31668 10106 31680
rect 15580 31668 15608 31699
rect 10100 31640 15608 31668
rect 10100 31628 10106 31640
rect 15746 31628 15752 31680
rect 15804 31677 15810 31680
rect 15804 31671 15823 31677
rect 15811 31637 15823 31671
rect 15856 31668 15884 31708
rect 15930 31696 15936 31748
rect 15988 31736 15994 31748
rect 16776 31736 16804 31776
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 17310 31764 17316 31816
rect 17368 31764 17374 31816
rect 15988 31708 16804 31736
rect 16853 31739 16911 31745
rect 15988 31696 15994 31708
rect 16853 31705 16865 31739
rect 16899 31736 16911 31739
rect 17420 31736 17448 31844
rect 17862 31764 17868 31816
rect 17920 31804 17926 31816
rect 18325 31807 18383 31813
rect 18325 31804 18337 31807
rect 17920 31776 18337 31804
rect 17920 31764 17926 31776
rect 18325 31773 18337 31776
rect 18371 31804 18383 31807
rect 18432 31804 18460 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 21082 31872 21088 31884
rect 19429 31835 19487 31841
rect 20272 31844 21088 31872
rect 20272 31813 20300 31844
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 22020 31881 22048 31912
rect 22646 31900 22652 31952
rect 22704 31940 22710 31952
rect 24581 31943 24639 31949
rect 24581 31940 24593 31943
rect 22704 31912 24593 31940
rect 22704 31900 22710 31912
rect 24581 31909 24593 31912
rect 24627 31909 24639 31943
rect 24581 31903 24639 31909
rect 22005 31875 22063 31881
rect 22005 31841 22017 31875
rect 22051 31841 22063 31875
rect 22005 31835 22063 31841
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 22664 31872 22692 31900
rect 22922 31872 22928 31884
rect 22603 31844 22692 31872
rect 22756 31844 22928 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 18371 31776 18460 31804
rect 18509 31807 18567 31813
rect 18371 31773 18383 31776
rect 18325 31767 18383 31773
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 20257 31807 20315 31813
rect 18555 31776 20208 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 16899 31708 17448 31736
rect 16899 31705 16911 31708
rect 16853 31699 16911 31705
rect 16666 31668 16672 31680
rect 15856 31640 16672 31668
rect 15804 31631 15823 31637
rect 15804 31628 15810 31631
rect 16666 31628 16672 31640
rect 16724 31668 16730 31680
rect 18322 31668 18328 31680
rect 16724 31640 18328 31668
rect 16724 31628 16730 31640
rect 18322 31628 18328 31640
rect 18380 31628 18386 31680
rect 20180 31668 20208 31776
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31804 20499 31807
rect 20806 31804 20812 31816
rect 20487 31776 20812 31804
rect 20487 31773 20499 31776
rect 20441 31767 20499 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 20993 31807 21051 31813
rect 20993 31773 21005 31807
rect 21039 31804 21051 31807
rect 21174 31804 21180 31816
rect 21039 31776 21180 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21174 31764 21180 31776
rect 21232 31764 21238 31816
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 21358 31804 21364 31816
rect 21315 31776 21364 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21358 31764 21364 31776
rect 21416 31764 21422 31816
rect 22756 31804 22784 31844
rect 22922 31832 22928 31844
rect 22980 31872 22986 31884
rect 23017 31875 23075 31881
rect 23017 31872 23029 31875
rect 22980 31844 23029 31872
rect 22980 31832 22986 31844
rect 23017 31841 23029 31844
rect 23063 31841 23075 31875
rect 23017 31835 23075 31841
rect 25038 31832 25044 31884
rect 25096 31832 25102 31884
rect 25130 31832 25136 31884
rect 25188 31832 25194 31884
rect 21468 31776 22784 31804
rect 21082 31696 21088 31748
rect 21140 31696 21146 31748
rect 21468 31668 21496 31776
rect 22830 31764 22836 31816
rect 22888 31764 22894 31816
rect 23750 31764 23756 31816
rect 23808 31764 23814 31816
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31773 26479 31807
rect 26421 31767 26479 31773
rect 23382 31696 23388 31748
rect 23440 31736 23446 31748
rect 23860 31736 23888 31767
rect 23440 31708 23888 31736
rect 26436 31736 26464 31767
rect 26602 31764 26608 31816
rect 26660 31764 26666 31816
rect 26694 31736 26700 31748
rect 26436 31708 26700 31736
rect 23440 31696 23446 31708
rect 26694 31696 26700 31708
rect 26752 31696 26758 31748
rect 27706 31736 27712 31748
rect 27554 31708 27712 31736
rect 27706 31696 27712 31708
rect 27764 31696 27770 31748
rect 20180 31640 21496 31668
rect 23474 31628 23480 31680
rect 23532 31628 23538 31680
rect 24762 31628 24768 31680
rect 24820 31668 24826 31680
rect 24949 31671 25007 31677
rect 24949 31668 24961 31671
rect 24820 31640 24961 31668
rect 24820 31628 24826 31640
rect 24949 31637 24961 31640
rect 24995 31637 25007 31671
rect 24949 31631 25007 31637
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 9493 31467 9551 31473
rect 9493 31433 9505 31467
rect 9539 31464 9551 31467
rect 9858 31464 9864 31476
rect 9539 31436 9864 31464
rect 9539 31433 9551 31436
rect 9493 31427 9551 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 14274 31464 14280 31476
rect 13587 31436 14280 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 14274 31424 14280 31436
rect 14332 31424 14338 31476
rect 15838 31424 15844 31476
rect 15896 31464 15902 31476
rect 16117 31467 16175 31473
rect 16117 31464 16129 31467
rect 15896 31436 16129 31464
rect 15896 31424 15902 31436
rect 16117 31433 16129 31436
rect 16163 31464 16175 31467
rect 17037 31467 17095 31473
rect 17037 31464 17049 31467
rect 16163 31436 17049 31464
rect 16163 31433 16175 31436
rect 16117 31427 16175 31433
rect 17037 31433 17049 31436
rect 17083 31433 17095 31467
rect 17037 31427 17095 31433
rect 17310 31424 17316 31476
rect 17368 31464 17374 31476
rect 17589 31467 17647 31473
rect 17589 31464 17601 31467
rect 17368 31436 17601 31464
rect 17368 31424 17374 31436
rect 17589 31433 17601 31436
rect 17635 31433 17647 31467
rect 17589 31427 17647 31433
rect 20806 31424 20812 31476
rect 20864 31473 20870 31476
rect 20864 31467 20892 31473
rect 20880 31433 20892 31467
rect 20864 31427 20892 31433
rect 24765 31467 24823 31473
rect 24765 31433 24777 31467
rect 24811 31464 24823 31467
rect 25130 31464 25136 31476
rect 24811 31436 25136 31464
rect 24811 31433 24823 31436
rect 24765 31427 24823 31433
rect 20864 31424 20870 31427
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 25869 31467 25927 31473
rect 25869 31433 25881 31467
rect 25915 31464 25927 31467
rect 26602 31464 26608 31476
rect 25915 31436 26608 31464
rect 25915 31433 25927 31436
rect 25869 31427 25927 31433
rect 26602 31424 26608 31436
rect 26660 31424 26666 31476
rect 27338 31424 27344 31476
rect 27396 31464 27402 31476
rect 28629 31467 28687 31473
rect 28629 31464 28641 31467
rect 27396 31436 28641 31464
rect 27396 31424 27402 31436
rect 28629 31433 28641 31436
rect 28675 31433 28687 31467
rect 28629 31427 28687 31433
rect 10042 31356 10048 31408
rect 10100 31396 10106 31408
rect 10321 31399 10379 31405
rect 10321 31396 10333 31399
rect 10100 31368 10333 31396
rect 10100 31356 10106 31368
rect 10321 31365 10333 31368
rect 10367 31365 10379 31399
rect 10321 31359 10379 31365
rect 10594 31356 10600 31408
rect 10652 31396 10658 31408
rect 10689 31399 10747 31405
rect 10689 31396 10701 31399
rect 10652 31368 10701 31396
rect 10652 31356 10658 31368
rect 10689 31365 10701 31368
rect 10735 31365 10747 31399
rect 10689 31359 10747 31365
rect 13188 31368 15608 31396
rect 8846 31288 8852 31340
rect 8904 31328 8910 31340
rect 9125 31331 9183 31337
rect 9125 31328 9137 31331
rect 8904 31300 9137 31328
rect 8904 31288 8910 31300
rect 9125 31297 9137 31300
rect 9171 31328 9183 31331
rect 9950 31328 9956 31340
rect 9171 31300 9956 31328
rect 9171 31297 9183 31300
rect 9125 31291 9183 31297
rect 9950 31288 9956 31300
rect 10008 31288 10014 31340
rect 10226 31288 10232 31340
rect 10284 31288 10290 31340
rect 12710 31288 12716 31340
rect 12768 31328 12774 31340
rect 13188 31337 13216 31368
rect 15580 31340 15608 31368
rect 15654 31356 15660 31408
rect 15712 31396 15718 31408
rect 16022 31396 16028 31408
rect 15712 31368 16028 31396
rect 15712 31356 15718 31368
rect 16022 31356 16028 31368
rect 16080 31396 16086 31408
rect 16080 31368 16344 31396
rect 16080 31356 16086 31368
rect 13173 31331 13231 31337
rect 13173 31328 13185 31331
rect 12768 31300 13185 31328
rect 12768 31288 12774 31300
rect 13173 31297 13185 31300
rect 13219 31297 13231 31331
rect 13173 31291 13231 31297
rect 14090 31288 14096 31340
rect 14148 31288 14154 31340
rect 14826 31288 14832 31340
rect 14884 31288 14890 31340
rect 14921 31331 14979 31337
rect 14921 31297 14933 31331
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9398 31260 9404 31272
rect 9263 31232 9404 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 9398 31220 9404 31232
rect 9456 31220 9462 31272
rect 9490 31220 9496 31272
rect 9548 31260 9554 31272
rect 10413 31263 10471 31269
rect 10413 31260 10425 31263
rect 9548 31232 10425 31260
rect 9548 31220 9554 31232
rect 10413 31229 10425 31232
rect 10459 31260 10471 31263
rect 12434 31260 12440 31272
rect 10459 31232 12440 31260
rect 10459 31229 10471 31232
rect 10413 31223 10471 31229
rect 12434 31220 12440 31232
rect 12492 31220 12498 31272
rect 13262 31220 13268 31272
rect 13320 31220 13326 31272
rect 14642 31220 14648 31272
rect 14700 31260 14706 31272
rect 14936 31260 14964 31291
rect 15562 31288 15568 31340
rect 15620 31328 15626 31340
rect 16316 31337 16344 31368
rect 16666 31356 16672 31408
rect 16724 31396 16730 31408
rect 16853 31399 16911 31405
rect 16853 31396 16865 31399
rect 16724 31368 16865 31396
rect 16724 31356 16730 31368
rect 16853 31365 16865 31368
rect 16899 31365 16911 31399
rect 22189 31399 22247 31405
rect 22189 31396 22201 31399
rect 16853 31359 16911 31365
rect 20640 31368 22201 31396
rect 16117 31331 16175 31337
rect 16117 31328 16129 31331
rect 15620 31300 16129 31328
rect 15620 31288 15626 31300
rect 16117 31297 16129 31300
rect 16163 31297 16175 31331
rect 16117 31291 16175 31297
rect 16301 31331 16359 31337
rect 16301 31297 16313 31331
rect 16347 31297 16359 31331
rect 16301 31291 16359 31297
rect 17126 31288 17132 31340
rect 17184 31288 17190 31340
rect 17586 31288 17592 31340
rect 17644 31288 17650 31340
rect 17678 31288 17684 31340
rect 17736 31328 17742 31340
rect 17773 31331 17831 31337
rect 17773 31328 17785 31331
rect 17736 31300 17785 31328
rect 17736 31288 17742 31300
rect 17773 31297 17785 31300
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 20640 31337 20668 31368
rect 22189 31365 22201 31368
rect 22235 31365 22247 31399
rect 24486 31396 24492 31408
rect 22189 31359 22247 31365
rect 22940 31368 24492 31396
rect 22940 31340 22968 31368
rect 24486 31356 24492 31368
rect 24544 31356 24550 31408
rect 24670 31356 24676 31408
rect 24728 31396 24734 31408
rect 24728 31368 27660 31396
rect 24728 31356 24734 31368
rect 20625 31331 20683 31337
rect 20625 31328 20637 31331
rect 20404 31300 20637 31328
rect 20404 31288 20410 31300
rect 20625 31297 20637 31300
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 21048 31300 21097 31328
rect 21048 31288 21054 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 22646 31288 22652 31340
rect 22704 31288 22710 31340
rect 22922 31288 22928 31340
rect 22980 31288 22986 31340
rect 23014 31288 23020 31340
rect 23072 31288 23078 31340
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31297 23351 31331
rect 23293 31291 23351 31297
rect 14700 31232 14964 31260
rect 14700 31220 14706 31232
rect 15746 31220 15752 31272
rect 15804 31260 15810 31272
rect 17144 31260 17172 31288
rect 21364 31272 21416 31278
rect 15804 31232 17172 31260
rect 15804 31220 15810 31232
rect 20530 31220 20536 31272
rect 20588 31220 20594 31272
rect 21450 31220 21456 31272
rect 21508 31260 21514 31272
rect 23308 31260 23336 31291
rect 23474 31288 23480 31340
rect 23532 31288 23538 31340
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31328 24271 31331
rect 24578 31328 24584 31340
rect 24259 31300 24584 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 24578 31288 24584 31300
rect 24636 31328 24642 31340
rect 24854 31328 24860 31340
rect 24636 31300 24860 31328
rect 24636 31288 24642 31300
rect 24854 31288 24860 31300
rect 24912 31288 24918 31340
rect 25240 31337 25268 31368
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25314 31288 25320 31340
rect 25372 31328 25378 31340
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25372 31300 25421 31328
rect 25372 31288 25378 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 25409 31291 25467 31297
rect 25682 31288 25688 31340
rect 25740 31288 25746 31340
rect 26694 31288 26700 31340
rect 26752 31328 26758 31340
rect 27338 31328 27344 31340
rect 26752 31300 27344 31328
rect 26752 31288 26758 31300
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27632 31337 27660 31368
rect 27617 31331 27675 31337
rect 27617 31297 27629 31331
rect 27663 31328 27675 31331
rect 28567 31331 28625 31337
rect 28567 31328 28579 31331
rect 27663 31300 28579 31328
rect 27663 31297 27675 31300
rect 27617 31291 27675 31297
rect 28567 31297 28579 31300
rect 28613 31297 28625 31331
rect 28567 31291 28625 31297
rect 21508 31232 23336 31260
rect 24489 31263 24547 31269
rect 21508 31220 21514 31232
rect 24489 31229 24501 31263
rect 24535 31260 24547 31263
rect 25590 31260 25596 31272
rect 24535 31232 25596 31260
rect 24535 31229 24547 31232
rect 24489 31223 24547 31229
rect 25590 31220 25596 31232
rect 25648 31260 25654 31272
rect 27157 31263 27215 31269
rect 27157 31260 27169 31263
rect 25648 31232 27169 31260
rect 25648 31220 25654 31232
rect 27157 31229 27169 31232
rect 27203 31229 27215 31263
rect 27157 31223 27215 31229
rect 29086 31220 29092 31272
rect 29144 31220 29150 31272
rect 21364 31214 21416 31220
rect 10686 31152 10692 31204
rect 10744 31192 10750 31204
rect 10873 31195 10931 31201
rect 10873 31192 10885 31195
rect 10744 31164 10885 31192
rect 10744 31152 10750 31164
rect 10873 31161 10885 31164
rect 10919 31161 10931 31195
rect 10873 31155 10931 31161
rect 16850 31152 16856 31204
rect 16908 31152 16914 31204
rect 25501 31195 25559 31201
rect 25501 31161 25513 31195
rect 25547 31161 25559 31195
rect 25501 31155 25559 31161
rect 14274 31084 14280 31136
rect 14332 31084 14338 31136
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 25516 31124 25544 31155
rect 25774 31124 25780 31136
rect 24627 31096 25780 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 25774 31084 25780 31096
rect 25832 31124 25838 31136
rect 28445 31127 28503 31133
rect 28445 31124 28457 31127
rect 25832 31096 28457 31124
rect 25832 31084 25838 31096
rect 28445 31093 28457 31096
rect 28491 31093 28503 31127
rect 28445 31087 28503 31093
rect 28994 31084 29000 31136
rect 29052 31084 29058 31136
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 9398 30880 9404 30932
rect 9456 30880 9462 30932
rect 10042 30880 10048 30932
rect 10100 30880 10106 30932
rect 10226 30880 10232 30932
rect 10284 30920 10290 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10284 30892 10701 30920
rect 10284 30880 10290 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 13262 30880 13268 30932
rect 13320 30920 13326 30932
rect 13541 30923 13599 30929
rect 13541 30920 13553 30923
rect 13320 30892 13553 30920
rect 13320 30880 13326 30892
rect 13541 30889 13553 30892
rect 13587 30889 13599 30923
rect 13541 30883 13599 30889
rect 20990 30880 20996 30932
rect 21048 30880 21054 30932
rect 22741 30923 22799 30929
rect 22741 30889 22753 30923
rect 22787 30920 22799 30923
rect 23014 30920 23020 30932
rect 22787 30892 23020 30920
rect 22787 30889 22799 30892
rect 22741 30883 22799 30889
rect 23014 30880 23020 30892
rect 23072 30880 23078 30932
rect 10060 30784 10088 30880
rect 14826 30852 14832 30864
rect 13464 30824 14832 30852
rect 9324 30756 10088 30784
rect 9324 30725 9352 30756
rect 10502 30744 10508 30796
rect 10560 30784 10566 30796
rect 13464 30793 13492 30824
rect 14826 30812 14832 30824
rect 14884 30852 14890 30864
rect 23109 30855 23167 30861
rect 14884 30824 16252 30852
rect 14884 30812 14890 30824
rect 13449 30787 13507 30793
rect 10560 30756 10824 30784
rect 10560 30744 10566 30756
rect 9309 30719 9367 30725
rect 9309 30685 9321 30719
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 9490 30676 9496 30728
rect 9548 30676 9554 30728
rect 9950 30676 9956 30728
rect 10008 30676 10014 30728
rect 10134 30676 10140 30728
rect 10192 30676 10198 30728
rect 10410 30676 10416 30728
rect 10468 30716 10474 30728
rect 10594 30716 10600 30728
rect 10468 30688 10600 30716
rect 10468 30676 10474 30688
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 10796 30725 10824 30756
rect 13449 30753 13461 30787
rect 13495 30753 13507 30787
rect 13449 30747 13507 30753
rect 13633 30787 13691 30793
rect 13633 30753 13645 30787
rect 13679 30784 13691 30787
rect 13679 30756 14964 30784
rect 13679 30753 13691 30756
rect 13633 30747 13691 30753
rect 14936 30728 14964 30756
rect 15746 30744 15752 30796
rect 15804 30744 15810 30796
rect 10781 30719 10839 30725
rect 10781 30685 10793 30719
rect 10827 30685 10839 30719
rect 10781 30679 10839 30685
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 14090 30716 14096 30728
rect 13771 30688 14096 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 14090 30676 14096 30688
rect 14148 30716 14154 30728
rect 14550 30716 14556 30728
rect 14148 30688 14556 30716
rect 14148 30676 14154 30688
rect 14550 30676 14556 30688
rect 14608 30716 14614 30728
rect 14645 30719 14703 30725
rect 14645 30716 14657 30719
rect 14608 30688 14657 30716
rect 14608 30676 14614 30688
rect 14645 30685 14657 30688
rect 14691 30685 14703 30719
rect 14645 30679 14703 30685
rect 14918 30676 14924 30728
rect 14976 30716 14982 30728
rect 15013 30719 15071 30725
rect 15013 30716 15025 30719
rect 14976 30688 15025 30716
rect 14976 30676 14982 30688
rect 15013 30685 15025 30688
rect 15059 30685 15071 30719
rect 15013 30679 15071 30685
rect 15562 30676 15568 30728
rect 15620 30676 15626 30728
rect 16022 30676 16028 30728
rect 16080 30676 16086 30728
rect 16224 30725 16252 30824
rect 23109 30821 23121 30855
rect 23155 30852 23167 30855
rect 23382 30852 23388 30864
rect 23155 30824 23388 30852
rect 23155 30821 23167 30824
rect 23109 30815 23167 30821
rect 23382 30812 23388 30824
rect 23440 30852 23446 30864
rect 27525 30855 27583 30861
rect 27525 30852 27537 30855
rect 23440 30824 27537 30852
rect 23440 30812 23446 30824
rect 27525 30821 27537 30824
rect 27571 30821 27583 30855
rect 27525 30815 27583 30821
rect 20625 30787 20683 30793
rect 20625 30753 20637 30787
rect 20671 30784 20683 30787
rect 23750 30784 23756 30796
rect 20671 30756 23756 30784
rect 20671 30753 20683 30756
rect 20625 30747 20683 30753
rect 22940 30728 22968 30756
rect 23750 30744 23756 30756
rect 23808 30784 23814 30796
rect 24670 30784 24676 30796
rect 23808 30756 24676 30784
rect 23808 30744 23814 30756
rect 24670 30744 24676 30756
rect 24728 30744 24734 30796
rect 25222 30744 25228 30796
rect 25280 30784 25286 30796
rect 29086 30784 29092 30796
rect 25280 30756 26280 30784
rect 25280 30744 25286 30756
rect 16209 30719 16267 30725
rect 16209 30685 16221 30719
rect 16255 30685 16267 30719
rect 16209 30679 16267 30685
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30716 20867 30719
rect 21450 30716 21456 30728
rect 20855 30688 21456 30716
rect 20855 30685 20867 30688
rect 20809 30679 20867 30685
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 22922 30676 22928 30728
rect 22980 30676 22986 30728
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 25038 30676 25044 30728
rect 25096 30676 25102 30728
rect 25590 30676 25596 30728
rect 25648 30676 25654 30728
rect 25774 30676 25780 30728
rect 25832 30676 25838 30728
rect 26252 30725 26280 30756
rect 28460 30756 29092 30784
rect 28460 30728 28488 30756
rect 29086 30744 29092 30756
rect 29144 30744 29150 30796
rect 26237 30719 26295 30725
rect 26237 30685 26249 30719
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 27706 30676 27712 30728
rect 27764 30676 27770 30728
rect 28077 30719 28135 30725
rect 28077 30685 28089 30719
rect 28123 30685 28135 30719
rect 28077 30679 28135 30685
rect 10612 30648 10640 30676
rect 17586 30648 17592 30660
rect 10612 30620 17592 30648
rect 17586 30608 17592 30620
rect 17644 30648 17650 30660
rect 20990 30648 20996 30660
rect 17644 30620 20996 30648
rect 17644 30608 17650 30620
rect 20990 30608 20996 30620
rect 21048 30608 21054 30660
rect 26142 30608 26148 30660
rect 26200 30608 26206 30660
rect 27614 30608 27620 30660
rect 27672 30648 27678 30660
rect 28092 30648 28120 30679
rect 28442 30676 28448 30728
rect 28500 30676 28506 30728
rect 28902 30676 28908 30728
rect 28960 30676 28966 30728
rect 28718 30648 28724 30660
rect 27672 30620 28724 30648
rect 27672 30608 27678 30620
rect 28718 30608 28724 30620
rect 28776 30608 28782 30660
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 28994 30336 29000 30388
rect 29052 30336 29058 30388
rect 29086 30336 29092 30388
rect 29144 30376 29150 30388
rect 29733 30379 29791 30385
rect 29733 30376 29745 30379
rect 29144 30348 29745 30376
rect 29144 30336 29150 30348
rect 29733 30345 29745 30348
rect 29779 30345 29791 30379
rect 29733 30339 29791 30345
rect 16022 30268 16028 30320
rect 16080 30308 16086 30320
rect 16080 30280 18814 30308
rect 16080 30268 16086 30280
rect 25038 30268 25044 30320
rect 25096 30308 25102 30320
rect 25682 30308 25688 30320
rect 25096 30280 25688 30308
rect 25096 30268 25102 30280
rect 25682 30268 25688 30280
rect 25740 30308 25746 30320
rect 27706 30308 27712 30320
rect 25740 30280 26096 30308
rect 25740 30268 25746 30280
rect 14274 30200 14280 30252
rect 14332 30200 14338 30252
rect 14918 30200 14924 30252
rect 14976 30200 14982 30252
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20162 30240 20168 30252
rect 19751 30212 20168 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20806 30240 20812 30252
rect 20303 30212 20812 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 20898 30200 20904 30252
rect 20956 30240 20962 30252
rect 20993 30243 21051 30249
rect 20993 30240 21005 30243
rect 20956 30212 21005 30240
rect 20956 30200 20962 30212
rect 20993 30209 21005 30212
rect 21039 30209 21051 30243
rect 20993 30203 21051 30209
rect 24670 30200 24676 30252
rect 24728 30200 24734 30252
rect 25130 30200 25136 30252
rect 25188 30200 25194 30252
rect 25222 30200 25228 30252
rect 25280 30240 25286 30252
rect 25317 30243 25375 30249
rect 25317 30240 25329 30243
rect 25280 30212 25329 30240
rect 25280 30200 25286 30212
rect 25317 30209 25329 30212
rect 25363 30209 25375 30243
rect 25317 30203 25375 30209
rect 25774 30200 25780 30252
rect 25832 30200 25838 30252
rect 26068 30249 26096 30280
rect 27356 30280 27712 30308
rect 27356 30249 27384 30280
rect 27706 30268 27712 30280
rect 27764 30268 27770 30320
rect 28074 30268 28080 30320
rect 28132 30268 28138 30320
rect 28537 30311 28595 30317
rect 28537 30277 28549 30311
rect 28583 30308 28595 30311
rect 29012 30308 29040 30336
rect 28583 30280 29040 30308
rect 28583 30277 28595 30280
rect 28537 30271 28595 30277
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 26053 30243 26111 30249
rect 26053 30209 26065 30243
rect 26099 30209 26111 30243
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 26053 30203 26111 30209
rect 26206 30212 27353 30240
rect 25590 30132 25596 30184
rect 25648 30172 25654 30184
rect 25884 30172 25912 30203
rect 26206 30184 26234 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 27522 30200 27528 30252
rect 27580 30240 27586 30252
rect 27617 30243 27675 30249
rect 27617 30240 27629 30243
rect 27580 30212 27629 30240
rect 27580 30200 27586 30212
rect 27617 30209 27629 30212
rect 27663 30240 27675 30243
rect 28442 30240 28448 30252
rect 27663 30212 28448 30240
rect 27663 30209 27675 30212
rect 27617 30203 27675 30209
rect 28442 30200 28448 30212
rect 28500 30200 28506 30252
rect 25648 30144 25912 30172
rect 25648 30132 25654 30144
rect 26142 30132 26148 30184
rect 26200 30132 26234 30184
rect 27433 30175 27491 30181
rect 27433 30141 27445 30175
rect 27479 30172 27491 30175
rect 28552 30172 28580 30271
rect 28718 30200 28724 30252
rect 28776 30200 28782 30252
rect 28994 30200 29000 30252
rect 29052 30200 29058 30252
rect 29178 30200 29184 30252
rect 29236 30200 29242 30252
rect 29638 30200 29644 30252
rect 29696 30200 29702 30252
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 27479 30144 28580 30172
rect 27479 30141 27491 30144
rect 27433 30135 27491 30141
rect 25774 30064 25780 30116
rect 25832 30104 25838 30116
rect 26206 30104 26234 30132
rect 25832 30076 26234 30104
rect 25832 30064 25838 30076
rect 28074 30064 28080 30116
rect 28132 30104 28138 30116
rect 29840 30104 29868 30203
rect 28132 30076 29868 30104
rect 28132 30064 28138 30076
rect 12894 29996 12900 30048
rect 12952 30036 12958 30048
rect 13449 30039 13507 30045
rect 13449 30036 13461 30039
rect 12952 30008 13461 30036
rect 12952 29996 12958 30008
rect 13449 30005 13461 30008
rect 13495 30005 13507 30039
rect 13449 29999 13507 30005
rect 20622 29996 20628 30048
rect 20680 30036 20686 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 20680 30008 20913 30036
rect 20680 29996 20686 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 20901 29999 20959 30005
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 14826 29792 14832 29844
rect 14884 29792 14890 29844
rect 25038 29792 25044 29844
rect 25096 29792 25102 29844
rect 25130 29792 25136 29844
rect 25188 29832 25194 29844
rect 25188 29804 28580 29832
rect 25188 29792 25194 29804
rect 9030 29724 9036 29776
rect 9088 29764 9094 29776
rect 10413 29767 10471 29773
rect 10413 29764 10425 29767
rect 9088 29736 10425 29764
rect 9088 29724 9094 29736
rect 10413 29733 10425 29736
rect 10459 29733 10471 29767
rect 10413 29727 10471 29733
rect 19720 29736 22094 29764
rect 10686 29696 10692 29708
rect 9968 29668 10692 29696
rect 9968 29637 9996 29668
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29597 9735 29631
rect 9677 29591 9735 29597
rect 9953 29631 10011 29637
rect 9953 29597 9965 29631
rect 9999 29597 10011 29631
rect 9953 29591 10011 29597
rect 9692 29560 9720 29591
rect 10410 29588 10416 29640
rect 10468 29588 10474 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 12894 29628 12900 29640
rect 10551 29600 12900 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10134 29560 10140 29572
rect 9692 29532 10140 29560
rect 10134 29520 10140 29532
rect 10192 29560 10198 29572
rect 10520 29560 10548 29591
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13173 29631 13231 29637
rect 13173 29597 13185 29631
rect 13219 29628 13231 29631
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 13219 29600 14933 29628
rect 13219 29597 13231 29600
rect 13173 29591 13231 29597
rect 14921 29597 14933 29600
rect 14967 29628 14979 29631
rect 15010 29628 15016 29640
rect 14967 29600 15016 29628
rect 14967 29597 14979 29600
rect 14921 29591 14979 29597
rect 10192 29532 10548 29560
rect 10192 29520 10198 29532
rect 10686 29520 10692 29572
rect 10744 29520 10750 29572
rect 13004 29560 13032 29591
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 19610 29588 19616 29640
rect 19668 29628 19674 29640
rect 19720 29628 19748 29736
rect 20441 29699 20499 29705
rect 20441 29665 20453 29699
rect 20487 29696 20499 29699
rect 20530 29696 20536 29708
rect 20487 29668 20536 29696
rect 20487 29665 20499 29668
rect 20441 29659 20499 29665
rect 20530 29656 20536 29668
rect 20588 29656 20594 29708
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21545 29699 21603 29705
rect 21545 29696 21557 29699
rect 20864 29668 21557 29696
rect 20864 29656 20870 29668
rect 21545 29665 21557 29668
rect 21591 29665 21603 29699
rect 22066 29696 22094 29736
rect 23198 29724 23204 29776
rect 23256 29764 23262 29776
rect 27341 29767 27399 29773
rect 27341 29764 27353 29767
rect 23256 29736 27353 29764
rect 23256 29724 23262 29736
rect 27341 29733 27353 29736
rect 27387 29733 27399 29767
rect 27341 29727 27399 29733
rect 27706 29724 27712 29776
rect 27764 29724 27770 29776
rect 27154 29696 27160 29708
rect 22066 29668 27160 29696
rect 21545 29659 21603 29665
rect 27154 29656 27160 29668
rect 27212 29656 27218 29708
rect 19668 29600 19748 29628
rect 20165 29631 20223 29637
rect 19668 29588 19674 29600
rect 20165 29597 20177 29631
rect 20211 29628 20223 29631
rect 20346 29628 20352 29640
rect 20211 29600 20352 29628
rect 20211 29597 20223 29600
rect 20165 29591 20223 29597
rect 20346 29588 20352 29600
rect 20404 29588 20410 29640
rect 20714 29588 20720 29640
rect 20772 29628 20778 29640
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20772 29600 21005 29628
rect 20772 29588 20778 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 14182 29560 14188 29572
rect 13004 29532 14188 29560
rect 14182 29520 14188 29532
rect 14240 29520 14246 29572
rect 15102 29520 15108 29572
rect 15160 29520 15166 29572
rect 20898 29520 20904 29572
rect 20956 29560 20962 29572
rect 21376 29560 21404 29591
rect 24762 29588 24768 29640
rect 24820 29588 24826 29640
rect 24854 29588 24860 29640
rect 24912 29588 24918 29640
rect 27522 29588 27528 29640
rect 27580 29588 27586 29640
rect 27614 29588 27620 29640
rect 27672 29588 27678 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 21634 29560 21640 29572
rect 20956 29532 21640 29560
rect 20956 29520 20962 29532
rect 21634 29520 21640 29532
rect 21692 29520 21698 29572
rect 27816 29560 27844 29591
rect 28350 29588 28356 29640
rect 28408 29588 28414 29640
rect 28552 29637 28580 29804
rect 28902 29764 28908 29776
rect 28736 29736 28908 29764
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28736 29560 28764 29736
rect 28902 29724 28908 29736
rect 28960 29764 28966 29776
rect 30009 29767 30067 29773
rect 30009 29764 30021 29767
rect 28960 29736 30021 29764
rect 28960 29724 28966 29736
rect 30009 29733 30021 29736
rect 30055 29733 30067 29767
rect 30009 29727 30067 29733
rect 28813 29699 28871 29705
rect 28813 29665 28825 29699
rect 28859 29696 28871 29699
rect 28994 29696 29000 29708
rect 28859 29668 29000 29696
rect 28859 29665 28871 29668
rect 28813 29659 28871 29665
rect 28994 29656 29000 29668
rect 29052 29696 29058 29708
rect 29052 29668 29960 29696
rect 29052 29656 29058 29668
rect 28902 29588 28908 29640
rect 28960 29588 28966 29640
rect 29178 29588 29184 29640
rect 29236 29628 29242 29640
rect 29932 29637 29960 29668
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29236 29600 29745 29628
rect 29236 29588 29242 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 27816 29532 28764 29560
rect 9306 29452 9312 29504
rect 9364 29492 9370 29504
rect 9493 29495 9551 29501
rect 9493 29492 9505 29495
rect 9364 29464 9505 29492
rect 9364 29452 9370 29464
rect 9493 29461 9505 29464
rect 9539 29461 9551 29495
rect 9493 29455 9551 29461
rect 9861 29495 9919 29501
rect 9861 29461 9873 29495
rect 9907 29492 9919 29495
rect 9950 29492 9956 29504
rect 9907 29464 9956 29492
rect 9907 29461 9919 29464
rect 9861 29455 9919 29461
rect 9950 29452 9956 29464
rect 10008 29492 10014 29504
rect 10410 29492 10416 29504
rect 10008 29464 10416 29492
rect 10008 29452 10014 29464
rect 10410 29452 10416 29464
rect 10468 29492 10474 29504
rect 12710 29492 12716 29504
rect 10468 29464 12716 29492
rect 10468 29452 10474 29464
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 12802 29452 12808 29504
rect 12860 29452 12866 29504
rect 19518 29452 19524 29504
rect 19576 29452 19582 29504
rect 21361 29495 21419 29501
rect 21361 29461 21373 29495
rect 21407 29492 21419 29495
rect 21450 29492 21456 29504
rect 21407 29464 21456 29492
rect 21407 29461 21419 29464
rect 21361 29455 21419 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 14550 29248 14556 29300
rect 14608 29248 14614 29300
rect 14918 29248 14924 29300
rect 14976 29288 14982 29300
rect 14976 29260 17724 29288
rect 14976 29248 14982 29260
rect 12912 29220 12940 29248
rect 12544 29192 12940 29220
rect 9030 29112 9036 29164
rect 9088 29112 9094 29164
rect 9306 29112 9312 29164
rect 9364 29112 9370 29164
rect 9490 29112 9496 29164
rect 9548 29112 9554 29164
rect 11882 29112 11888 29164
rect 11940 29112 11946 29164
rect 12544 29161 12572 29192
rect 15102 29180 15108 29232
rect 15160 29220 15166 29232
rect 17696 29229 17724 29260
rect 20162 29248 20168 29300
rect 20220 29248 20226 29300
rect 21358 29248 21364 29300
rect 21416 29288 21422 29300
rect 22097 29291 22155 29297
rect 22097 29288 22109 29291
rect 21416 29260 22109 29288
rect 21416 29248 21422 29260
rect 22097 29257 22109 29260
rect 22143 29257 22155 29291
rect 22097 29251 22155 29257
rect 27154 29248 27160 29300
rect 27212 29288 27218 29300
rect 27522 29288 27528 29300
rect 27212 29260 27528 29288
rect 27212 29248 27218 29260
rect 27522 29248 27528 29260
rect 27580 29248 27586 29300
rect 27614 29248 27620 29300
rect 27672 29288 27678 29300
rect 27893 29291 27951 29297
rect 27893 29288 27905 29291
rect 27672 29260 27905 29288
rect 27672 29248 27678 29260
rect 27893 29257 27905 29260
rect 27939 29257 27951 29291
rect 27893 29251 27951 29257
rect 28350 29248 28356 29300
rect 28408 29288 28414 29300
rect 28921 29291 28979 29297
rect 28921 29288 28933 29291
rect 28408 29260 28933 29288
rect 28408 29248 28414 29260
rect 28921 29257 28933 29260
rect 28967 29257 28979 29291
rect 28921 29251 28979 29257
rect 29089 29291 29147 29297
rect 29089 29257 29101 29291
rect 29135 29288 29147 29291
rect 29178 29288 29184 29300
rect 29135 29260 29184 29288
rect 29135 29257 29147 29260
rect 29089 29251 29147 29257
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 15381 29223 15439 29229
rect 15381 29220 15393 29223
rect 15160 29192 15393 29220
rect 15160 29180 15166 29192
rect 15381 29189 15393 29192
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 17681 29223 17739 29229
rect 17681 29189 17693 29223
rect 17727 29189 17739 29223
rect 20530 29220 20536 29232
rect 17681 29183 17739 29189
rect 20364 29192 20536 29220
rect 12529 29155 12587 29161
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29152 12679 29155
rect 12710 29152 12716 29164
rect 12667 29124 12716 29152
rect 12667 29121 12679 29124
rect 12621 29115 12679 29121
rect 12710 29112 12716 29124
rect 12768 29112 12774 29164
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 12897 29155 12955 29161
rect 12897 29152 12909 29155
rect 12860 29124 12909 29152
rect 12860 29112 12866 29124
rect 12897 29121 12909 29124
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13354 29152 13360 29164
rect 13219 29124 13360 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 13354 29112 13360 29124
rect 13412 29112 13418 29164
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29152 14795 29155
rect 15120 29152 15148 29180
rect 14783 29124 15148 29152
rect 14783 29121 14795 29124
rect 14737 29115 14795 29121
rect 15562 29112 15568 29164
rect 15620 29112 15626 29164
rect 15749 29155 15807 29161
rect 15749 29121 15761 29155
rect 15795 29152 15807 29155
rect 16390 29152 16396 29164
rect 15795 29124 16396 29152
rect 15795 29121 15807 29124
rect 15749 29115 15807 29121
rect 16390 29112 16396 29124
rect 16448 29112 16454 29164
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29152 19211 29155
rect 19334 29152 19340 29164
rect 19199 29124 19340 29152
rect 19199 29121 19211 29124
rect 19153 29115 19211 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 19518 29112 19524 29164
rect 19576 29112 19582 29164
rect 20364 29161 20392 29192
rect 20530 29180 20536 29192
rect 20588 29220 20594 29232
rect 20588 29192 21404 29220
rect 20588 29180 20594 29192
rect 20349 29155 20407 29161
rect 20349 29121 20361 29155
rect 20395 29121 20407 29155
rect 20349 29115 20407 29121
rect 20438 29112 20444 29164
rect 20496 29112 20502 29164
rect 20622 29112 20628 29164
rect 20680 29112 20686 29164
rect 20714 29112 20720 29164
rect 20772 29112 20778 29164
rect 21376 29161 21404 29192
rect 21634 29180 21640 29232
rect 21692 29220 21698 29232
rect 21692 29192 22600 29220
rect 21692 29180 21698 29192
rect 21177 29155 21235 29161
rect 21177 29121 21189 29155
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29152 22339 29155
rect 22370 29152 22376 29164
rect 22327 29124 22376 29152
rect 22327 29121 22339 29124
rect 22281 29115 22339 29121
rect 12434 29044 12440 29096
rect 12492 29044 12498 29096
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29084 14979 29087
rect 15010 29084 15016 29096
rect 14967 29056 15016 29084
rect 14967 29053 14979 29056
rect 14921 29047 14979 29053
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 20456 29016 20484 29112
rect 21192 29016 21220 29115
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22572 29161 22600 29192
rect 25222 29180 25228 29232
rect 25280 29180 25286 29232
rect 27249 29223 27307 29229
rect 27249 29189 27261 29223
rect 27295 29220 27307 29223
rect 28721 29223 28779 29229
rect 28721 29220 28733 29223
rect 27295 29192 28120 29220
rect 27295 29189 27307 29192
rect 27249 29183 27307 29189
rect 28092 29164 28120 29192
rect 28184 29192 28733 29220
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 22738 29112 22744 29164
rect 22796 29112 22802 29164
rect 23474 29112 23480 29164
rect 23532 29152 23538 29164
rect 24486 29152 24492 29164
rect 23532 29124 24492 29152
rect 23532 29112 23538 29124
rect 24486 29112 24492 29124
rect 24544 29152 24550 29164
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 24544 29124 25329 29152
rect 24544 29112 24550 29124
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29152 25651 29155
rect 26050 29152 26056 29164
rect 25639 29124 26056 29152
rect 25639 29121 25651 29124
rect 25593 29115 25651 29121
rect 26050 29112 26056 29124
rect 26108 29112 26114 29164
rect 27154 29112 27160 29164
rect 27212 29112 27218 29164
rect 27338 29112 27344 29164
rect 27396 29112 27402 29164
rect 28074 29112 28080 29164
rect 28132 29112 28138 29164
rect 26786 29044 26792 29096
rect 26844 29084 26850 29096
rect 28184 29084 28212 29192
rect 28721 29189 28733 29192
rect 28767 29189 28779 29223
rect 28721 29183 28779 29189
rect 26844 29056 28212 29084
rect 28261 29087 28319 29093
rect 26844 29044 26850 29056
rect 28261 29053 28273 29087
rect 28307 29084 28319 29087
rect 29638 29084 29644 29096
rect 28307 29056 29644 29084
rect 28307 29053 28319 29056
rect 28261 29047 28319 29053
rect 20456 28988 21220 29016
rect 21266 28976 21272 29028
rect 21324 28976 21330 29028
rect 22373 29019 22431 29025
rect 22373 29016 22385 29019
rect 22066 28988 22385 29016
rect 8938 28908 8944 28960
rect 8996 28948 9002 28960
rect 9401 28951 9459 28957
rect 9401 28948 9413 28951
rect 8996 28920 9413 28948
rect 8996 28908 9002 28920
rect 9401 28917 9413 28920
rect 9447 28917 9459 28951
rect 9401 28911 9459 28917
rect 20714 28908 20720 28960
rect 20772 28948 20778 28960
rect 22066 28948 22094 28988
rect 22373 28985 22385 28988
rect 22419 28985 22431 29019
rect 22373 28979 22431 28985
rect 22465 29019 22523 29025
rect 22465 28985 22477 29019
rect 22511 29016 22523 29019
rect 23198 29016 23204 29028
rect 22511 28988 23204 29016
rect 22511 28985 22523 28988
rect 22465 28979 22523 28985
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 28276 29016 28304 29047
rect 29638 29044 29644 29056
rect 29696 29044 29702 29096
rect 27488 28988 28304 29016
rect 27488 28976 27494 28988
rect 20772 28920 22094 28948
rect 20772 28908 20778 28920
rect 28902 28908 28908 28960
rect 28960 28908 28966 28960
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 21174 28704 21180 28756
rect 21232 28704 21238 28756
rect 28813 28747 28871 28753
rect 28813 28713 28825 28747
rect 28859 28744 28871 28747
rect 28902 28744 28908 28756
rect 28859 28716 28908 28744
rect 28859 28713 28871 28716
rect 28813 28707 28871 28713
rect 28902 28704 28908 28716
rect 28960 28704 28966 28756
rect 12434 28636 12440 28688
rect 12492 28676 12498 28688
rect 12802 28676 12808 28688
rect 12492 28648 12808 28676
rect 12492 28636 12498 28648
rect 12802 28636 12808 28648
rect 12860 28636 12866 28688
rect 15197 28679 15255 28685
rect 15197 28676 15209 28679
rect 13464 28648 15209 28676
rect 9490 28608 9496 28620
rect 9324 28580 9496 28608
rect 9324 28549 9352 28580
rect 9490 28568 9496 28580
rect 9548 28608 9554 28620
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 9548 28580 10977 28608
rect 9548 28568 9554 28580
rect 10965 28577 10977 28580
rect 11011 28577 11023 28611
rect 10965 28571 11023 28577
rect 11609 28611 11667 28617
rect 11609 28577 11621 28611
rect 11655 28608 11667 28611
rect 11882 28608 11888 28620
rect 11655 28580 11888 28608
rect 11655 28577 11667 28580
rect 11609 28571 11667 28577
rect 11882 28568 11888 28580
rect 11940 28608 11946 28620
rect 12526 28608 12532 28620
rect 11940 28580 12532 28608
rect 11940 28568 11946 28580
rect 12526 28568 12532 28580
rect 12584 28608 12590 28620
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12584 28580 13185 28608
rect 12584 28568 12590 28580
rect 13173 28577 13185 28580
rect 13219 28577 13231 28611
rect 13173 28571 13231 28577
rect 13354 28568 13360 28620
rect 13412 28608 13418 28620
rect 13464 28608 13492 28648
rect 15197 28645 15209 28648
rect 15243 28645 15255 28679
rect 27338 28676 27344 28688
rect 15197 28639 15255 28645
rect 24044 28648 27344 28676
rect 13412 28580 13492 28608
rect 13412 28568 13418 28580
rect 15010 28568 15016 28620
rect 15068 28608 15074 28620
rect 15068 28580 19932 28608
rect 15068 28568 15074 28580
rect 19904 28552 19932 28580
rect 20806 28568 20812 28620
rect 20864 28608 20870 28620
rect 20864 28580 21036 28608
rect 20864 28568 20870 28580
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 9309 28503 9367 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 9030 28432 9036 28484
rect 9088 28472 9094 28484
rect 9600 28472 9628 28503
rect 10686 28500 10692 28552
rect 10744 28540 10750 28552
rect 11241 28543 11299 28549
rect 11241 28540 11253 28543
rect 10744 28512 11253 28540
rect 10744 28500 10750 28512
rect 11241 28509 11253 28512
rect 11287 28509 11299 28543
rect 11241 28503 11299 28509
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28540 12403 28543
rect 12434 28540 12440 28552
rect 12391 28512 12440 28540
rect 12391 28509 12403 28512
rect 12345 28503 12403 28509
rect 9088 28444 9628 28472
rect 12084 28472 12112 28503
rect 12434 28500 12440 28512
rect 12492 28500 12498 28552
rect 13081 28543 13139 28549
rect 13081 28509 13093 28543
rect 13127 28509 13139 28543
rect 13081 28503 13139 28509
rect 12618 28472 12624 28484
rect 12084 28444 12624 28472
rect 9088 28432 9094 28444
rect 12618 28432 12624 28444
rect 12676 28432 12682 28484
rect 13096 28472 13124 28503
rect 13262 28500 13268 28552
rect 13320 28500 13326 28552
rect 14550 28500 14556 28552
rect 14608 28500 14614 28552
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28540 14979 28543
rect 15102 28540 15108 28552
rect 14967 28512 15108 28540
rect 14967 28509 14979 28512
rect 14921 28503 14979 28509
rect 15102 28500 15108 28512
rect 15160 28500 15166 28552
rect 15378 28500 15384 28552
rect 15436 28500 15442 28552
rect 15746 28500 15752 28552
rect 15804 28540 15810 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 15804 28512 16313 28540
rect 15804 28500 15810 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 16390 28500 16396 28552
rect 16448 28540 16454 28552
rect 16669 28543 16727 28549
rect 16669 28540 16681 28543
rect 16448 28512 16681 28540
rect 16448 28500 16454 28512
rect 16669 28509 16681 28512
rect 16715 28540 16727 28543
rect 19610 28540 19616 28552
rect 16715 28512 19616 28540
rect 16715 28509 16727 28512
rect 16669 28503 16727 28509
rect 19610 28500 19616 28512
rect 19668 28500 19674 28552
rect 19886 28500 19892 28552
rect 19944 28500 19950 28552
rect 19978 28500 19984 28552
rect 20036 28500 20042 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 20088 28512 20637 28540
rect 15930 28472 15936 28484
rect 12820 28444 15936 28472
rect 9122 28364 9128 28416
rect 9180 28364 9186 28416
rect 9306 28364 9312 28416
rect 9364 28404 9370 28416
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 9364 28376 9505 28404
rect 9364 28364 9370 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 9493 28367 9551 28373
rect 12342 28364 12348 28416
rect 12400 28404 12406 28416
rect 12820 28404 12848 28444
rect 15930 28432 15936 28444
rect 15988 28432 15994 28484
rect 18414 28432 18420 28484
rect 18472 28472 18478 28484
rect 20088 28472 20116 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 20625 28503 20683 28509
rect 20714 28500 20720 28552
rect 20772 28500 20778 28552
rect 20898 28500 20904 28552
rect 20956 28500 20962 28552
rect 21008 28549 21036 28580
rect 20993 28543 21051 28549
rect 20993 28509 21005 28543
rect 21039 28540 21051 28543
rect 23293 28543 23351 28549
rect 21039 28512 22094 28540
rect 21039 28509 21051 28512
rect 20993 28503 21051 28509
rect 18472 28444 20116 28472
rect 18472 28432 18478 28444
rect 12400 28376 12848 28404
rect 12400 28364 12406 28376
rect 12894 28364 12900 28416
rect 12952 28364 12958 28416
rect 20088 28404 20116 28444
rect 20165 28475 20223 28481
rect 20165 28441 20177 28475
rect 20211 28472 20223 28475
rect 20732 28472 20760 28500
rect 20211 28444 20760 28472
rect 22066 28472 22094 28512
rect 23293 28509 23305 28543
rect 23339 28509 23351 28543
rect 23293 28503 23351 28509
rect 23308 28472 23336 28503
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 23937 28543 23995 28549
rect 23937 28540 23949 28543
rect 23440 28512 23949 28540
rect 23440 28500 23446 28512
rect 23937 28509 23949 28512
rect 23983 28540 23995 28543
rect 24044 28540 24072 28648
rect 27338 28636 27344 28648
rect 27396 28636 27402 28688
rect 26237 28611 26295 28617
rect 26237 28577 26249 28611
rect 26283 28608 26295 28611
rect 26694 28608 26700 28620
rect 26283 28580 26700 28608
rect 26283 28577 26295 28580
rect 26237 28571 26295 28577
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 28350 28608 28356 28620
rect 28014 28580 28356 28608
rect 28350 28568 28356 28580
rect 28408 28568 28414 28620
rect 27890 28540 27896 28552
rect 23983 28512 24072 28540
rect 27738 28512 27896 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28718 28500 28724 28552
rect 28776 28500 28782 28552
rect 23658 28472 23664 28484
rect 22066 28444 22494 28472
rect 23308 28444 23664 28472
rect 20211 28441 20223 28444
rect 20165 28435 20223 28441
rect 23658 28432 23664 28444
rect 23716 28472 23722 28484
rect 24670 28472 24676 28484
rect 23716 28444 24676 28472
rect 23716 28432 23722 28444
rect 24670 28432 24676 28444
rect 24728 28432 24734 28484
rect 22738 28404 22744 28416
rect 20088 28376 22744 28404
rect 22738 28364 22744 28376
rect 22796 28364 22802 28416
rect 27246 28364 27252 28416
rect 27304 28364 27310 28416
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 8113 28203 8171 28209
rect 8113 28169 8125 28203
rect 8159 28200 8171 28203
rect 8938 28200 8944 28212
rect 8159 28172 8944 28200
rect 8159 28169 8171 28172
rect 8113 28163 8171 28169
rect 8938 28160 8944 28172
rect 8996 28160 9002 28212
rect 13354 28160 13360 28212
rect 13412 28160 13418 28212
rect 15378 28160 15384 28212
rect 15436 28160 15442 28212
rect 19610 28200 19616 28212
rect 19260 28172 19616 28200
rect 8846 28132 8852 28144
rect 7944 28104 8852 28132
rect 7944 28073 7972 28104
rect 8846 28092 8852 28104
rect 8904 28092 8910 28144
rect 9140 28104 9904 28132
rect 9140 28076 9168 28104
rect 7929 28067 7987 28073
rect 7929 28033 7941 28067
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28064 8263 28067
rect 9033 28067 9091 28073
rect 9033 28064 9045 28067
rect 8251 28036 9045 28064
rect 8251 28033 8263 28036
rect 8205 28027 8263 28033
rect 9033 28033 9045 28036
rect 9079 28064 9091 28067
rect 9122 28064 9128 28076
rect 9079 28036 9128 28064
rect 9079 28033 9091 28036
rect 9033 28027 9091 28033
rect 9122 28024 9128 28036
rect 9180 28024 9186 28076
rect 9876 28073 9904 28104
rect 12618 28092 12624 28144
rect 12676 28132 12682 28144
rect 13372 28132 13400 28160
rect 15010 28132 15016 28144
rect 12676 28104 13400 28132
rect 14016 28104 15016 28132
rect 12676 28092 12682 28104
rect 9677 28067 9735 28073
rect 9677 28033 9689 28067
rect 9723 28033 9735 28067
rect 9677 28027 9735 28033
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 8754 27956 8760 28008
rect 8812 27956 8818 28008
rect 8846 27956 8852 28008
rect 8904 27956 8910 28008
rect 8938 27956 8944 28008
rect 8996 27996 9002 28008
rect 9692 27996 9720 28027
rect 10686 28024 10692 28076
rect 10744 28064 10750 28076
rect 11885 28067 11943 28073
rect 11885 28064 11897 28067
rect 10744 28036 11897 28064
rect 10744 28024 10750 28036
rect 11885 28033 11897 28036
rect 11931 28064 11943 28067
rect 12342 28064 12348 28076
rect 11931 28036 12348 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12342 28024 12348 28036
rect 12400 28024 12406 28076
rect 12526 28024 12532 28076
rect 12584 28024 12590 28076
rect 12912 28073 12940 28104
rect 14016 28076 14044 28104
rect 15010 28092 15016 28104
rect 15068 28092 15074 28144
rect 15562 28092 15568 28144
rect 15620 28132 15626 28144
rect 15933 28135 15991 28141
rect 15933 28132 15945 28135
rect 15620 28104 15945 28132
rect 15620 28092 15626 28104
rect 15933 28101 15945 28104
rect 15979 28132 15991 28135
rect 16022 28132 16028 28144
rect 15979 28104 16028 28132
rect 15979 28101 15991 28104
rect 15933 28095 15991 28101
rect 16022 28092 16028 28104
rect 16080 28092 16086 28144
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13262 28024 13268 28076
rect 13320 28064 13326 28076
rect 13357 28067 13415 28073
rect 13357 28064 13369 28067
rect 13320 28036 13369 28064
rect 13320 28024 13326 28036
rect 13357 28033 13369 28036
rect 13403 28064 13415 28067
rect 13817 28067 13875 28073
rect 13817 28064 13829 28067
rect 13403 28036 13829 28064
rect 13403 28033 13415 28036
rect 13357 28027 13415 28033
rect 13817 28033 13829 28036
rect 13863 28033 13875 28067
rect 13817 28027 13875 28033
rect 13998 28024 14004 28076
rect 14056 28024 14062 28076
rect 14182 28024 14188 28076
rect 14240 28024 14246 28076
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28064 15439 28067
rect 15746 28064 15752 28076
rect 15427 28036 15752 28064
rect 15427 28033 15439 28036
rect 15381 28027 15439 28033
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 19260 28073 19288 28172
rect 19610 28160 19616 28172
rect 19668 28160 19674 28212
rect 19886 28160 19892 28212
rect 19944 28200 19950 28212
rect 22281 28203 22339 28209
rect 19944 28172 22094 28200
rect 19944 28160 19950 28172
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 20625 28135 20683 28141
rect 19392 28104 19472 28132
rect 19392 28092 19398 28104
rect 19444 28073 19472 28104
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 20898 28132 20904 28144
rect 20671 28104 20904 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 20898 28092 20904 28104
rect 20956 28092 20962 28144
rect 22066 28132 22094 28172
rect 22281 28169 22293 28203
rect 22327 28200 22339 28203
rect 22370 28200 22376 28212
rect 22327 28172 22376 28200
rect 22327 28169 22339 28172
rect 22281 28163 22339 28169
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 23198 28160 23204 28212
rect 23256 28160 23262 28212
rect 26602 28132 26608 28144
rect 22066 28104 26608 28132
rect 26602 28092 26608 28104
rect 26660 28092 26666 28144
rect 27338 28092 27344 28144
rect 27396 28132 27402 28144
rect 30193 28135 30251 28141
rect 30193 28132 30205 28135
rect 27396 28104 30205 28132
rect 27396 28092 27402 28104
rect 30193 28101 30205 28104
rect 30239 28132 30251 28135
rect 31110 28132 31116 28144
rect 30239 28104 31116 28132
rect 30239 28101 30251 28104
rect 30193 28095 30251 28101
rect 31110 28092 31116 28104
rect 31168 28092 31174 28144
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 19429 28067 19487 28073
rect 19429 28033 19441 28067
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28064 20591 28067
rect 23658 28064 23664 28076
rect 20579 28036 22094 28064
rect 20579 28033 20591 28036
rect 20533 28027 20591 28033
rect 8996 27968 9720 27996
rect 8996 27956 9002 27968
rect 12434 27956 12440 28008
rect 12492 27956 12498 28008
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 14608 27968 15301 27996
rect 14608 27956 14614 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 19337 27999 19395 28005
rect 19337 27965 19349 27999
rect 19383 27996 19395 27999
rect 19978 27996 19984 28008
rect 19383 27968 19984 27996
rect 19383 27965 19395 27968
rect 19337 27959 19395 27965
rect 19978 27956 19984 27968
rect 20036 27996 20042 28008
rect 20272 27996 20300 28027
rect 20036 27968 20300 27996
rect 20036 27956 20042 27968
rect 7745 27863 7803 27869
rect 7745 27829 7757 27863
rect 7791 27860 7803 27863
rect 9122 27860 9128 27872
rect 7791 27832 9128 27860
rect 7791 27829 7803 27832
rect 7745 27823 7803 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9217 27863 9275 27869
rect 9217 27829 9229 27863
rect 9263 27860 9275 27863
rect 9306 27860 9312 27872
rect 9263 27832 9312 27860
rect 9263 27829 9275 27832
rect 9217 27823 9275 27829
rect 9306 27820 9312 27832
rect 9364 27860 9370 27872
rect 9582 27860 9588 27872
rect 9364 27832 9588 27860
rect 9364 27820 9370 27832
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 9766 27820 9772 27872
rect 9824 27820 9830 27872
rect 22066 27860 22094 28036
rect 22664 28036 23664 28064
rect 22465 27931 22523 27937
rect 22465 27897 22477 27931
rect 22511 27928 22523 27931
rect 22664 27928 22692 28036
rect 23658 28024 23664 28036
rect 23716 28024 23722 28076
rect 25038 28024 25044 28076
rect 25096 28024 25102 28076
rect 25406 28024 25412 28076
rect 25464 28064 25470 28076
rect 25685 28067 25743 28073
rect 25685 28064 25697 28067
rect 25464 28036 25697 28064
rect 25464 28024 25470 28036
rect 25685 28033 25697 28036
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27249 28067 27307 28073
rect 27249 28064 27261 28067
rect 27120 28036 27261 28064
rect 27120 28024 27126 28036
rect 27249 28033 27261 28036
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28064 27583 28067
rect 27706 28064 27712 28076
rect 27571 28036 27712 28064
rect 27571 28033 27583 28036
rect 27525 28027 27583 28033
rect 27706 28024 27712 28036
rect 27764 28024 27770 28076
rect 30006 28024 30012 28076
rect 30064 28024 30070 28076
rect 30285 28067 30343 28073
rect 30285 28033 30297 28067
rect 30331 28064 30343 28067
rect 32674 28064 32680 28076
rect 30331 28036 32680 28064
rect 30331 28033 30343 28036
rect 30285 28027 30343 28033
rect 32674 28024 32680 28036
rect 32732 28024 32738 28076
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27965 22799 27999
rect 22741 27959 22799 27965
rect 22511 27900 22692 27928
rect 22756 27928 22784 27959
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 26050 27956 26056 28008
rect 26108 27956 26114 28008
rect 26510 27956 26516 28008
rect 26568 27996 26574 28008
rect 27157 27999 27215 28005
rect 27157 27996 27169 27999
rect 26568 27968 27169 27996
rect 26568 27956 26574 27968
rect 27157 27965 27169 27968
rect 27203 27965 27215 27999
rect 27157 27959 27215 27965
rect 23382 27928 23388 27940
rect 22756 27900 23388 27928
rect 22511 27897 22523 27900
rect 22465 27891 22523 27897
rect 23382 27888 23388 27900
rect 23440 27888 23446 27940
rect 24857 27931 24915 27937
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25866 27928 25872 27940
rect 24903 27900 25872 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25866 27888 25872 27900
rect 25924 27888 25930 27940
rect 24670 27860 24676 27872
rect 22066 27832 24676 27860
rect 24670 27820 24676 27832
rect 24728 27820 24734 27872
rect 29822 27820 29828 27872
rect 29880 27820 29886 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 16022 27548 16028 27600
rect 16080 27588 16086 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 16080 27560 16865 27588
rect 16080 27548 16086 27560
rect 16853 27557 16865 27560
rect 16899 27557 16911 27591
rect 16853 27551 16911 27557
rect 24854 27548 24860 27600
rect 24912 27588 24918 27600
rect 25225 27591 25283 27597
rect 25225 27588 25237 27591
rect 24912 27560 25237 27588
rect 24912 27548 24918 27560
rect 25225 27557 25237 27560
rect 25271 27557 25283 27591
rect 26050 27588 26056 27600
rect 25225 27551 25283 27557
rect 25424 27560 26056 27588
rect 9030 27480 9036 27532
rect 9088 27520 9094 27532
rect 9217 27523 9275 27529
rect 9217 27520 9229 27523
rect 9088 27492 9229 27520
rect 9088 27480 9094 27492
rect 9217 27489 9229 27492
rect 9263 27489 9275 27523
rect 9217 27483 9275 27489
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 12805 27523 12863 27529
rect 12805 27520 12817 27523
rect 12584 27492 12817 27520
rect 12584 27480 12590 27492
rect 12805 27489 12817 27492
rect 12851 27489 12863 27523
rect 13998 27520 14004 27532
rect 12805 27483 12863 27489
rect 13188 27492 14004 27520
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 9180 27424 9321 27452
rect 9180 27412 9186 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 13188 27461 13216 27492
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 17218 27520 17224 27532
rect 15948 27492 17224 27520
rect 9677 27455 9735 27461
rect 9677 27452 9689 27455
rect 9640 27424 9689 27452
rect 9640 27412 9646 27424
rect 9677 27421 9689 27424
rect 9723 27421 9735 27455
rect 9677 27415 9735 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 14182 27452 14188 27464
rect 13403 27424 14188 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 15948 27461 15976 27492
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 20898 27520 20904 27532
rect 18156 27492 20904 27520
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 8202 27344 8208 27396
rect 8260 27384 8266 27396
rect 10137 27387 10195 27393
rect 10137 27384 10149 27387
rect 8260 27356 10149 27384
rect 8260 27344 8266 27356
rect 10137 27353 10149 27356
rect 10183 27384 10195 27387
rect 12342 27384 12348 27396
rect 10183 27356 12348 27384
rect 10183 27353 10195 27356
rect 10137 27347 10195 27353
rect 12342 27344 12348 27356
rect 12400 27344 12406 27396
rect 12710 27344 12716 27396
rect 12768 27384 12774 27396
rect 14369 27387 14427 27393
rect 14369 27384 14381 27387
rect 12768 27356 14381 27384
rect 12768 27344 12774 27356
rect 14369 27353 14381 27356
rect 14415 27353 14427 27387
rect 14369 27347 14427 27353
rect 14936 27316 14964 27415
rect 16022 27412 16028 27464
rect 16080 27412 16086 27464
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27452 16267 27455
rect 18156 27452 18184 27492
rect 20898 27480 20904 27492
rect 20956 27480 20962 27532
rect 20990 27480 20996 27532
rect 21048 27520 21054 27532
rect 21910 27520 21916 27532
rect 21048 27492 21916 27520
rect 21048 27480 21054 27492
rect 21910 27480 21916 27492
rect 21968 27520 21974 27532
rect 25038 27520 25044 27532
rect 21968 27492 25044 27520
rect 21968 27480 21974 27492
rect 25038 27480 25044 27492
rect 25096 27520 25102 27532
rect 25314 27520 25320 27532
rect 25096 27492 25320 27520
rect 25096 27480 25102 27492
rect 25314 27480 25320 27492
rect 25372 27480 25378 27532
rect 16255 27424 18184 27452
rect 16255 27421 16267 27424
rect 16209 27415 16267 27421
rect 18230 27412 18236 27464
rect 18288 27412 18294 27464
rect 22002 27412 22008 27464
rect 22060 27412 22066 27464
rect 25424 27461 25452 27560
rect 26050 27548 26056 27560
rect 26108 27548 26114 27600
rect 26620 27560 27476 27588
rect 26510 27520 26516 27532
rect 25976 27492 26516 27520
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 16393 27387 16451 27393
rect 16393 27353 16405 27387
rect 16439 27384 16451 27387
rect 17966 27387 18024 27393
rect 17966 27384 17978 27387
rect 16439 27356 17978 27384
rect 16439 27353 16451 27356
rect 16393 27347 16451 27353
rect 17966 27353 17978 27356
rect 18012 27353 18024 27387
rect 17966 27347 18024 27353
rect 20254 27344 20260 27396
rect 20312 27384 20318 27396
rect 22296 27384 22324 27415
rect 25682 27412 25688 27464
rect 25740 27412 25746 27464
rect 25976 27461 26004 27492
rect 26510 27480 26516 27492
rect 26568 27480 26574 27532
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27421 26019 27455
rect 25961 27415 26019 27421
rect 20312 27356 22324 27384
rect 20312 27344 20318 27356
rect 25590 27344 25596 27396
rect 25648 27384 25654 27396
rect 25976 27384 26004 27415
rect 26142 27412 26148 27464
rect 26200 27452 26206 27464
rect 26620 27461 26648 27560
rect 27448 27461 27476 27560
rect 27890 27548 27896 27600
rect 27948 27548 27954 27600
rect 28445 27523 28503 27529
rect 28445 27520 28457 27523
rect 27724 27492 28457 27520
rect 27724 27464 27752 27492
rect 28445 27489 28457 27492
rect 28491 27489 28503 27523
rect 28445 27483 28503 27489
rect 26605 27455 26663 27461
rect 26605 27452 26617 27455
rect 26200 27424 26617 27452
rect 26200 27412 26206 27424
rect 26605 27421 26617 27424
rect 26651 27421 26663 27455
rect 26605 27415 26663 27421
rect 26881 27455 26939 27461
rect 26881 27421 26893 27455
rect 26927 27421 26939 27455
rect 26881 27415 26939 27421
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 25648 27356 26004 27384
rect 25648 27344 25654 27356
rect 19794 27316 19800 27328
rect 14936 27288 19800 27316
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 21910 27276 21916 27328
rect 21968 27316 21974 27328
rect 22097 27319 22155 27325
rect 22097 27316 22109 27319
rect 21968 27288 22109 27316
rect 21968 27276 21974 27288
rect 22097 27285 22109 27288
rect 22143 27285 22155 27319
rect 22097 27279 22155 27285
rect 22370 27276 22376 27328
rect 22428 27316 22434 27328
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 22428 27288 22477 27316
rect 22428 27276 22434 27288
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 22465 27279 22523 27285
rect 25866 27276 25872 27328
rect 25924 27316 25930 27328
rect 26896 27316 26924 27415
rect 27522 27412 27528 27464
rect 27580 27412 27586 27464
rect 27706 27412 27712 27464
rect 27764 27412 27770 27464
rect 28353 27455 28411 27461
rect 28353 27421 28365 27455
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27421 28595 27455
rect 28537 27415 28595 27421
rect 29825 27455 29883 27461
rect 29825 27421 29837 27455
rect 29871 27452 29883 27455
rect 29914 27452 29920 27464
rect 29871 27424 29920 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 27540 27384 27568 27412
rect 28368 27384 28396 27415
rect 27540 27356 28396 27384
rect 25924 27288 26924 27316
rect 25924 27276 25930 27288
rect 27062 27276 27068 27328
rect 27120 27316 27126 27328
rect 27525 27319 27583 27325
rect 27525 27316 27537 27319
rect 27120 27288 27537 27316
rect 27120 27276 27126 27288
rect 27525 27285 27537 27288
rect 27571 27285 27583 27319
rect 28552 27316 28580 27415
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 30092 27387 30150 27393
rect 30092 27353 30104 27387
rect 30138 27384 30150 27387
rect 32214 27384 32220 27396
rect 30138 27356 32220 27384
rect 30138 27353 30150 27356
rect 30092 27347 30150 27353
rect 32214 27344 32220 27356
rect 32272 27344 32278 27396
rect 28718 27316 28724 27328
rect 28552 27288 28724 27316
rect 27525 27279 27583 27285
rect 28718 27276 28724 27288
rect 28776 27316 28782 27328
rect 31205 27319 31263 27325
rect 31205 27316 31217 27319
rect 28776 27288 31217 27316
rect 28776 27276 28782 27288
rect 31205 27285 31217 27288
rect 31251 27316 31263 27319
rect 32582 27316 32588 27328
rect 31251 27288 32588 27316
rect 31251 27285 31263 27288
rect 31205 27279 31263 27285
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12894 27112 12900 27124
rect 12124 27084 12900 27112
rect 12124 27072 12130 27084
rect 12894 27072 12900 27084
rect 12952 27072 12958 27124
rect 18230 27072 18236 27124
rect 18288 27112 18294 27124
rect 19521 27115 19579 27121
rect 19521 27112 19533 27115
rect 18288 27084 19533 27112
rect 18288 27072 18294 27084
rect 19521 27081 19533 27084
rect 19567 27081 19579 27115
rect 19521 27075 19579 27081
rect 19794 27072 19800 27124
rect 19852 27112 19858 27124
rect 19852 27084 22094 27112
rect 19852 27072 19858 27084
rect 8297 27047 8355 27053
rect 8297 27013 8309 27047
rect 8343 27044 8355 27047
rect 9122 27044 9128 27056
rect 8343 27016 9128 27044
rect 8343 27013 8355 27016
rect 8297 27007 8355 27013
rect 9122 27004 9128 27016
rect 9180 27044 9186 27056
rect 10594 27044 10600 27056
rect 9180 27016 10600 27044
rect 9180 27004 9186 27016
rect 10594 27004 10600 27016
rect 10652 27004 10658 27056
rect 12710 27044 12716 27056
rect 11900 27016 12716 27044
rect 8202 26936 8208 26988
rect 8260 26936 8266 26988
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 8527 26948 9229 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9217 26945 9229 26948
rect 9263 26976 9275 26979
rect 9766 26976 9772 26988
rect 9263 26948 9772 26976
rect 9263 26945 9275 26948
rect 9217 26939 9275 26945
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 11900 26985 11928 27016
rect 12710 27004 12716 27016
rect 12768 27044 12774 27056
rect 13446 27044 13452 27056
rect 12768 27016 13452 27044
rect 12768 27004 12774 27016
rect 13446 27004 13452 27016
rect 13504 27044 13510 27056
rect 13504 27016 13676 27044
rect 13504 27004 13510 27016
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 12066 26936 12072 26988
rect 12124 26936 12130 26988
rect 12161 26979 12219 26985
rect 12161 26945 12173 26979
rect 12207 26976 12219 26979
rect 12434 26976 12440 26988
rect 12207 26948 12440 26976
rect 12207 26945 12219 26948
rect 12161 26939 12219 26945
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 13648 26985 13676 27016
rect 14182 27004 14188 27056
rect 14240 27044 14246 27056
rect 15473 27047 15531 27053
rect 15473 27044 15485 27047
rect 14240 27016 15485 27044
rect 14240 27004 14246 27016
rect 15473 27013 15485 27016
rect 15519 27013 15531 27047
rect 22066 27044 22094 27084
rect 31110 27072 31116 27124
rect 31168 27072 31174 27124
rect 22649 27047 22707 27053
rect 22066 27016 22140 27044
rect 15473 27007 15531 27013
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26945 13691 26979
rect 13633 26939 13691 26945
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26976 15899 26979
rect 16390 26976 16396 26988
rect 15887 26948 16396 26976
rect 15887 26945 15899 26948
rect 15841 26939 15899 26945
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18322 26976 18328 26988
rect 18279 26948 18328 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 20898 26936 20904 26988
rect 20956 26976 20962 26988
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 20956 26948 21005 26976
rect 20956 26936 20962 26948
rect 20993 26945 21005 26948
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26945 21235 26979
rect 21177 26939 21235 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 21358 26976 21364 26988
rect 21315 26948 21364 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 8481 26843 8539 26849
rect 8481 26809 8493 26843
rect 8527 26840 8539 26843
rect 9048 26840 9076 26871
rect 9122 26868 9128 26920
rect 9180 26868 9186 26920
rect 9309 26911 9367 26917
rect 9309 26877 9321 26911
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 9324 26840 9352 26871
rect 8527 26812 9076 26840
rect 9140 26812 9352 26840
rect 21008 26840 21036 26939
rect 21192 26908 21220 26939
rect 21358 26936 21364 26948
rect 21416 26976 21422 26988
rect 22002 26976 22008 26988
rect 21416 26948 22008 26976
rect 21416 26936 21422 26948
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 22112 26985 22140 27016
rect 22649 27013 22661 27047
rect 22695 27044 22707 27047
rect 22922 27044 22928 27056
rect 22695 27016 22928 27044
rect 22695 27013 22707 27016
rect 22649 27007 22707 27013
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 22664 26908 22692 27007
rect 22922 27004 22928 27016
rect 22980 27044 22986 27056
rect 25406 27044 25412 27056
rect 22980 27016 25412 27044
rect 22980 27004 22986 27016
rect 25406 27004 25412 27016
rect 25464 27004 25470 27056
rect 26142 27044 26148 27056
rect 25792 27016 26148 27044
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 24820 26948 24961 26976
rect 24820 26936 24826 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 24949 26939 25007 26945
rect 25130 26936 25136 26988
rect 25188 26936 25194 26988
rect 25590 26936 25596 26988
rect 25648 26936 25654 26988
rect 25792 26985 25820 27016
rect 26142 27004 26148 27016
rect 26200 27044 26206 27056
rect 27525 27047 27583 27053
rect 27525 27044 27537 27047
rect 26200 27016 27537 27044
rect 26200 27004 26206 27016
rect 27525 27013 27537 27016
rect 27571 27013 27583 27047
rect 27525 27007 27583 27013
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 25866 26936 25872 26988
rect 25924 26936 25930 26988
rect 27246 26936 27252 26988
rect 27304 26936 27310 26988
rect 27430 26936 27436 26988
rect 27488 26936 27494 26988
rect 29822 26936 29828 26988
rect 29880 26976 29886 26988
rect 30009 26979 30067 26985
rect 30009 26976 30021 26979
rect 29880 26948 30021 26976
rect 29880 26936 29886 26948
rect 30009 26945 30021 26948
rect 30055 26945 30067 26979
rect 30009 26939 30067 26945
rect 21192 26880 22692 26908
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 26421 26911 26479 26917
rect 26421 26908 26433 26911
rect 26200 26880 26433 26908
rect 26200 26868 26206 26880
rect 26421 26877 26433 26880
rect 26467 26908 26479 26911
rect 28350 26908 28356 26920
rect 26467 26880 28356 26908
rect 26467 26877 26479 26880
rect 26421 26871 26479 26877
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 29733 26911 29791 26917
rect 29733 26877 29745 26911
rect 29779 26908 29791 26911
rect 29914 26908 29920 26920
rect 29779 26880 29920 26908
rect 29779 26877 29791 26880
rect 29733 26871 29791 26877
rect 29914 26868 29920 26880
rect 29972 26868 29978 26920
rect 21634 26840 21640 26852
rect 21008 26812 21640 26840
rect 8527 26809 8539 26812
rect 8481 26803 8539 26809
rect 8754 26732 8760 26784
rect 8812 26772 8818 26784
rect 9140 26772 9168 26812
rect 21634 26800 21640 26812
rect 21692 26800 21698 26852
rect 27154 26800 27160 26852
rect 27212 26840 27218 26852
rect 27522 26840 27528 26852
rect 27212 26812 27528 26840
rect 27212 26800 27218 26812
rect 27522 26800 27528 26812
rect 27580 26800 27586 26852
rect 8812 26744 9168 26772
rect 8812 26732 8818 26744
rect 9214 26732 9220 26784
rect 9272 26772 9278 26784
rect 9493 26775 9551 26781
rect 9493 26772 9505 26775
rect 9272 26744 9505 26772
rect 9272 26732 9278 26744
rect 9493 26741 9505 26744
rect 9539 26741 9551 26775
rect 9493 26735 9551 26741
rect 11146 26732 11152 26784
rect 11204 26772 11210 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 11204 26744 11713 26772
rect 11204 26732 11210 26744
rect 11701 26741 11713 26744
rect 11747 26741 11759 26775
rect 11701 26735 11759 26741
rect 12618 26732 12624 26784
rect 12676 26772 12682 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 12676 26744 13645 26772
rect 12676 26732 12682 26744
rect 13633 26741 13645 26744
rect 13679 26772 13691 26775
rect 18414 26772 18420 26784
rect 13679 26744 18420 26772
rect 13679 26741 13691 26744
rect 13633 26735 13691 26741
rect 18414 26732 18420 26744
rect 18472 26732 18478 26784
rect 20809 26775 20867 26781
rect 20809 26741 20821 26775
rect 20855 26772 20867 26775
rect 20898 26772 20904 26784
rect 20855 26744 20904 26772
rect 20855 26741 20867 26744
rect 20809 26735 20867 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12434 26568 12440 26580
rect 12391 26540 12440 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 13354 26568 13360 26580
rect 12952 26540 13360 26568
rect 12952 26528 12958 26540
rect 13354 26528 13360 26540
rect 13412 26568 13418 26580
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 13412 26540 13461 26568
rect 13412 26528 13418 26540
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 13449 26531 13507 26537
rect 15654 26528 15660 26580
rect 15712 26568 15718 26580
rect 16669 26571 16727 26577
rect 16669 26568 16681 26571
rect 15712 26540 16681 26568
rect 15712 26528 15718 26540
rect 16669 26537 16681 26540
rect 16715 26568 16727 26571
rect 17126 26568 17132 26580
rect 16715 26540 17132 26568
rect 16715 26537 16727 26540
rect 16669 26531 16727 26537
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 25130 26528 25136 26580
rect 25188 26568 25194 26580
rect 25225 26571 25283 26577
rect 25225 26568 25237 26571
rect 25188 26540 25237 26568
rect 25188 26528 25194 26540
rect 25225 26537 25237 26540
rect 25271 26537 25283 26571
rect 25225 26531 25283 26537
rect 27062 26528 27068 26580
rect 27120 26528 27126 26580
rect 32214 26528 32220 26580
rect 32272 26528 32278 26580
rect 9306 26460 9312 26512
rect 9364 26500 9370 26512
rect 9401 26503 9459 26509
rect 9401 26500 9413 26503
rect 9364 26472 9413 26500
rect 9364 26460 9370 26472
rect 9401 26469 9413 26472
rect 9447 26469 9459 26503
rect 13265 26503 13323 26509
rect 13265 26500 13277 26503
rect 9401 26463 9459 26469
rect 12084 26472 13277 26500
rect 11146 26392 11152 26444
rect 11204 26392 11210 26444
rect 11701 26435 11759 26441
rect 11701 26401 11713 26435
rect 11747 26432 11759 26435
rect 12084 26432 12112 26472
rect 13265 26469 13277 26472
rect 13311 26469 13323 26503
rect 13265 26463 13323 26469
rect 26694 26460 26700 26512
rect 26752 26500 26758 26512
rect 26752 26472 27752 26500
rect 26752 26460 26758 26472
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11747 26404 12112 26432
rect 12406 26404 12725 26432
rect 11747 26401 11759 26404
rect 11701 26395 11759 26401
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 12406 26364 12434 26404
rect 12713 26401 12725 26404
rect 12759 26432 12771 26435
rect 14734 26432 14740 26444
rect 12759 26404 14740 26432
rect 12759 26401 12771 26404
rect 12713 26395 12771 26401
rect 14734 26392 14740 26404
rect 14792 26392 14798 26444
rect 18049 26435 18107 26441
rect 18049 26401 18061 26435
rect 18095 26432 18107 26435
rect 18230 26432 18236 26444
rect 18095 26404 18236 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19392 26404 19840 26432
rect 19392 26392 19398 26404
rect 11379 26336 12434 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 12618 26324 12624 26376
rect 12676 26324 12682 26376
rect 19812 26373 19840 26404
rect 24578 26392 24584 26444
rect 24636 26432 24642 26444
rect 27724 26441 27752 26472
rect 28626 26460 28632 26512
rect 28684 26500 28690 26512
rect 31297 26503 31355 26509
rect 31297 26500 31309 26503
rect 28684 26472 31309 26500
rect 28684 26460 28690 26472
rect 31297 26469 31309 26472
rect 31343 26469 31355 26503
rect 31297 26463 31355 26469
rect 27709 26435 27767 26441
rect 24636 26404 27568 26432
rect 24636 26392 24642 26404
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 20070 26364 20076 26376
rect 19935 26336 20076 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 9030 26256 9036 26308
rect 9088 26296 9094 26308
rect 9125 26299 9183 26305
rect 9125 26296 9137 26299
rect 9088 26268 9137 26296
rect 9088 26256 9094 26268
rect 9125 26265 9137 26268
rect 9171 26296 9183 26299
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 9171 26268 11621 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 11609 26265 11621 26268
rect 11655 26265 11667 26299
rect 11609 26259 11667 26265
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13446 26305 13452 26308
rect 13417 26299 13452 26305
rect 13417 26296 13429 26299
rect 12584 26268 13429 26296
rect 12584 26256 12590 26268
rect 13417 26265 13429 26268
rect 13417 26259 13452 26265
rect 13446 26256 13452 26259
rect 13504 26256 13510 26308
rect 13538 26256 13544 26308
rect 13596 26296 13602 26308
rect 13633 26299 13691 26305
rect 13633 26296 13645 26299
rect 13596 26268 13645 26296
rect 13596 26256 13602 26268
rect 13633 26265 13645 26268
rect 13679 26265 13691 26299
rect 13633 26259 13691 26265
rect 16850 26256 16856 26308
rect 16908 26296 16914 26308
rect 17782 26299 17840 26305
rect 17782 26296 17794 26299
rect 16908 26268 17794 26296
rect 16908 26256 16914 26268
rect 17782 26265 17794 26268
rect 17828 26265 17840 26299
rect 17782 26259 17840 26265
rect 18230 26256 18236 26308
rect 18288 26296 18294 26308
rect 19429 26299 19487 26305
rect 19429 26296 19441 26299
rect 18288 26268 19441 26296
rect 18288 26256 18294 26268
rect 19429 26265 19441 26268
rect 19475 26265 19487 26299
rect 19628 26296 19656 26327
rect 20070 26324 20076 26336
rect 20128 26364 20134 26376
rect 21358 26364 21364 26376
rect 20128 26336 21364 26364
rect 20128 26324 20134 26336
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 25314 26324 25320 26376
rect 25372 26364 25378 26376
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 25372 26336 25421 26364
rect 25372 26324 25378 26336
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25498 26324 25504 26376
rect 25556 26324 25562 26376
rect 25590 26324 25596 26376
rect 25648 26324 25654 26376
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 25915 26336 26464 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 20254 26296 20260 26308
rect 19628 26268 20260 26296
rect 19429 26259 19487 26265
rect 20254 26256 20260 26268
rect 20312 26256 20318 26308
rect 22554 26256 22560 26308
rect 22612 26256 22618 26308
rect 22738 26256 22744 26308
rect 22796 26296 22802 26308
rect 25700 26296 25728 26327
rect 22796 26268 25728 26296
rect 22796 26256 22802 26268
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9585 26231 9643 26237
rect 9585 26228 9597 26231
rect 9364 26200 9597 26228
rect 9364 26188 9370 26200
rect 9585 26197 9597 26200
rect 9631 26197 9643 26231
rect 9585 26191 9643 26197
rect 21085 26231 21143 26237
rect 21085 26197 21097 26231
rect 21131 26228 21143 26231
rect 21174 26228 21180 26240
rect 21131 26200 21180 26228
rect 21131 26197 21143 26200
rect 21085 26191 21143 26197
rect 21174 26188 21180 26200
rect 21232 26188 21238 26240
rect 26436 26228 26464 26336
rect 26510 26324 26516 26376
rect 26568 26324 26574 26376
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26620 26296 26648 26327
rect 26786 26324 26792 26376
rect 26844 26324 26850 26376
rect 26878 26324 26884 26376
rect 26936 26324 26942 26376
rect 27540 26373 27568 26404
rect 27709 26401 27721 26435
rect 27755 26401 27767 26435
rect 27709 26395 27767 26401
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 32398 26324 32404 26376
rect 32456 26324 32462 26376
rect 32582 26324 32588 26376
rect 32640 26324 32646 26376
rect 32674 26324 32680 26376
rect 32732 26324 32738 26376
rect 27614 26296 27620 26308
rect 26620 26268 27620 26296
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 29086 26256 29092 26308
rect 29144 26296 29150 26308
rect 30009 26299 30067 26305
rect 30009 26296 30021 26299
rect 29144 26268 30021 26296
rect 29144 26256 29150 26268
rect 30009 26265 30021 26268
rect 30055 26265 30067 26299
rect 30009 26259 30067 26265
rect 26602 26228 26608 26240
rect 26436 26200 26608 26228
rect 26602 26188 26608 26200
rect 26660 26188 26666 26240
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 9272 25996 10640 26024
rect 9272 25984 9278 25996
rect 10505 25959 10563 25965
rect 10505 25956 10517 25959
rect 9508 25928 10517 25956
rect 9306 25848 9312 25900
rect 9364 25888 9370 25900
rect 9508 25897 9536 25928
rect 10505 25925 10517 25928
rect 10551 25925 10563 25959
rect 10505 25919 10563 25925
rect 9493 25891 9551 25897
rect 9493 25888 9505 25891
rect 9364 25860 9505 25888
rect 9364 25848 9370 25860
rect 9493 25857 9505 25860
rect 9539 25857 9551 25891
rect 9709 25891 9767 25897
rect 9709 25888 9721 25891
rect 9493 25851 9551 25857
rect 9692 25857 9721 25888
rect 9755 25857 9767 25891
rect 9692 25851 9767 25857
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25888 10471 25891
rect 10612 25888 10640 25996
rect 12342 25984 12348 26036
rect 12400 25984 12406 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12492 25996 13124 26024
rect 12492 25984 12498 25996
rect 12066 25916 12072 25968
rect 12124 25916 12130 25968
rect 12253 25959 12311 25965
rect 12253 25925 12265 25959
rect 12299 25956 12311 25959
rect 12526 25956 12532 25968
rect 12299 25928 12532 25956
rect 12299 25925 12311 25928
rect 12253 25919 12311 25925
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 13096 25965 13124 25996
rect 16850 25984 16856 26036
rect 16908 25984 16914 26036
rect 17126 25984 17132 26036
rect 17184 26024 17190 26036
rect 17221 26027 17279 26033
rect 17221 26024 17233 26027
rect 17184 25996 17233 26024
rect 17184 25984 17190 25996
rect 17221 25993 17233 25996
rect 17267 25993 17279 26027
rect 17221 25987 17279 25993
rect 25593 26027 25651 26033
rect 25593 25993 25605 26027
rect 25639 26024 25651 26027
rect 25682 26024 25688 26036
rect 25639 25996 25688 26024
rect 25639 25993 25651 25996
rect 25593 25987 25651 25993
rect 25682 25984 25688 25996
rect 25740 25984 25746 26036
rect 27157 26027 27215 26033
rect 27157 25993 27169 26027
rect 27203 26024 27215 26027
rect 27246 26024 27252 26036
rect 27203 25996 27252 26024
rect 27203 25993 27215 25996
rect 27157 25987 27215 25993
rect 27246 25984 27252 25996
rect 27304 25984 27310 26036
rect 29914 25984 29920 26036
rect 29972 25984 29978 26036
rect 13081 25959 13139 25965
rect 13081 25925 13093 25959
rect 13127 25925 13139 25959
rect 13081 25919 13139 25925
rect 13354 25916 13360 25968
rect 13412 25916 13418 25968
rect 21361 25959 21419 25965
rect 21361 25925 21373 25959
rect 21407 25956 21419 25959
rect 21910 25956 21916 25968
rect 21407 25928 21916 25956
rect 21407 25925 21419 25928
rect 21361 25919 21419 25925
rect 21910 25916 21916 25928
rect 21968 25916 21974 25968
rect 24581 25959 24639 25965
rect 24581 25925 24593 25959
rect 24627 25956 24639 25959
rect 25133 25959 25191 25965
rect 25133 25956 25145 25959
rect 24627 25928 25145 25956
rect 24627 25925 24639 25928
rect 24581 25919 24639 25925
rect 25133 25925 25145 25928
rect 25179 25956 25191 25959
rect 25498 25956 25504 25968
rect 25179 25928 25504 25956
rect 25179 25925 25191 25928
rect 25133 25919 25191 25925
rect 25498 25916 25504 25928
rect 25556 25916 25562 25968
rect 26786 25916 26792 25968
rect 26844 25956 26850 25968
rect 26844 25928 27568 25956
rect 26844 25916 26850 25928
rect 10459 25860 10640 25888
rect 10459 25857 10471 25860
rect 10413 25851 10471 25857
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9272 25792 9597 25820
rect 9272 25780 9278 25792
rect 9585 25789 9597 25792
rect 9631 25789 9643 25823
rect 9585 25783 9643 25789
rect 9692 25752 9720 25851
rect 10686 25848 10692 25900
rect 10744 25848 10750 25900
rect 12342 25848 12348 25900
rect 12400 25888 12406 25900
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 12400 25860 13277 25888
rect 12400 25848 12406 25860
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 9953 25823 10011 25829
rect 9953 25789 9965 25823
rect 9999 25820 10011 25823
rect 13280 25820 13308 25851
rect 13446 25848 13452 25900
rect 13504 25897 13510 25900
rect 13504 25888 13512 25897
rect 13504 25860 13549 25888
rect 13504 25851 13512 25860
rect 13504 25848 13510 25851
rect 17034 25848 17040 25900
rect 17092 25848 17098 25900
rect 17218 25848 17224 25900
rect 17276 25888 17282 25900
rect 17313 25891 17371 25897
rect 17313 25888 17325 25891
rect 17276 25860 17325 25888
rect 17276 25848 17282 25860
rect 17313 25857 17325 25860
rect 17359 25888 17371 25891
rect 17678 25888 17684 25900
rect 17359 25860 17684 25888
rect 17359 25857 17371 25860
rect 17313 25851 17371 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 19610 25848 19616 25900
rect 19668 25848 19674 25900
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 14642 25820 14648 25832
rect 9999 25792 12434 25820
rect 13280 25792 14648 25820
rect 9999 25789 10011 25792
rect 9953 25783 10011 25789
rect 10689 25755 10747 25761
rect 10689 25752 10701 25755
rect 9692 25724 10701 25752
rect 10689 25721 10701 25724
rect 10735 25721 10747 25755
rect 12406 25752 12434 25792
rect 14642 25780 14648 25792
rect 14700 25780 14706 25832
rect 14458 25752 14464 25764
rect 12406 25724 14464 25752
rect 10689 25715 10747 25721
rect 14458 25712 14464 25724
rect 14516 25712 14522 25764
rect 20824 25752 20852 25851
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21232 25860 22017 25888
rect 21232 25848 21238 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25888 22339 25891
rect 22370 25888 22376 25900
rect 22327 25860 22376 25888
rect 22327 25857 22339 25860
rect 22281 25851 22339 25857
rect 22370 25848 22376 25860
rect 22428 25848 22434 25900
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 24489 25891 24547 25897
rect 24489 25888 24501 25891
rect 23624 25860 24501 25888
rect 23624 25848 23630 25860
rect 24489 25857 24501 25860
rect 24535 25857 24547 25891
rect 24489 25851 24547 25857
rect 23474 25820 23480 25832
rect 21468 25792 23480 25820
rect 21468 25752 21496 25792
rect 23474 25780 23480 25792
rect 23532 25780 23538 25832
rect 24504 25820 24532 25851
rect 24670 25848 24676 25900
rect 24728 25888 24734 25900
rect 24854 25888 24860 25900
rect 24728 25860 24860 25888
rect 24728 25848 24734 25860
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 26510 25848 26516 25900
rect 26568 25848 26574 25900
rect 26878 25848 26884 25900
rect 26936 25888 26942 25900
rect 27540 25897 27568 25928
rect 27433 25891 27491 25897
rect 27433 25888 27445 25891
rect 26936 25860 27445 25888
rect 26936 25848 26942 25860
rect 27433 25857 27445 25860
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25857 27583 25891
rect 27525 25851 27583 25857
rect 28626 25848 28632 25900
rect 28684 25848 28690 25900
rect 31938 25848 31944 25900
rect 31996 25888 32002 25900
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31996 25860 32505 25888
rect 31996 25848 32002 25860
rect 32493 25857 32505 25860
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 32674 25848 32680 25900
rect 32732 25848 32738 25900
rect 32766 25848 32772 25900
rect 32824 25848 32830 25900
rect 25222 25820 25228 25832
rect 24504 25792 25228 25820
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 20824 25724 21496 25752
rect 25130 25712 25136 25764
rect 25188 25752 25194 25764
rect 25409 25755 25467 25761
rect 25409 25752 25421 25755
rect 25188 25724 25421 25752
rect 25188 25712 25194 25724
rect 25409 25721 25421 25724
rect 25455 25752 25467 25755
rect 26896 25752 26924 25848
rect 27062 25780 27068 25832
rect 27120 25820 27126 25832
rect 27341 25823 27399 25829
rect 27341 25820 27353 25823
rect 27120 25792 27353 25820
rect 27120 25780 27126 25792
rect 27341 25789 27353 25792
rect 27387 25789 27399 25823
rect 27341 25783 27399 25789
rect 27614 25780 27620 25832
rect 27672 25820 27678 25832
rect 28258 25820 28264 25832
rect 27672 25792 28264 25820
rect 27672 25780 27678 25792
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 25455 25724 26924 25752
rect 25455 25721 25467 25724
rect 25409 25715 25467 25721
rect 12621 25687 12679 25693
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 12710 25684 12716 25696
rect 12667 25656 12716 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 13078 25644 13084 25696
rect 13136 25644 13142 25696
rect 18322 25644 18328 25696
rect 18380 25644 18386 25696
rect 25866 25644 25872 25696
rect 25924 25684 25930 25696
rect 26050 25684 26056 25696
rect 25924 25656 26056 25684
rect 25924 25644 25930 25656
rect 26050 25644 26056 25656
rect 26108 25684 26114 25696
rect 26329 25687 26387 25693
rect 26329 25684 26341 25687
rect 26108 25656 26341 25684
rect 26108 25644 26114 25656
rect 26329 25653 26341 25656
rect 26375 25653 26387 25687
rect 26329 25647 26387 25653
rect 32306 25644 32312 25696
rect 32364 25644 32370 25696
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 15654 25480 15660 25492
rect 15427 25452 15660 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 15654 25440 15660 25452
rect 15712 25440 15718 25492
rect 19794 25440 19800 25492
rect 19852 25440 19858 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 26053 25483 26111 25489
rect 26053 25480 26065 25483
rect 25648 25452 26065 25480
rect 25648 25440 25654 25452
rect 26053 25449 26065 25452
rect 26099 25449 26111 25483
rect 26053 25443 26111 25449
rect 26237 25483 26295 25489
rect 26237 25449 26249 25483
rect 26283 25480 26295 25483
rect 26694 25480 26700 25492
rect 26283 25452 26700 25480
rect 26283 25449 26295 25452
rect 26237 25443 26295 25449
rect 26694 25440 26700 25452
rect 26752 25440 26758 25492
rect 28258 25440 28264 25492
rect 28316 25440 28322 25492
rect 13078 25344 13084 25356
rect 12544 25316 13084 25344
rect 3326 25236 3332 25288
rect 3384 25276 3390 25288
rect 3421 25279 3479 25285
rect 3421 25276 3433 25279
rect 3384 25248 3433 25276
rect 3384 25236 3390 25248
rect 3421 25245 3433 25248
rect 3467 25245 3479 25279
rect 3421 25239 3479 25245
rect 4062 25236 4068 25288
rect 4120 25236 4126 25288
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25276 4399 25279
rect 4798 25276 4804 25288
rect 4387 25248 4804 25276
rect 4387 25245 4399 25248
rect 4341 25239 4399 25245
rect 4798 25236 4804 25248
rect 4856 25236 4862 25288
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 6822 25276 6828 25288
rect 6779 25248 6828 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 6822 25236 6828 25248
rect 6880 25236 6886 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 7466 25276 7472 25288
rect 6963 25248 7472 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 7466 25236 7472 25248
rect 7524 25236 7530 25288
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 12544 25285 12572 25316
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 15672 25344 15700 25440
rect 16298 25372 16304 25424
rect 16356 25372 16362 25424
rect 26602 25372 26608 25424
rect 26660 25412 26666 25424
rect 26660 25384 28396 25412
rect 26660 25372 26666 25384
rect 15672 25316 16344 25344
rect 12253 25279 12311 25285
rect 12253 25276 12265 25279
rect 10744 25248 12265 25276
rect 10744 25236 10750 25248
rect 12253 25245 12265 25248
rect 12299 25276 12311 25279
rect 12529 25279 12587 25285
rect 12299 25248 12434 25276
rect 12299 25245 12311 25248
rect 12253 25239 12311 25245
rect 3970 25168 3976 25220
rect 4028 25168 4034 25220
rect 12406 25208 12434 25248
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12529 25239 12587 25245
rect 12710 25236 12716 25288
rect 12768 25236 12774 25288
rect 15378 25236 15384 25288
rect 15436 25236 15442 25288
rect 15930 25276 15936 25288
rect 15488 25248 15936 25276
rect 15396 25208 15424 25236
rect 12406 25180 15424 25208
rect 2866 25100 2872 25152
rect 2924 25140 2930 25152
rect 3329 25143 3387 25149
rect 3329 25140 3341 25143
rect 2924 25112 3341 25140
rect 2924 25100 2930 25112
rect 3329 25109 3341 25112
rect 3375 25109 3387 25143
rect 3329 25103 3387 25109
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 5592 25112 6745 25140
rect 5592 25100 5598 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6733 25103 6791 25109
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 13446 25140 13452 25152
rect 12115 25112 13452 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 15194 25100 15200 25152
rect 15252 25100 15258 25152
rect 15365 25143 15423 25149
rect 15365 25109 15377 25143
rect 15411 25140 15423 25143
rect 15488 25140 15516 25248
rect 15930 25236 15936 25248
rect 15988 25276 15994 25288
rect 16316 25285 16344 25316
rect 21174 25304 21180 25356
rect 21232 25304 21238 25356
rect 26206 25316 26740 25344
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15988 25248 16037 25276
rect 15988 25236 15994 25248
rect 16025 25245 16037 25248
rect 16071 25245 16083 25279
rect 16025 25239 16083 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 20898 25236 20904 25288
rect 20956 25285 20962 25288
rect 20956 25276 20968 25285
rect 20956 25248 21001 25276
rect 20956 25239 20968 25248
rect 20956 25236 20962 25239
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 26206 25276 26234 25316
rect 24872 25248 26234 25276
rect 26712 25276 26740 25316
rect 27338 25276 27344 25288
rect 26712 25248 27344 25276
rect 24872 25220 24900 25248
rect 27338 25236 27344 25248
rect 27396 25236 27402 25288
rect 28368 25285 28396 25384
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25276 28411 25279
rect 28902 25276 28908 25288
rect 28399 25248 28908 25276
rect 28399 25245 28411 25248
rect 28353 25239 28411 25245
rect 15565 25211 15623 25217
rect 15565 25177 15577 25211
rect 15611 25177 15623 25211
rect 15565 25171 15623 25177
rect 15411 25112 15516 25140
rect 15580 25140 15608 25171
rect 21082 25168 21088 25220
rect 21140 25208 21146 25220
rect 21637 25211 21695 25217
rect 21637 25208 21649 25211
rect 21140 25180 21649 25208
rect 21140 25168 21146 25180
rect 21637 25177 21649 25180
rect 21683 25177 21695 25211
rect 21637 25171 21695 25177
rect 24854 25168 24860 25220
rect 24912 25168 24918 25220
rect 25222 25168 25228 25220
rect 25280 25208 25286 25220
rect 26237 25211 26295 25217
rect 26237 25208 26249 25211
rect 25280 25180 26249 25208
rect 25280 25168 25286 25180
rect 26237 25177 26249 25180
rect 26283 25177 26295 25211
rect 26237 25171 26295 25177
rect 26510 25168 26516 25220
rect 26568 25208 26574 25220
rect 27448 25208 27476 25239
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 30098 25236 30104 25288
rect 30156 25236 30162 25288
rect 30374 25217 30380 25220
rect 26568 25180 27476 25208
rect 26568 25168 26574 25180
rect 15746 25140 15752 25152
rect 15580 25112 15752 25140
rect 15411 25109 15423 25112
rect 15365 25103 15423 25109
rect 15746 25100 15752 25112
rect 15804 25140 15810 25152
rect 16117 25143 16175 25149
rect 16117 25140 16129 25143
rect 15804 25112 16129 25140
rect 15804 25100 15810 25112
rect 16117 25109 16129 25112
rect 16163 25140 16175 25143
rect 18414 25140 18420 25152
rect 16163 25112 18420 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 18414 25100 18420 25112
rect 18472 25100 18478 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22612 25112 22937 25140
rect 22612 25100 22618 25112
rect 22925 25109 22937 25112
rect 22971 25109 22983 25143
rect 22925 25103 22983 25109
rect 27062 25100 27068 25152
rect 27120 25100 27126 25152
rect 27448 25140 27476 25180
rect 30368 25171 30380 25217
rect 30374 25168 30380 25171
rect 30432 25168 30438 25220
rect 30926 25140 30932 25152
rect 27448 25112 30932 25140
rect 30926 25100 30932 25112
rect 30984 25140 30990 25152
rect 31481 25143 31539 25149
rect 31481 25140 31493 25143
rect 30984 25112 31493 25140
rect 30984 25100 30990 25112
rect 31481 25109 31493 25112
rect 31527 25109 31539 25143
rect 31481 25103 31539 25109
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 17034 24896 17040 24948
rect 17092 24936 17098 24948
rect 17092 24908 23428 24936
rect 17092 24896 17098 24908
rect 5074 24828 5080 24880
rect 5132 24868 5138 24880
rect 5261 24871 5319 24877
rect 5261 24868 5273 24871
rect 5132 24840 5273 24868
rect 5132 24828 5138 24840
rect 5261 24837 5273 24840
rect 5307 24837 5319 24871
rect 5261 24831 5319 24837
rect 15212 24840 15884 24868
rect 15212 24812 15240 24840
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 2363 24772 3924 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24732 2651 24735
rect 2774 24732 2780 24744
rect 2639 24704 2780 24732
rect 2639 24701 2651 24704
rect 2593 24695 2651 24701
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 3896 24664 3924 24772
rect 3970 24760 3976 24812
rect 4028 24800 4034 24812
rect 4028 24772 4646 24800
rect 4028 24760 4034 24772
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 6917 24803 6975 24809
rect 6917 24800 6929 24803
rect 6880 24772 6929 24800
rect 6880 24760 6886 24772
rect 6917 24769 6929 24772
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 15013 24803 15071 24809
rect 15013 24769 15025 24803
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24800 15163 24803
rect 15194 24800 15200 24812
rect 15151 24772 15200 24800
rect 15151 24769 15163 24772
rect 15105 24763 15163 24769
rect 4706 24692 4712 24744
rect 4764 24692 4770 24744
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8386 24732 8392 24744
rect 7975 24704 8392 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 15028 24732 15056 24763
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15856 24809 15884 24840
rect 21100 24840 21404 24868
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16298 24800 16304 24812
rect 16071 24772 16304 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 15470 24732 15476 24744
rect 15028 24704 15476 24732
rect 15470 24692 15476 24704
rect 15528 24692 15534 24744
rect 6730 24664 6736 24676
rect 3896 24636 6736 24664
rect 6730 24624 6736 24636
rect 6788 24624 6794 24676
rect 15197 24667 15255 24673
rect 15197 24633 15209 24667
rect 15243 24664 15255 24667
rect 16040 24664 16068 24763
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 17678 24760 17684 24812
rect 17736 24800 17742 24812
rect 18141 24803 18199 24809
rect 17736 24772 18092 24800
rect 17736 24760 17742 24772
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17865 24735 17923 24741
rect 17865 24732 17877 24735
rect 17368 24704 17877 24732
rect 17368 24692 17374 24704
rect 17865 24701 17877 24704
rect 17911 24701 17923 24735
rect 18064 24732 18092 24772
rect 18141 24769 18153 24803
rect 18187 24800 18199 24803
rect 18230 24800 18236 24812
rect 18187 24772 18236 24800
rect 18187 24769 18199 24772
rect 18141 24763 18199 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 20806 24800 20812 24812
rect 18708 24772 20812 24800
rect 18708 24732 18736 24772
rect 20806 24760 20812 24772
rect 20864 24800 20870 24812
rect 21100 24809 21128 24840
rect 21376 24812 21404 24840
rect 20993 24803 21051 24809
rect 20993 24800 21005 24803
rect 20864 24772 21005 24800
rect 20864 24760 20870 24772
rect 20993 24769 21005 24772
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21085 24763 21143 24769
rect 21192 24772 21281 24800
rect 18064 24704 18736 24732
rect 17865 24695 17923 24701
rect 19334 24692 19340 24744
rect 19392 24692 19398 24744
rect 20898 24692 20904 24744
rect 20956 24732 20962 24744
rect 21192 24732 21220 24772
rect 21269 24769 21281 24772
rect 21315 24769 21327 24803
rect 21269 24763 21327 24769
rect 21358 24760 21364 24812
rect 21416 24760 21422 24812
rect 21453 24803 21511 24809
rect 21453 24769 21465 24803
rect 21499 24800 21511 24803
rect 22261 24803 22319 24809
rect 22261 24800 22273 24803
rect 21499 24772 22273 24800
rect 21499 24769 21511 24772
rect 21453 24763 21511 24769
rect 22261 24769 22273 24772
rect 22307 24769 22319 24803
rect 23400 24800 23428 24908
rect 25130 24896 25136 24948
rect 25188 24896 25194 24948
rect 27062 24868 27068 24880
rect 26160 24840 27068 24868
rect 23566 24800 23572 24812
rect 23400 24772 23572 24800
rect 22261 24763 22319 24769
rect 23566 24760 23572 24772
rect 23624 24760 23630 24812
rect 25222 24760 25228 24812
rect 25280 24760 25286 24812
rect 25314 24760 25320 24812
rect 25372 24760 25378 24812
rect 26160 24809 26188 24840
rect 27062 24828 27068 24840
rect 27120 24828 27126 24880
rect 28629 24871 28687 24877
rect 28629 24837 28641 24871
rect 28675 24837 28687 24871
rect 28629 24831 28687 24837
rect 28813 24871 28871 24877
rect 28813 24837 28825 24871
rect 28859 24837 28871 24871
rect 28813 24831 28871 24837
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24769 26203 24803
rect 28644 24800 28672 24831
rect 26145 24763 26203 24769
rect 26344 24772 28672 24800
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 20956 24704 21220 24732
rect 21284 24704 22017 24732
rect 20956 24692 20962 24704
rect 21284 24676 21312 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 26344 24732 26372 24772
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 28828 24800 28856 24831
rect 28776 24772 28856 24800
rect 28776 24760 28782 24772
rect 29086 24760 29092 24812
rect 29144 24760 29150 24812
rect 30368 24803 30426 24809
rect 30368 24769 30380 24803
rect 30414 24800 30426 24803
rect 32306 24800 32312 24812
rect 30414 24772 32312 24800
rect 30414 24769 30426 24772
rect 30368 24763 30426 24769
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 22005 24695 22063 24701
rect 23032 24704 26372 24732
rect 26421 24735 26479 24741
rect 15243 24636 16068 24664
rect 15243 24633 15255 24636
rect 15197 24627 15255 24633
rect 21266 24624 21272 24676
rect 21324 24624 21330 24676
rect 3881 24599 3939 24605
rect 3881 24565 3893 24599
rect 3927 24596 3939 24599
rect 4062 24596 4068 24608
rect 3927 24568 4068 24596
rect 3927 24565 3939 24568
rect 3881 24559 3939 24565
rect 4062 24556 4068 24568
rect 4120 24596 4126 24608
rect 4338 24596 4344 24608
rect 4120 24568 4344 24596
rect 4120 24556 4126 24568
rect 4338 24556 4344 24568
rect 4396 24556 4402 24608
rect 14918 24556 14924 24608
rect 14976 24596 14982 24608
rect 16025 24599 16083 24605
rect 16025 24596 16037 24599
rect 14976 24568 16037 24596
rect 14976 24556 14982 24568
rect 16025 24565 16037 24568
rect 16071 24565 16083 24599
rect 16025 24559 16083 24565
rect 21542 24556 21548 24608
rect 21600 24596 21606 24608
rect 23032 24596 23060 24704
rect 26421 24701 26433 24735
rect 26467 24732 26479 24735
rect 27154 24732 27160 24744
rect 26467 24704 27160 24732
rect 26467 24701 26479 24704
rect 26421 24695 26479 24701
rect 27154 24692 27160 24704
rect 27212 24692 27218 24744
rect 30098 24692 30104 24744
rect 30156 24692 30162 24744
rect 26329 24667 26387 24673
rect 26329 24633 26341 24667
rect 26375 24664 26387 24667
rect 26602 24664 26608 24676
rect 26375 24636 26608 24664
rect 26375 24633 26387 24636
rect 26329 24627 26387 24633
rect 26602 24624 26608 24636
rect 26660 24624 26666 24676
rect 31481 24667 31539 24673
rect 31481 24633 31493 24667
rect 31527 24664 31539 24667
rect 32674 24664 32680 24676
rect 31527 24636 32680 24664
rect 31527 24633 31539 24636
rect 31481 24627 31539 24633
rect 21600 24568 23060 24596
rect 23385 24599 23443 24605
rect 21600 24556 21606 24568
rect 23385 24565 23397 24599
rect 23431 24596 23443 24599
rect 23474 24596 23480 24608
rect 23431 24568 23480 24596
rect 23431 24565 23443 24568
rect 23385 24559 23443 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 25958 24556 25964 24608
rect 26016 24556 26022 24608
rect 28810 24556 28816 24608
rect 28868 24556 28874 24608
rect 28902 24556 28908 24608
rect 28960 24596 28966 24608
rect 31496 24596 31524 24627
rect 32674 24624 32680 24636
rect 32732 24624 32738 24676
rect 28960 24568 31524 24596
rect 28960 24556 28966 24568
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 2774 24352 2780 24404
rect 2832 24352 2838 24404
rect 6822 24352 6828 24404
rect 6880 24352 6886 24404
rect 20898 24392 20904 24404
rect 17880 24364 20904 24392
rect 2317 24327 2375 24333
rect 2317 24293 2329 24327
rect 2363 24324 2375 24327
rect 5261 24327 5319 24333
rect 5261 24324 5273 24327
rect 2363 24296 2912 24324
rect 2363 24293 2375 24296
rect 2317 24287 2375 24293
rect 2774 24256 2780 24268
rect 2056 24228 2780 24256
rect 2056 24197 2084 24228
rect 2774 24216 2780 24228
rect 2832 24216 2838 24268
rect 2041 24191 2099 24197
rect 2041 24157 2053 24191
rect 2087 24157 2099 24191
rect 2041 24151 2099 24157
rect 2314 24080 2320 24132
rect 2372 24080 2378 24132
rect 2884 24120 2912 24296
rect 2976 24296 5273 24324
rect 2976 24268 3004 24296
rect 5261 24293 5273 24296
rect 5307 24293 5319 24327
rect 5261 24287 5319 24293
rect 2958 24216 2964 24268
rect 3016 24216 3022 24268
rect 4157 24259 4215 24265
rect 4157 24256 4169 24259
rect 3068 24228 4169 24256
rect 3068 24197 3096 24228
rect 4157 24225 4169 24228
rect 4203 24225 4215 24259
rect 4157 24219 4215 24225
rect 4341 24259 4399 24265
rect 4341 24225 4353 24259
rect 4387 24256 4399 24259
rect 5074 24256 5080 24268
rect 4387 24228 5080 24256
rect 4387 24225 4399 24228
rect 4341 24219 4399 24225
rect 5074 24216 5080 24228
rect 5132 24256 5138 24268
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 5132 24228 5181 24256
rect 5132 24216 5138 24228
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 7282 24256 7288 24268
rect 5169 24219 5227 24225
rect 5460 24228 7288 24256
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 4433 24191 4491 24197
rect 4433 24157 4445 24191
rect 4479 24157 4491 24191
rect 4433 24151 4491 24157
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24157 4583 24191
rect 4525 24151 4583 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24188 4675 24191
rect 5460 24188 5488 24228
rect 7282 24216 7288 24228
rect 7340 24216 7346 24268
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 13504 24228 14780 24256
rect 13504 24216 13510 24228
rect 4663 24160 5488 24188
rect 4663 24157 4675 24160
rect 4617 24151 4675 24157
rect 3329 24123 3387 24129
rect 3329 24120 3341 24123
rect 2884 24092 3341 24120
rect 3329 24089 3341 24092
rect 3375 24089 3387 24123
rect 3329 24083 3387 24089
rect 3418 24080 3424 24132
rect 3476 24080 3482 24132
rect 2133 24055 2191 24061
rect 2133 24021 2145 24055
rect 2179 24052 2191 24055
rect 4246 24052 4252 24064
rect 2179 24024 4252 24052
rect 2179 24021 2191 24024
rect 2133 24015 2191 24021
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 4448 24052 4476 24151
rect 4540 24120 4568 24151
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24157 5779 24191
rect 5721 24151 5779 24157
rect 5552 24120 5580 24148
rect 4540 24092 5580 24120
rect 5736 24120 5764 24151
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7561 24191 7619 24197
rect 7561 24188 7573 24191
rect 7064 24160 7573 24188
rect 7064 24148 7070 24160
rect 7561 24157 7573 24160
rect 7607 24188 7619 24191
rect 8202 24188 8208 24200
rect 7607 24160 8208 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 8202 24148 8208 24160
rect 8260 24148 8266 24200
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24188 8539 24191
rect 9306 24188 9312 24200
rect 8527 24160 9312 24188
rect 8527 24157 8539 24160
rect 8481 24151 8539 24157
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 11974 24188 11980 24200
rect 11931 24160 11980 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24188 12127 24191
rect 12434 24188 12440 24200
rect 12115 24160 12440 24188
rect 12115 24157 12127 24160
rect 12069 24151 12127 24157
rect 12434 24148 12440 24160
rect 12492 24188 12498 24200
rect 13262 24188 13268 24200
rect 12492 24160 13268 24188
rect 12492 24148 12498 24160
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 7834 24120 7840 24132
rect 5736 24092 7840 24120
rect 5736 24052 5764 24092
rect 7834 24080 7840 24092
rect 7892 24080 7898 24132
rect 14476 24120 14504 24151
rect 14550 24148 14556 24200
rect 14608 24148 14614 24200
rect 14752 24197 14780 24228
rect 15010 24216 15016 24268
rect 15068 24256 15074 24268
rect 15841 24259 15899 24265
rect 15841 24256 15853 24259
rect 15068 24228 15853 24256
rect 15068 24216 15074 24228
rect 15841 24225 15853 24228
rect 15887 24225 15899 24259
rect 15841 24219 15899 24225
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 14826 24148 14832 24200
rect 14884 24148 14890 24200
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24157 15715 24191
rect 15657 24151 15715 24157
rect 15672 24120 15700 24151
rect 16390 24148 16396 24200
rect 16448 24188 16454 24200
rect 17880 24197 17908 24364
rect 20898 24352 20904 24364
rect 20956 24392 20962 24404
rect 21818 24392 21824 24404
rect 20956 24364 21824 24392
rect 20956 24352 20962 24364
rect 21818 24352 21824 24364
rect 21876 24392 21882 24404
rect 22833 24395 22891 24401
rect 21876 24364 22416 24392
rect 21876 24352 21882 24364
rect 22388 24324 22416 24364
rect 22833 24361 22845 24395
rect 22879 24392 22891 24395
rect 24578 24392 24584 24404
rect 22879 24364 24584 24392
rect 22879 24361 22891 24364
rect 22833 24355 22891 24361
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 30561 24395 30619 24401
rect 30561 24392 30573 24395
rect 30432 24364 30573 24392
rect 30432 24352 30438 24364
rect 30561 24361 30573 24364
rect 30607 24361 30619 24395
rect 30561 24355 30619 24361
rect 30006 24324 30012 24336
rect 22388 24296 30012 24324
rect 30006 24284 30012 24296
rect 30064 24284 30070 24336
rect 20993 24259 21051 24265
rect 20993 24225 21005 24259
rect 21039 24256 21051 24259
rect 21082 24256 21088 24268
rect 21039 24228 21088 24256
rect 21039 24225 21051 24228
rect 20993 24219 21051 24225
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 32398 24256 32404 24268
rect 23900 24228 32404 24256
rect 23900 24216 23906 24228
rect 32398 24216 32404 24228
rect 32456 24216 32462 24268
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16448 24160 17049 24188
rect 16448 24148 16454 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17865 24191 17923 24197
rect 17865 24157 17877 24191
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 17236 24120 17264 24151
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 18141 24191 18199 24197
rect 18141 24188 18153 24191
rect 18012 24160 18153 24188
rect 18012 24148 18018 24160
rect 18141 24157 18153 24160
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 20622 24148 20628 24200
rect 20680 24148 20686 24200
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 18049 24123 18107 24129
rect 18049 24120 18061 24123
rect 14476 24092 15608 24120
rect 15672 24092 17172 24120
rect 17236 24092 18061 24120
rect 4448 24024 5764 24052
rect 5810 24012 5816 24064
rect 5868 24052 5874 24064
rect 10502 24052 10508 24064
rect 5868 24024 10508 24052
rect 5868 24012 5874 24024
rect 10502 24012 10508 24024
rect 10560 24012 10566 24064
rect 12069 24055 12127 24061
rect 12069 24021 12081 24055
rect 12115 24052 12127 24055
rect 12618 24052 12624 24064
rect 12115 24024 12624 24052
rect 12115 24021 12127 24024
rect 12069 24015 12127 24021
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12894 24012 12900 24064
rect 12952 24052 12958 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 12952 24024 14289 24052
rect 12952 24012 12958 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 15470 24012 15476 24064
rect 15528 24012 15534 24064
rect 15580 24052 15608 24092
rect 17144 24064 17172 24092
rect 18049 24089 18061 24092
rect 18095 24120 18107 24123
rect 18690 24120 18696 24132
rect 18095 24092 18696 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18690 24080 18696 24092
rect 18748 24080 18754 24132
rect 19702 24080 19708 24132
rect 19760 24120 19766 24132
rect 20824 24120 20852 24151
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21324 24160 21465 24188
rect 21324 24148 21330 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 19760 24092 20852 24120
rect 21720 24123 21778 24129
rect 19760 24080 19766 24092
rect 21720 24089 21732 24123
rect 21766 24120 21778 24123
rect 23293 24123 23351 24129
rect 23293 24120 23305 24123
rect 21766 24092 23305 24120
rect 21766 24089 21778 24092
rect 21720 24083 21778 24089
rect 23293 24089 23305 24092
rect 23339 24089 23351 24123
rect 23768 24120 23796 24151
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 25866 24188 25872 24200
rect 25455 24160 25872 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 30834 24188 30840 24200
rect 30791 24160 30840 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 30834 24148 30840 24160
rect 30892 24148 30898 24200
rect 30926 24148 30932 24200
rect 30984 24148 30990 24200
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24188 31079 24191
rect 32766 24188 32772 24200
rect 31067 24160 32772 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 23293 24083 23351 24089
rect 23584 24092 23796 24120
rect 25240 24120 25268 24148
rect 25240 24092 25452 24120
rect 15654 24052 15660 24064
rect 15580 24024 15660 24052
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 17126 24012 17132 24064
rect 17184 24012 17190 24064
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 17644 24024 17693 24052
rect 17644 24012 17650 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 17681 24015 17739 24021
rect 20806 24012 20812 24064
rect 20864 24052 20870 24064
rect 23584 24052 23612 24092
rect 20864 24024 23612 24052
rect 20864 24012 20870 24024
rect 23658 24012 23664 24064
rect 23716 24012 23722 24064
rect 25314 24012 25320 24064
rect 25372 24012 25378 24064
rect 25424 24052 25452 24092
rect 25498 24080 25504 24132
rect 25556 24120 25562 24132
rect 31036 24120 31064 24151
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 25556 24092 31064 24120
rect 25556 24080 25562 24092
rect 26786 24052 26792 24064
rect 25424 24024 26792 24052
rect 26786 24012 26792 24024
rect 26844 24012 26850 24064
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 2314 23808 2320 23860
rect 2372 23848 2378 23860
rect 5077 23851 5135 23857
rect 5077 23848 5089 23851
rect 2372 23820 5089 23848
rect 2372 23808 2378 23820
rect 5077 23817 5089 23820
rect 5123 23817 5135 23851
rect 5077 23811 5135 23817
rect 5184 23820 7788 23848
rect 4617 23783 4675 23789
rect 4617 23749 4629 23783
rect 4663 23780 4675 23783
rect 4706 23780 4712 23792
rect 4663 23752 4712 23780
rect 4663 23749 4675 23752
rect 4617 23743 4675 23749
rect 4706 23740 4712 23752
rect 4764 23740 4770 23792
rect 4798 23740 4804 23792
rect 4856 23780 4862 23792
rect 5184 23780 5212 23820
rect 5810 23780 5816 23792
rect 4856 23752 5212 23780
rect 5276 23752 5816 23780
rect 4856 23740 4862 23752
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23712 3755 23715
rect 4522 23712 4528 23724
rect 3743 23684 4528 23712
rect 3743 23681 3755 23684
rect 3697 23675 3755 23681
rect 2792 23576 2820 23675
rect 4522 23672 4528 23684
rect 4580 23672 4586 23724
rect 5276 23653 5304 23752
rect 5810 23740 5816 23752
rect 5868 23740 5874 23792
rect 5445 23715 5503 23721
rect 5445 23681 5457 23715
rect 5491 23681 5503 23715
rect 5445 23675 5503 23681
rect 5537 23715 5595 23721
rect 5537 23681 5549 23715
rect 5583 23712 5595 23715
rect 7190 23712 7196 23724
rect 5583 23684 7196 23712
rect 5583 23681 5595 23684
rect 5537 23675 5595 23681
rect 5261 23647 5319 23653
rect 5261 23644 5273 23647
rect 3988 23616 5273 23644
rect 3326 23576 3332 23588
rect 2792 23548 3332 23576
rect 3326 23536 3332 23548
rect 3384 23576 3390 23588
rect 3988 23576 4016 23616
rect 5261 23613 5273 23616
rect 5307 23613 5319 23647
rect 5261 23607 5319 23613
rect 5353 23647 5411 23653
rect 5353 23613 5365 23647
rect 5399 23613 5411 23647
rect 5353 23607 5411 23613
rect 3384 23548 4016 23576
rect 3384 23536 3390 23548
rect 4338 23536 4344 23588
rect 4396 23576 4402 23588
rect 5368 23576 5396 23607
rect 4396 23548 5396 23576
rect 4396 23536 4402 23548
rect 4890 23468 4896 23520
rect 4948 23508 4954 23520
rect 5460 23508 5488 23675
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 7760 23712 7788 23820
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 15286 23848 15292 23860
rect 15151 23820 15292 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15286 23808 15292 23820
rect 15344 23848 15350 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15344 23820 15945 23848
rect 15344 23808 15350 23820
rect 15933 23817 15945 23820
rect 15979 23817 15991 23851
rect 15933 23811 15991 23817
rect 18230 23808 18236 23860
rect 18288 23848 18294 23860
rect 18414 23848 18420 23860
rect 18288 23820 18420 23848
rect 18288 23808 18294 23820
rect 18414 23808 18420 23820
rect 18472 23848 18478 23860
rect 21358 23848 21364 23860
rect 18472 23820 21364 23848
rect 18472 23808 18478 23820
rect 21358 23808 21364 23820
rect 21416 23848 21422 23860
rect 25222 23848 25228 23860
rect 21416 23820 25228 23848
rect 21416 23808 21422 23820
rect 8386 23740 8392 23792
rect 8444 23780 8450 23792
rect 8444 23752 9904 23780
rect 8444 23740 8450 23752
rect 9876 23721 9904 23752
rect 15010 23740 15016 23792
rect 15068 23780 15074 23792
rect 16117 23783 16175 23789
rect 16117 23780 16129 23783
rect 15068 23752 16129 23780
rect 15068 23740 15074 23752
rect 16117 23749 16129 23752
rect 16163 23749 16175 23783
rect 16117 23743 16175 23749
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23780 20039 23783
rect 20898 23780 20904 23792
rect 20027 23752 20904 23780
rect 20027 23749 20039 23752
rect 19981 23743 20039 23749
rect 20898 23740 20904 23752
rect 20956 23780 20962 23792
rect 21910 23780 21916 23792
rect 20956 23752 21916 23780
rect 20956 23740 20962 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22112 23789 22140 23820
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 30098 23808 30104 23860
rect 30156 23808 30162 23860
rect 22097 23783 22155 23789
rect 22097 23749 22109 23783
rect 22143 23749 22155 23783
rect 22097 23743 22155 23749
rect 28626 23740 28632 23792
rect 28684 23740 28690 23792
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 7760 23684 9229 23712
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10042 23672 10048 23724
rect 10100 23672 10106 23724
rect 12894 23672 12900 23724
rect 12952 23672 12958 23724
rect 13262 23672 13268 23724
rect 13320 23672 13326 23724
rect 14369 23715 14427 23721
rect 14369 23681 14381 23715
rect 14415 23712 14427 23715
rect 15470 23712 15476 23724
rect 14415 23684 15476 23712
rect 14415 23681 14427 23684
rect 14369 23675 14427 23681
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23712 16359 23715
rect 17126 23712 17132 23724
rect 16347 23684 17132 23712
rect 16347 23681 16359 23684
rect 16301 23675 16359 23681
rect 17126 23672 17132 23684
rect 17184 23672 17190 23724
rect 19518 23672 19524 23724
rect 19576 23712 19582 23724
rect 20441 23715 20499 23721
rect 20441 23712 20453 23715
rect 19576 23684 20453 23712
rect 19576 23672 19582 23684
rect 20441 23681 20453 23684
rect 20487 23681 20499 23715
rect 20441 23675 20499 23681
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6788 23616 6837 23644
rect 6788 23604 6794 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 7098 23604 7104 23656
rect 7156 23604 7162 23656
rect 8294 23604 8300 23656
rect 8352 23644 8358 23656
rect 8481 23647 8539 23653
rect 8481 23644 8493 23647
rect 8352 23616 8493 23644
rect 8352 23604 8358 23616
rect 8481 23613 8493 23616
rect 8527 23644 8539 23647
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 8527 23616 9413 23644
rect 8527 23613 8539 23616
rect 8481 23607 8539 23613
rect 9401 23613 9413 23616
rect 9447 23644 9459 23647
rect 9582 23644 9588 23656
rect 9447 23616 9588 23644
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 9582 23604 9588 23616
rect 9640 23604 9646 23656
rect 10502 23604 10508 23656
rect 10560 23644 10566 23656
rect 12253 23647 12311 23653
rect 12253 23644 12265 23647
rect 10560 23616 12265 23644
rect 10560 23604 10566 23616
rect 12253 23613 12265 23616
rect 12299 23613 12311 23647
rect 12253 23607 12311 23613
rect 12989 23647 13047 23653
rect 12989 23613 13001 23647
rect 13035 23613 13047 23647
rect 12989 23607 13047 23613
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 9953 23579 10011 23585
rect 9953 23576 9965 23579
rect 7892 23548 9965 23576
rect 7892 23536 7898 23548
rect 9953 23545 9965 23548
rect 9999 23545 10011 23579
rect 13004 23576 13032 23607
rect 13170 23604 13176 23656
rect 13228 23604 13234 23656
rect 14642 23604 14648 23656
rect 14700 23644 14706 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 14700 23616 14841 23644
rect 14700 23604 14706 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 14829 23607 14887 23613
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 15289 23647 15347 23653
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 15378 23644 15384 23656
rect 15335 23616 15384 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 15378 23604 15384 23616
rect 15436 23644 15442 23656
rect 16482 23644 16488 23656
rect 15436 23616 16488 23644
rect 15436 23604 15442 23616
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 14182 23576 14188 23588
rect 13004 23548 14188 23576
rect 9953 23539 10011 23545
rect 14182 23536 14188 23548
rect 14240 23536 14246 23588
rect 14277 23579 14335 23585
rect 14277 23545 14289 23579
rect 14323 23576 14335 23579
rect 15212 23576 15240 23604
rect 14323 23548 15240 23576
rect 18693 23579 18751 23585
rect 14323 23545 14335 23548
rect 14277 23539 14335 23545
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 19702 23576 19708 23588
rect 18739 23548 19708 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 20456 23576 20484 23675
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 21542 23712 21548 23724
rect 20772 23684 21548 23712
rect 20772 23672 20778 23684
rect 21542 23672 21548 23684
rect 21600 23672 21606 23724
rect 22649 23715 22707 23721
rect 22649 23681 22661 23715
rect 22695 23712 22707 23715
rect 23474 23712 23480 23724
rect 22695 23684 23480 23712
rect 22695 23681 22707 23684
rect 22649 23675 22707 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 23658 23672 23664 23724
rect 23716 23712 23722 23724
rect 24854 23712 24860 23724
rect 23716 23684 24860 23712
rect 23716 23672 23722 23684
rect 24854 23672 24860 23684
rect 24912 23712 24918 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 24912 23684 25513 23712
rect 24912 23672 24918 23684
rect 25501 23681 25513 23684
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 20806 23604 20812 23656
rect 20864 23604 20870 23656
rect 28810 23576 28816 23588
rect 20456 23548 28816 23576
rect 28810 23536 28816 23548
rect 28868 23536 28874 23588
rect 4948 23480 5488 23508
rect 4948 23468 4954 23480
rect 7466 23468 7472 23520
rect 7524 23508 7530 23520
rect 9033 23511 9091 23517
rect 9033 23508 9045 23511
rect 7524 23480 9045 23508
rect 7524 23468 7530 23480
rect 9033 23477 9045 23480
rect 9079 23477 9091 23511
rect 9033 23471 9091 23477
rect 15470 23468 15476 23520
rect 15528 23468 15534 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25409 23511 25467 23517
rect 25409 23508 25421 23511
rect 25004 23480 25421 23508
rect 25004 23468 25010 23480
rect 25409 23477 25421 23480
rect 25455 23477 25467 23511
rect 25409 23471 25467 23477
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3237 23307 3295 23313
rect 3237 23304 3249 23307
rect 2924 23276 3249 23304
rect 2924 23264 2930 23276
rect 3237 23273 3249 23276
rect 3283 23273 3295 23307
rect 3237 23267 3295 23273
rect 3329 23307 3387 23313
rect 3329 23273 3341 23307
rect 3375 23304 3387 23307
rect 3418 23304 3424 23316
rect 3375 23276 3424 23304
rect 3375 23273 3387 23276
rect 3329 23267 3387 23273
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 4157 23307 4215 23313
rect 4157 23273 4169 23307
rect 4203 23304 4215 23307
rect 4430 23304 4436 23316
rect 4203 23276 4436 23304
rect 4203 23273 4215 23276
rect 4157 23267 4215 23273
rect 4430 23264 4436 23276
rect 4488 23304 4494 23316
rect 4798 23304 4804 23316
rect 4488 23276 4804 23304
rect 4488 23264 4494 23276
rect 4798 23264 4804 23276
rect 4856 23264 4862 23316
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7098 23304 7104 23316
rect 6963 23276 7104 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 10318 23304 10324 23316
rect 8220 23276 10324 23304
rect 4890 23196 4896 23248
rect 4948 23236 4954 23248
rect 8220 23236 8248 23276
rect 10318 23264 10324 23276
rect 10376 23264 10382 23316
rect 11974 23264 11980 23316
rect 12032 23264 12038 23316
rect 18690 23264 18696 23316
rect 18748 23264 18754 23316
rect 21910 23264 21916 23316
rect 21968 23264 21974 23316
rect 31846 23264 31852 23316
rect 31904 23304 31910 23316
rect 33134 23304 33140 23316
rect 31904 23276 33140 23304
rect 31904 23264 31910 23276
rect 33134 23264 33140 23276
rect 33192 23264 33198 23316
rect 4948 23208 8248 23236
rect 4948 23196 4954 23208
rect 3421 23171 3479 23177
rect 3421 23137 3433 23171
rect 3467 23168 3479 23171
rect 3970 23168 3976 23180
rect 3467 23140 3976 23168
rect 3467 23137 3479 23140
rect 3421 23131 3479 23137
rect 3970 23128 3976 23140
rect 4028 23128 4034 23180
rect 8220 23177 8248 23208
rect 8662 23196 8668 23248
rect 8720 23236 8726 23248
rect 9125 23239 9183 23245
rect 9125 23236 9137 23239
rect 8720 23208 9137 23236
rect 8720 23196 8726 23208
rect 9125 23205 9137 23208
rect 9171 23205 9183 23239
rect 9125 23199 9183 23205
rect 8113 23171 8171 23177
rect 8113 23168 8125 23171
rect 7208 23140 8125 23168
rect 7208 23112 7236 23140
rect 8113 23137 8125 23140
rect 8159 23137 8171 23171
rect 8113 23131 8171 23137
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23137 8263 23171
rect 8205 23131 8263 23137
rect 8294 23128 8300 23180
rect 8352 23128 8358 23180
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23168 8447 23171
rect 8478 23168 8484 23180
rect 8435 23140 8484 23168
rect 8435 23137 8447 23140
rect 8389 23131 8447 23137
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 8573 23171 8631 23177
rect 8573 23137 8585 23171
rect 8619 23137 8631 23171
rect 8573 23131 8631 23137
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23168 11851 23171
rect 11992 23168 12020 23264
rect 15565 23239 15623 23245
rect 15565 23205 15577 23239
rect 15611 23236 15623 23239
rect 16117 23239 16175 23245
rect 16117 23236 16129 23239
rect 15611 23208 16129 23236
rect 15611 23205 15623 23208
rect 15565 23199 15623 23205
rect 16117 23205 16129 23208
rect 16163 23205 16175 23239
rect 16117 23199 16175 23205
rect 19610 23196 19616 23248
rect 19668 23236 19674 23248
rect 19705 23239 19763 23245
rect 19705 23236 19717 23239
rect 19668 23208 19717 23236
rect 19668 23196 19674 23208
rect 19705 23205 19717 23208
rect 19751 23205 19763 23239
rect 19705 23199 19763 23205
rect 19978 23196 19984 23248
rect 20036 23236 20042 23248
rect 28718 23236 28724 23248
rect 20036 23208 28724 23236
rect 20036 23196 20042 23208
rect 28718 23196 28724 23208
rect 28776 23196 28782 23248
rect 11839 23140 12020 23168
rect 11839 23137 11851 23140
rect 11793 23131 11851 23137
rect 3142 23060 3148 23112
rect 3200 23060 3206 23112
rect 7098 23060 7104 23112
rect 7156 23060 7162 23112
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 7558 23060 7564 23112
rect 7616 23060 7622 23112
rect 8588 23100 8616 23131
rect 14918 23128 14924 23180
rect 14976 23168 14982 23180
rect 15105 23171 15163 23177
rect 15105 23168 15117 23171
rect 14976 23140 15117 23168
rect 14976 23128 14982 23140
rect 15105 23137 15117 23140
rect 15151 23137 15163 23171
rect 15105 23131 15163 23137
rect 15194 23128 15200 23180
rect 15252 23128 15258 23180
rect 15286 23128 15292 23180
rect 15344 23128 15350 23180
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 15528 23140 16497 23168
rect 15528 23128 15534 23140
rect 16485 23137 16497 23140
rect 16531 23137 16543 23171
rect 16485 23131 16543 23137
rect 17310 23128 17316 23180
rect 17368 23128 17374 23180
rect 24946 23128 24952 23180
rect 25004 23128 25010 23180
rect 25314 23128 25320 23180
rect 25372 23128 25378 23180
rect 31386 23128 31392 23180
rect 31444 23168 31450 23180
rect 32674 23168 32680 23180
rect 31444 23140 32680 23168
rect 31444 23128 31450 23140
rect 32674 23128 32680 23140
rect 32732 23128 32738 23180
rect 33134 23128 33140 23180
rect 33192 23168 33198 23180
rect 33192 23140 33824 23168
rect 33192 23128 33198 23140
rect 8588 23072 8800 23100
rect 4338 22992 4344 23044
rect 4396 22992 4402 23044
rect 7285 23035 7343 23041
rect 7285 23001 7297 23035
rect 7331 23001 7343 23035
rect 7285 22995 7343 23001
rect 7423 23035 7481 23041
rect 7423 23001 7435 23035
rect 7469 23032 7481 23035
rect 8662 23032 8668 23044
rect 7469 23004 8668 23032
rect 7469 23001 7481 23004
rect 7423 22995 7481 23001
rect 3970 22924 3976 22976
rect 4028 22924 4034 22976
rect 4141 22967 4199 22973
rect 4141 22933 4153 22967
rect 4187 22964 4199 22967
rect 4706 22964 4712 22976
rect 4187 22936 4712 22964
rect 4187 22933 4199 22936
rect 4141 22927 4199 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 7300 22964 7328 22995
rect 8662 22992 8668 23004
rect 8720 22992 8726 23044
rect 8772 23032 8800 23072
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9364 23072 9413 23100
rect 9364 23060 9370 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 12066 23060 12072 23112
rect 12124 23060 12130 23112
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 12176 23072 12541 23100
rect 9125 23035 9183 23041
rect 9125 23032 9137 23035
rect 8772 23004 9137 23032
rect 9125 23001 9137 23004
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 9824 23004 10626 23032
rect 9824 22992 9830 23004
rect 11514 22992 11520 23044
rect 11572 23032 11578 23044
rect 12176 23032 12204 23072
rect 12529 23069 12541 23072
rect 12575 23069 12587 23103
rect 12529 23063 12587 23069
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 15010 23100 15016 23112
rect 14700 23072 15016 23100
rect 14700 23060 14706 23072
rect 15010 23060 15016 23072
rect 15068 23100 15074 23112
rect 17586 23109 17592 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15068 23072 15393 23100
rect 15068 23060 15074 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 17580 23100 17592 23109
rect 17547 23072 17592 23100
rect 15381 23063 15439 23069
rect 17580 23063 17592 23072
rect 17586 23060 17592 23063
rect 17644 23060 17650 23112
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 19702 23060 19708 23112
rect 19760 23060 19766 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20806 23100 20812 23112
rect 20671 23072 20812 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 24854 23060 24860 23112
rect 24912 23060 24918 23112
rect 27522 23060 27528 23112
rect 27580 23060 27586 23112
rect 28074 23060 28080 23112
rect 28132 23060 28138 23112
rect 28258 23060 28264 23112
rect 28316 23060 28322 23112
rect 31754 23060 31760 23112
rect 31812 23060 31818 23112
rect 32030 23060 32036 23112
rect 32088 23060 32094 23112
rect 32398 23060 32404 23112
rect 32456 23100 32462 23112
rect 32769 23103 32827 23109
rect 32769 23100 32781 23103
rect 32456 23072 32781 23100
rect 32456 23060 32462 23072
rect 32769 23069 32781 23072
rect 32815 23069 32827 23103
rect 32769 23063 32827 23069
rect 33318 23060 33324 23112
rect 33376 23100 33382 23112
rect 33796 23109 33824 23140
rect 33597 23103 33655 23109
rect 33597 23100 33609 23103
rect 33376 23072 33609 23100
rect 33376 23060 33382 23072
rect 33597 23069 33609 23072
rect 33643 23069 33655 23103
rect 33597 23063 33655 23069
rect 33781 23103 33839 23109
rect 33781 23069 33793 23103
rect 33827 23069 33839 23103
rect 33781 23063 33839 23069
rect 13265 23035 13323 23041
rect 13265 23032 13277 23035
rect 11572 23004 12204 23032
rect 12406 23004 13277 23032
rect 11572 22992 11578 23004
rect 7834 22964 7840 22976
rect 7300 22936 7840 22964
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 9309 22967 9367 22973
rect 9309 22964 9321 22967
rect 8260 22936 9321 22964
rect 8260 22924 8266 22936
rect 9309 22933 9321 22936
rect 9355 22964 9367 22967
rect 10226 22964 10232 22976
rect 9355 22936 10232 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 10410 22924 10416 22976
rect 10468 22964 10474 22976
rect 10870 22964 10876 22976
rect 10468 22936 10876 22964
rect 10468 22924 10474 22936
rect 10870 22924 10876 22936
rect 10928 22964 10934 22976
rect 12406 22964 12434 23004
rect 13265 23001 13277 23004
rect 13311 23001 13323 23035
rect 13265 22995 13323 23001
rect 24673 23035 24731 23041
rect 24673 23001 24685 23035
rect 24719 23032 24731 23035
rect 25314 23032 25320 23044
rect 24719 23004 25320 23032
rect 24719 23001 24731 23004
rect 24673 22995 24731 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 27614 22992 27620 23044
rect 27672 23032 27678 23044
rect 27801 23035 27859 23041
rect 27801 23032 27813 23035
rect 27672 23004 27813 23032
rect 27672 22992 27678 23004
rect 27801 23001 27813 23004
rect 27847 23001 27859 23035
rect 27801 22995 27859 23001
rect 10928 22936 12434 22964
rect 10928 22924 10934 22936
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 16025 22967 16083 22973
rect 16025 22964 16037 22967
rect 14700 22936 16037 22964
rect 14700 22924 14706 22936
rect 16025 22933 16037 22936
rect 16071 22933 16083 22967
rect 16025 22927 16083 22933
rect 25130 22924 25136 22976
rect 25188 22924 25194 22976
rect 25222 22924 25228 22976
rect 25280 22924 25286 22976
rect 29730 22924 29736 22976
rect 29788 22964 29794 22976
rect 31021 22967 31079 22973
rect 31021 22964 31033 22967
rect 29788 22936 31033 22964
rect 29788 22924 29794 22936
rect 31021 22933 31033 22936
rect 31067 22933 31079 22967
rect 31021 22927 31079 22933
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 33689 22967 33747 22973
rect 33689 22964 33701 22967
rect 33560 22936 33701 22964
rect 33560 22924 33566 22936
rect 33689 22933 33701 22936
rect 33735 22933 33747 22967
rect 33689 22927 33747 22933
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 7558 22760 7564 22772
rect 7239 22732 7564 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 10042 22760 10048 22772
rect 7892 22732 10048 22760
rect 7892 22720 7898 22732
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 8312 22701 8340 22732
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 31846 22760 31852 22772
rect 14568 22732 31852 22760
rect 8113 22695 8171 22701
rect 8113 22692 8125 22695
rect 7156 22664 8125 22692
rect 7156 22652 7162 22664
rect 8113 22661 8125 22664
rect 8159 22661 8171 22695
rect 8113 22655 8171 22661
rect 8297 22695 8355 22701
rect 8297 22661 8309 22695
rect 8343 22661 8355 22695
rect 8297 22655 8355 22661
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 8481 22695 8539 22701
rect 8481 22692 8493 22695
rect 8444 22664 8493 22692
rect 8444 22652 8450 22664
rect 8481 22661 8493 22664
rect 8527 22661 8539 22695
rect 8481 22655 8539 22661
rect 9306 22652 9312 22704
rect 9364 22692 9370 22704
rect 9677 22695 9735 22701
rect 9364 22664 9628 22692
rect 9364 22652 9370 22664
rect 4246 22584 4252 22636
rect 4304 22624 4310 22636
rect 4433 22627 4491 22633
rect 4433 22624 4445 22627
rect 4304 22596 4445 22624
rect 4304 22584 4310 22596
rect 4433 22593 4445 22596
rect 4479 22624 4491 22627
rect 7006 22624 7012 22636
rect 4479 22596 7012 22624
rect 4479 22593 4491 22596
rect 4433 22587 4491 22593
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7466 22624 7472 22636
rect 7423 22596 7472 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22593 9551 22627
rect 9600 22624 9628 22664
rect 9677 22661 9689 22695
rect 9723 22692 9735 22695
rect 9766 22692 9772 22704
rect 9723 22664 9772 22692
rect 9723 22661 9735 22664
rect 9677 22655 9735 22661
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 12529 22695 12587 22701
rect 12529 22692 12541 22695
rect 9876 22664 12541 22692
rect 9876 22624 9904 22664
rect 12529 22661 12541 22664
rect 12575 22661 12587 22695
rect 14369 22695 14427 22701
rect 14369 22692 14381 22695
rect 12529 22655 12587 22661
rect 13280 22664 14381 22692
rect 9600 22596 9904 22624
rect 10321 22627 10379 22633
rect 9493 22587 9551 22593
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 10410 22624 10416 22636
rect 10367 22596 10416 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 4522 22448 4528 22500
rect 4580 22488 4586 22500
rect 7576 22488 7604 22587
rect 7668 22556 7696 22587
rect 7668 22528 8524 22556
rect 8496 22500 8524 22528
rect 4580 22460 7604 22488
rect 4580 22448 4586 22460
rect 8478 22448 8484 22500
rect 8536 22448 8542 22500
rect 9416 22488 9444 22587
rect 9508 22556 9536 22587
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 11698 22584 11704 22636
rect 11756 22584 11762 22636
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 12434 22624 12440 22636
rect 11931 22596 12440 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 13280 22633 13308 22664
rect 14369 22661 14381 22664
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12676 22596 12909 22624
rect 12676 22584 12682 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 9508 22528 10977 22556
rect 10965 22525 10977 22528
rect 11011 22556 11023 22559
rect 11790 22556 11796 22568
rect 11011 22528 11796 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 11974 22488 11980 22500
rect 9416 22460 11980 22488
rect 11974 22448 11980 22460
rect 12032 22448 12038 22500
rect 12894 22448 12900 22500
rect 12952 22488 12958 22500
rect 13372 22488 13400 22587
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13504 22596 13645 22624
rect 13504 22584 13510 22596
rect 13633 22593 13645 22596
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 14568 22624 14596 22732
rect 31846 22720 31852 22732
rect 31904 22720 31910 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32401 22763 32459 22769
rect 32401 22760 32413 22763
rect 32088 22732 32413 22760
rect 32088 22720 32094 22732
rect 32401 22729 32413 22732
rect 32447 22729 32459 22763
rect 32401 22723 32459 22729
rect 15010 22652 15016 22704
rect 15068 22692 15074 22704
rect 18138 22692 18144 22704
rect 15068 22664 18144 22692
rect 15068 22652 15074 22664
rect 13955 22596 14596 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 15286 22584 15292 22636
rect 15344 22584 15350 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22593 15531 22627
rect 15473 22587 15531 22593
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22624 15623 22627
rect 15654 22624 15660 22636
rect 15611 22596 15660 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 14369 22559 14427 22565
rect 14369 22556 14381 22559
rect 14240 22528 14381 22556
rect 14240 22516 14246 22528
rect 14369 22525 14381 22528
rect 14415 22525 14427 22559
rect 15488 22556 15516 22587
rect 15654 22584 15660 22596
rect 15712 22624 15718 22636
rect 16298 22624 16304 22636
rect 15712 22596 16304 22624
rect 15712 22584 15718 22596
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 17126 22584 17132 22636
rect 17184 22624 17190 22636
rect 17512 22633 17540 22664
rect 18138 22652 18144 22664
rect 18196 22652 18202 22704
rect 18601 22695 18659 22701
rect 18601 22661 18613 22695
rect 18647 22692 18659 22695
rect 18690 22692 18696 22704
rect 18647 22664 18696 22692
rect 18647 22661 18659 22664
rect 18601 22655 18659 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 20162 22652 20168 22704
rect 20220 22692 20226 22704
rect 20622 22692 20628 22704
rect 20220 22664 20628 22692
rect 20220 22652 20226 22664
rect 20622 22652 20628 22664
rect 20680 22692 20686 22704
rect 23753 22695 23811 22701
rect 20680 22664 23704 22692
rect 20680 22652 20686 22664
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 17184 22596 17325 22624
rect 17184 22584 17190 22596
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22593 17555 22627
rect 19978 22624 19984 22636
rect 17497 22587 17555 22593
rect 18064 22596 19984 22624
rect 15930 22556 15936 22568
rect 15488 22528 15936 22556
rect 14369 22519 14427 22525
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 16316 22556 16344 22584
rect 18064 22556 18092 22596
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22624 20407 22627
rect 20530 22624 20536 22636
rect 20395 22596 20536 22624
rect 20395 22593 20407 22596
rect 20349 22587 20407 22593
rect 16316 22528 18092 22556
rect 18138 22516 18144 22568
rect 18196 22516 18202 22568
rect 18230 22516 18236 22568
rect 18288 22516 18294 22568
rect 12952 22460 13400 22488
rect 17405 22491 17463 22497
rect 12952 22448 12958 22460
rect 17405 22457 17417 22491
rect 17451 22488 17463 22491
rect 18046 22488 18052 22500
rect 17451 22460 18052 22488
rect 17451 22457 17463 22460
rect 17405 22451 17463 22457
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 18156 22488 18184 22516
rect 20088 22488 20116 22587
rect 18156 22460 20116 22488
rect 20272 22488 20300 22587
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 22020 22633 22048 22664
rect 23676 22633 23704 22664
rect 23753 22661 23765 22695
rect 23799 22692 23811 22695
rect 25222 22692 25228 22704
rect 23799 22664 25228 22692
rect 23799 22661 23811 22664
rect 23753 22655 23811 22661
rect 25222 22652 25228 22664
rect 25280 22652 25286 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 27672 22664 29960 22692
rect 27672 22652 27678 22664
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22624 22063 22627
rect 22189 22627 22247 22633
rect 22051 22596 22085 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22624 24915 22627
rect 27154 22624 27160 22636
rect 24903 22596 27160 22624
rect 24903 22593 24915 22596
rect 24857 22587 24915 22593
rect 22005 22491 22063 22497
rect 22005 22488 22017 22491
rect 20272 22460 22017 22488
rect 22005 22457 22017 22460
rect 22051 22457 22063 22491
rect 22204 22488 22232 22587
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 28166 22584 28172 22636
rect 28224 22584 28230 22636
rect 28258 22584 28264 22636
rect 28316 22624 28322 22636
rect 29932 22633 29960 22664
rect 28813 22627 28871 22633
rect 28813 22624 28825 22627
rect 28316 22596 28825 22624
rect 28316 22584 28322 22596
rect 28813 22593 28825 22596
rect 28859 22624 28871 22627
rect 29917 22627 29975 22633
rect 28859 22596 29868 22624
rect 28859 22593 28871 22596
rect 28813 22587 28871 22593
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 23900 22528 24777 22556
rect 23900 22516 23906 22528
rect 24765 22525 24777 22528
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 25133 22559 25191 22565
rect 25133 22525 25145 22559
rect 25179 22556 25191 22559
rect 26142 22556 26148 22568
rect 25179 22528 26148 22556
rect 25179 22525 25191 22528
rect 25133 22519 25191 22525
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 29730 22516 29736 22568
rect 29788 22516 29794 22568
rect 25774 22488 25780 22500
rect 22204 22460 25780 22488
rect 22005 22451 22063 22457
rect 25774 22448 25780 22460
rect 25832 22448 25838 22500
rect 27982 22448 27988 22500
rect 28040 22488 28046 22500
rect 29748 22488 29776 22516
rect 28040 22460 29776 22488
rect 29840 22488 29868 22596
rect 29917 22593 29929 22627
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 30101 22627 30159 22633
rect 30101 22593 30113 22627
rect 30147 22624 30159 22627
rect 31297 22627 31355 22633
rect 31297 22624 31309 22627
rect 30147 22596 31309 22624
rect 30147 22593 30159 22596
rect 30101 22587 30159 22593
rect 31297 22593 31309 22596
rect 31343 22593 31355 22627
rect 31297 22587 31355 22593
rect 31021 22559 31079 22565
rect 31021 22525 31033 22559
rect 31067 22525 31079 22559
rect 31021 22519 31079 22525
rect 31036 22488 31064 22519
rect 31110 22516 31116 22568
rect 31168 22516 31174 22568
rect 31202 22516 31208 22568
rect 31260 22516 31266 22568
rect 32048 22488 32076 22720
rect 33045 22695 33103 22701
rect 33045 22661 33057 22695
rect 33091 22692 33103 22695
rect 33134 22692 33140 22704
rect 33091 22664 33140 22692
rect 33091 22661 33103 22664
rect 33045 22655 33103 22661
rect 33134 22652 33140 22664
rect 33192 22652 33198 22704
rect 33502 22652 33508 22704
rect 33560 22652 33566 22704
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 33686 22584 33692 22636
rect 33744 22584 33750 22636
rect 32398 22516 32404 22568
rect 32456 22556 32462 22568
rect 32539 22559 32597 22565
rect 32539 22556 32551 22559
rect 32456 22528 32551 22556
rect 32456 22516 32462 22528
rect 32539 22525 32551 22528
rect 32585 22525 32597 22559
rect 32539 22519 32597 22525
rect 32953 22559 33011 22565
rect 32953 22525 32965 22559
rect 32999 22556 33011 22559
rect 33318 22556 33324 22568
rect 32999 22528 33324 22556
rect 32999 22525 33011 22528
rect 32953 22519 33011 22525
rect 33318 22516 33324 22528
rect 33376 22516 33382 22568
rect 29840 22460 30972 22488
rect 31036 22460 32076 22488
rect 28040 22448 28046 22460
rect 4338 22380 4344 22432
rect 4396 22420 4402 22432
rect 9214 22420 9220 22432
rect 4396 22392 9220 22420
rect 4396 22380 4402 22392
rect 9214 22380 9220 22392
rect 9272 22380 9278 22432
rect 10226 22380 10232 22432
rect 10284 22420 10290 22432
rect 10410 22420 10416 22432
rect 10284 22392 10416 22420
rect 10284 22380 10290 22392
rect 10410 22380 10416 22392
rect 10468 22380 10474 22432
rect 11793 22423 11851 22429
rect 11793 22389 11805 22423
rect 11839 22420 11851 22423
rect 12986 22420 12992 22432
rect 11839 22392 12992 22420
rect 11839 22389 11851 22392
rect 11793 22383 11851 22389
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 14553 22423 14611 22429
rect 14553 22389 14565 22423
rect 14599 22420 14611 22423
rect 15105 22423 15163 22429
rect 15105 22420 15117 22423
rect 14599 22392 15117 22420
rect 14599 22389 14611 22392
rect 14553 22383 14611 22389
rect 15105 22389 15117 22392
rect 15151 22389 15163 22423
rect 15105 22383 15163 22389
rect 17954 22380 17960 22432
rect 18012 22380 18018 22432
rect 19794 22380 19800 22432
rect 19852 22380 19858 22432
rect 24578 22380 24584 22432
rect 24636 22380 24642 22432
rect 26970 22380 26976 22432
rect 27028 22420 27034 22432
rect 27341 22423 27399 22429
rect 27341 22420 27353 22423
rect 27028 22392 27353 22420
rect 27028 22380 27034 22392
rect 27341 22389 27353 22392
rect 27387 22389 27399 22423
rect 27341 22383 27399 22389
rect 30834 22380 30840 22432
rect 30892 22380 30898 22432
rect 30944 22420 30972 22460
rect 33781 22423 33839 22429
rect 33781 22420 33793 22423
rect 30944 22392 33793 22420
rect 33781 22389 33793 22392
rect 33827 22389 33839 22423
rect 33781 22383 33839 22389
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 4982 22176 4988 22228
rect 5040 22216 5046 22228
rect 11514 22216 11520 22228
rect 5040 22188 11520 22216
rect 5040 22176 5046 22188
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 11698 22176 11704 22228
rect 11756 22225 11762 22228
rect 11756 22219 11771 22225
rect 11759 22185 11771 22219
rect 11756 22179 11771 22185
rect 11756 22176 11762 22179
rect 15286 22176 15292 22228
rect 15344 22216 15350 22228
rect 15344 22188 22094 22216
rect 15344 22176 15350 22188
rect 12434 22108 12440 22160
rect 12492 22148 12498 22160
rect 12809 22151 12867 22157
rect 12809 22148 12821 22151
rect 12492 22120 12821 22148
rect 12492 22108 12498 22120
rect 12809 22117 12821 22120
rect 12855 22117 12867 22151
rect 12809 22111 12867 22117
rect 17954 22108 17960 22160
rect 18012 22108 18018 22160
rect 19242 22108 19248 22160
rect 19300 22148 19306 22160
rect 21634 22148 21640 22160
rect 19300 22120 21640 22148
rect 19300 22108 19306 22120
rect 21634 22108 21640 22120
rect 21692 22108 21698 22160
rect 22066 22148 22094 22188
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 23201 22219 23259 22225
rect 23201 22216 23213 22219
rect 22704 22188 23213 22216
rect 22704 22176 22710 22188
rect 23201 22185 23213 22188
rect 23247 22185 23259 22219
rect 23201 22179 23259 22185
rect 33505 22219 33563 22225
rect 33505 22185 33517 22219
rect 33551 22216 33563 22219
rect 33686 22216 33692 22228
rect 33551 22188 33692 22216
rect 33551 22185 33563 22188
rect 33505 22179 33563 22185
rect 33686 22176 33692 22188
rect 33744 22176 33750 22228
rect 23017 22151 23075 22157
rect 23017 22148 23029 22151
rect 22066 22120 23029 22148
rect 23017 22117 23029 22120
rect 23063 22117 23075 22151
rect 30374 22148 30380 22160
rect 23017 22111 23075 22117
rect 24964 22120 25360 22148
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 10229 22083 10287 22089
rect 10229 22080 10241 22083
rect 3200 22052 10241 22080
rect 3200 22040 3206 22052
rect 10229 22049 10241 22052
rect 10275 22080 10287 22083
rect 11054 22080 11060 22092
rect 10275 22052 11060 22080
rect 10275 22049 10287 22052
rect 10229 22043 10287 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11664 22052 11989 22080
rect 11664 22040 11670 22052
rect 11977 22049 11989 22052
rect 12023 22080 12035 22083
rect 12066 22080 12072 22092
rect 12023 22052 12072 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 17773 22083 17831 22089
rect 17773 22049 17785 22083
rect 17819 22080 17831 22083
rect 17972 22080 18000 22108
rect 24964 22080 24992 22120
rect 17819 22052 18000 22080
rect 18064 22052 24992 22080
rect 25041 22083 25099 22089
rect 17819 22049 17831 22052
rect 17773 22043 17831 22049
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 7156 21984 7205 22012
rect 7156 21972 7162 21984
rect 7193 21981 7205 21984
rect 7239 22012 7251 22015
rect 7466 22012 7472 22024
rect 7239 21984 7472 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9306 22012 9312 22024
rect 8619 21984 9312 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 11698 21944 11704 21956
rect 11270 21916 11704 21944
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 12728 21944 12756 21975
rect 12894 21972 12900 22024
rect 12952 21972 12958 22024
rect 12986 21972 12992 22024
rect 13044 21972 13050 22024
rect 17954 21972 17960 22024
rect 18012 21972 18018 22024
rect 18064 21944 18092 22052
rect 25041 22049 25053 22083
rect 25087 22080 25099 22083
rect 25222 22080 25228 22092
rect 25087 22052 25228 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 25332 22080 25360 22120
rect 26896 22120 27108 22148
rect 26896 22080 26924 22120
rect 25332 22052 26924 22080
rect 26970 22040 26976 22092
rect 27028 22040 27034 22092
rect 27080 22080 27108 22120
rect 30024 22120 30380 22148
rect 29914 22080 29920 22092
rect 27080 22052 29920 22080
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 30024 22089 30052 22120
rect 30374 22108 30380 22120
rect 30432 22148 30438 22160
rect 30834 22148 30840 22160
rect 30432 22120 30840 22148
rect 30432 22108 30438 22120
rect 30834 22108 30840 22120
rect 30892 22108 30898 22160
rect 30009 22083 30067 22089
rect 30009 22049 30021 22083
rect 30055 22080 30067 22083
rect 30055 22052 30089 22080
rect 31404 22052 32628 22080
rect 30055 22049 30067 22052
rect 30009 22043 30067 22049
rect 18230 21972 18236 22024
rect 18288 21972 18294 22024
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 19426 22012 19432 22024
rect 18371 21984 19432 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 18340 21944 18368 21975
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 22012 20867 22015
rect 20898 22012 20904 22024
rect 20855 21984 20904 22012
rect 20855 21981 20867 21984
rect 20809 21975 20867 21981
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23201 22015 23259 22021
rect 23201 22012 23213 22015
rect 22980 21984 23213 22012
rect 22980 21972 22986 21984
rect 23201 21981 23213 21984
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 22012 23443 22015
rect 24578 22012 24584 22024
rect 23431 21984 24584 22012
rect 23431 21981 23443 21984
rect 23385 21975 23443 21981
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24762 21972 24768 22024
rect 24820 21972 24826 22024
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 25958 22012 25964 22024
rect 24995 21984 25964 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 12728 21916 18092 21944
rect 18156 21916 18368 21944
rect 7190 21836 7196 21888
rect 7248 21836 7254 21888
rect 8478 21836 8484 21888
rect 8536 21836 8542 21888
rect 10686 21836 10692 21888
rect 10744 21876 10750 21888
rect 12529 21879 12587 21885
rect 12529 21876 12541 21879
rect 10744 21848 12541 21876
rect 10744 21836 10750 21848
rect 12529 21845 12541 21848
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 16482 21836 16488 21888
rect 16540 21876 16546 21888
rect 18156 21876 18184 21916
rect 19610 21904 19616 21956
rect 19668 21944 19674 21956
rect 19797 21947 19855 21953
rect 19797 21944 19809 21947
rect 19668 21916 19809 21944
rect 19668 21904 19674 21916
rect 19797 21913 19809 21916
rect 19843 21913 19855 21947
rect 19797 21907 19855 21913
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21944 20223 21947
rect 20254 21944 20260 21956
rect 20211 21916 20260 21944
rect 20211 21913 20223 21916
rect 20165 21907 20223 21913
rect 20254 21904 20260 21916
rect 20312 21944 20318 21956
rect 21082 21944 21088 21956
rect 20312 21916 21088 21944
rect 20312 21904 20318 21916
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 24872 21944 24900 21975
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 21981 26111 22015
rect 26053 21975 26111 21981
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 26988 22012 27016 22040
rect 26283 21984 27016 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 25130 21944 25136 21956
rect 24872 21916 25136 21944
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 16540 21848 18184 21876
rect 16540 21836 16546 21848
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 25096 21848 25237 21876
rect 25096 21836 25102 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 26068 21876 26096 21975
rect 27062 21972 27068 22024
rect 27120 22012 27126 22024
rect 27249 22015 27307 22021
rect 27249 22012 27261 22015
rect 27120 21984 27261 22012
rect 27120 21972 27126 21984
rect 27249 21981 27261 21984
rect 27295 22012 27307 22015
rect 27338 22012 27344 22024
rect 27295 21984 27344 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 27847 21984 28641 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 28629 21981 28641 21984
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 21981 30159 22015
rect 30101 21975 30159 21981
rect 26145 21947 26203 21953
rect 26145 21913 26157 21947
rect 26191 21944 26203 21947
rect 27522 21944 27528 21956
rect 26191 21916 27528 21944
rect 26191 21913 26203 21916
rect 26145 21907 26203 21913
rect 27522 21904 27528 21916
rect 27580 21944 27586 21956
rect 28261 21947 28319 21953
rect 28261 21944 28273 21947
rect 27580 21916 28273 21944
rect 27580 21904 27586 21916
rect 28261 21913 28273 21916
rect 28307 21913 28319 21947
rect 28261 21907 28319 21913
rect 28442 21904 28448 21956
rect 28500 21904 28506 21956
rect 30116 21944 30144 21975
rect 31018 21972 31024 22024
rect 31076 21972 31082 22024
rect 31202 21972 31208 22024
rect 31260 22012 31266 22024
rect 31404 22021 31432 22052
rect 32600 22024 32628 22052
rect 33134 22040 33140 22092
rect 33192 22040 33198 22092
rect 31389 22015 31447 22021
rect 31389 22012 31401 22015
rect 31260 21984 31401 22012
rect 31260 21972 31266 21984
rect 31389 21981 31401 21984
rect 31435 21981 31447 22015
rect 31389 21975 31447 21981
rect 31570 21972 31576 22024
rect 31628 22012 31634 22024
rect 32033 22015 32091 22021
rect 32033 22012 32045 22015
rect 31628 21984 32045 22012
rect 31628 21972 31634 21984
rect 32033 21981 32045 21984
rect 32079 21981 32091 22015
rect 32033 21975 32091 21981
rect 32398 21972 32404 22024
rect 32456 21972 32462 22024
rect 32582 21972 32588 22024
rect 32640 21972 32646 22024
rect 33318 21972 33324 22024
rect 33376 21972 33382 22024
rect 30282 21944 30288 21956
rect 30116 21916 30288 21944
rect 30282 21904 30288 21916
rect 30340 21944 30346 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30340 21916 31125 21944
rect 30340 21904 30346 21916
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 32125 21947 32183 21953
rect 32125 21944 32137 21947
rect 31113 21907 31171 21913
rect 31726 21916 32137 21944
rect 26970 21876 26976 21888
rect 26068 21848 26976 21876
rect 25225 21839 25283 21845
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 27062 21836 27068 21888
rect 27120 21876 27126 21888
rect 27709 21879 27767 21885
rect 27709 21876 27721 21879
rect 27120 21848 27721 21876
rect 27120 21836 27126 21848
rect 27709 21845 27721 21848
rect 27755 21845 27767 21879
rect 27709 21839 27767 21845
rect 29730 21836 29736 21888
rect 29788 21836 29794 21888
rect 31018 21836 31024 21888
rect 31076 21876 31082 21888
rect 31726 21876 31754 21916
rect 32125 21913 32137 21916
rect 32171 21913 32183 21947
rect 32125 21907 32183 21913
rect 31076 21848 31754 21876
rect 31076 21836 31082 21848
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 9858 21632 9864 21684
rect 9916 21672 9922 21684
rect 27062 21672 27068 21684
rect 9916 21644 12434 21672
rect 9916 21632 9922 21644
rect 11698 21564 11704 21616
rect 11756 21564 11762 21616
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 2915 21508 3801 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 3789 21505 3801 21508
rect 3835 21536 3847 21539
rect 3970 21536 3976 21548
rect 3835 21508 3976 21536
rect 3835 21505 3847 21508
rect 3789 21499 3847 21505
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21536 4123 21539
rect 4522 21536 4528 21548
rect 4111 21508 4528 21536
rect 4111 21505 4123 21508
rect 4065 21499 4123 21505
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 11790 21496 11796 21548
rect 11848 21496 11854 21548
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12406 21536 12434 21644
rect 22066 21644 27068 21672
rect 22066 21604 22094 21644
rect 27062 21632 27068 21644
rect 27120 21632 27126 21684
rect 27154 21632 27160 21684
rect 27212 21632 27218 21684
rect 29086 21672 29092 21684
rect 28092 21644 29092 21672
rect 28092 21604 28120 21644
rect 29086 21632 29092 21644
rect 29144 21632 29150 21684
rect 30282 21632 30288 21684
rect 30340 21632 30346 21684
rect 31665 21675 31723 21681
rect 31665 21641 31677 21675
rect 31711 21672 31723 21675
rect 31754 21672 31760 21684
rect 31711 21644 31760 21672
rect 31711 21641 31723 21644
rect 31665 21635 31723 21641
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 28442 21604 28448 21616
rect 20548 21576 22094 21604
rect 24596 21576 28120 21604
rect 28184 21576 28448 21604
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 12406 21508 14473 21536
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14599 21508 15301 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15838 21536 15844 21548
rect 15519 21508 15844 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 15838 21496 15844 21508
rect 15896 21536 15902 21548
rect 17678 21536 17684 21548
rect 15896 21508 17684 21536
rect 15896 21496 15902 21508
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 19518 21496 19524 21548
rect 19576 21496 19582 21548
rect 19794 21496 19800 21548
rect 19852 21496 19858 21548
rect 20548 21545 20576 21576
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 2958 21428 2964 21480
rect 3016 21428 3022 21480
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21468 3203 21471
rect 3191 21440 4016 21468
rect 3191 21437 3203 21440
rect 3145 21431 3203 21437
rect 2976 21400 3004 21428
rect 3988 21409 4016 21440
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 20640 21468 20668 21499
rect 18288 21440 20668 21468
rect 18288 21428 18294 21440
rect 3881 21403 3939 21409
rect 3881 21400 3893 21403
rect 2976 21372 3893 21400
rect 3881 21369 3893 21372
rect 3927 21369 3939 21403
rect 3881 21363 3939 21369
rect 3973 21403 4031 21409
rect 3973 21369 3985 21403
rect 4019 21400 4031 21403
rect 4062 21400 4068 21412
rect 4019 21372 4068 21400
rect 4019 21369 4031 21372
rect 3973 21363 4031 21369
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 22020 21400 22048 21499
rect 22278 21496 22284 21548
rect 22336 21496 22342 21548
rect 22370 21428 22376 21480
rect 22428 21428 22434 21480
rect 23198 21428 23204 21480
rect 23256 21428 23262 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 23566 21468 23572 21480
rect 23523 21440 23572 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24596 21477 24624 21576
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 27982 21536 27988 21548
rect 27571 21508 27988 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 28184 21545 28212 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 30374 21604 30380 21616
rect 30208 21576 30380 21604
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 29730 21536 29736 21548
rect 28399 21508 29736 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23992 21440 24593 21468
rect 23992 21428 23998 21440
rect 24581 21437 24593 21440
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 27433 21471 27491 21477
rect 27433 21437 27445 21471
rect 27479 21468 27491 21471
rect 27614 21468 27620 21480
rect 27479 21440 27620 21468
rect 27479 21437 27491 21440
rect 27433 21431 27491 21437
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 28184 21400 28212 21499
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 30208 21545 30236 21576
rect 30374 21564 30380 21576
rect 30432 21564 30438 21616
rect 30469 21607 30527 21613
rect 30469 21573 30481 21607
rect 30515 21604 30527 21607
rect 31018 21604 31024 21616
rect 30515 21576 31024 21604
rect 30515 21573 30527 21576
rect 30469 21567 30527 21573
rect 31018 21564 31024 21576
rect 31076 21564 31082 21616
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21505 30251 21539
rect 30193 21499 30251 21505
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31481 21539 31539 21545
rect 31481 21536 31493 21539
rect 31168 21508 31493 21536
rect 31168 21496 31174 21508
rect 31481 21505 31493 21508
rect 31527 21505 31539 21539
rect 31481 21499 31539 21505
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21536 31723 21539
rect 32582 21536 32588 21548
rect 31711 21508 32588 21536
rect 31711 21505 31723 21508
rect 31665 21499 31723 21505
rect 32582 21496 32588 21508
rect 32640 21496 32646 21548
rect 19208 21372 22094 21400
rect 19208 21360 19214 21372
rect 3050 21292 3056 21344
rect 3108 21292 3114 21344
rect 3602 21292 3608 21344
rect 3660 21292 3666 21344
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 16666 21332 16672 21344
rect 15519 21304 16672 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 16666 21292 16672 21304
rect 16724 21292 16730 21344
rect 19426 21292 19432 21344
rect 19484 21292 19490 21344
rect 22066 21332 22094 21372
rect 24504 21372 28212 21400
rect 23842 21332 23848 21344
rect 22066 21304 23848 21332
rect 23842 21292 23848 21304
rect 23900 21332 23906 21344
rect 24504 21332 24532 21372
rect 23900 21304 24532 21332
rect 23900 21292 23906 21304
rect 27890 21292 27896 21344
rect 27948 21332 27954 21344
rect 28353 21335 28411 21341
rect 28353 21332 28365 21335
rect 27948 21304 28365 21332
rect 27948 21292 27954 21304
rect 28353 21301 28365 21304
rect 28399 21301 28411 21335
rect 28353 21295 28411 21301
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 30469 21335 30527 21341
rect 30469 21332 30481 21335
rect 28500 21304 30481 21332
rect 28500 21292 28506 21304
rect 30469 21301 30481 21304
rect 30515 21301 30527 21335
rect 30469 21295 30527 21301
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 12952 21100 13461 21128
rect 12952 21088 12958 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21097 14795 21131
rect 14737 21091 14795 21097
rect 16117 21131 16175 21137
rect 16117 21097 16129 21131
rect 16163 21128 16175 21131
rect 17310 21128 17316 21140
rect 16163 21100 17316 21128
rect 16163 21097 16175 21100
rect 16117 21091 16175 21097
rect 14752 21060 14780 21091
rect 17310 21088 17316 21100
rect 17368 21088 17374 21140
rect 21266 21088 21272 21140
rect 21324 21088 21330 21140
rect 23566 21088 23572 21140
rect 23624 21088 23630 21140
rect 23842 21088 23848 21140
rect 23900 21128 23906 21140
rect 31938 21128 31944 21140
rect 23900 21100 31944 21128
rect 23900 21088 23906 21100
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 32398 21088 32404 21140
rect 32456 21088 32462 21140
rect 25866 21060 25872 21072
rect 14752 21032 25872 21060
rect 25866 21020 25872 21032
rect 25924 21020 25930 21072
rect 31110 21020 31116 21072
rect 31168 21060 31174 21072
rect 31297 21063 31355 21069
rect 31297 21060 31309 21063
rect 31168 21032 31309 21060
rect 31168 21020 31174 21032
rect 31297 21029 31309 21032
rect 31343 21029 31355 21063
rect 31297 21023 31355 21029
rect 4522 20952 4528 21004
rect 4580 20992 4586 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 4580 20964 7389 20992
rect 4580 20952 4586 20964
rect 7377 20961 7389 20964
rect 7423 20992 7435 20995
rect 7466 20992 7472 21004
rect 7423 20964 7472 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 11882 20992 11888 21004
rect 10612 20964 11888 20992
rect 3234 20884 3240 20936
rect 3292 20884 3298 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 3510 20924 3516 20936
rect 3467 20896 3516 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 3510 20884 3516 20896
rect 3568 20884 3574 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7340 20896 7573 20924
rect 7340 20884 7346 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 7650 20884 7656 20936
rect 7708 20884 7714 20936
rect 10410 20884 10416 20936
rect 10468 20884 10474 20936
rect 10612 20933 10640 20964
rect 11882 20952 11888 20964
rect 11940 20992 11946 21004
rect 19426 20992 19432 21004
rect 11940 20964 19432 20992
rect 11940 20952 11946 20964
rect 19426 20952 19432 20964
rect 19484 20952 19490 21004
rect 19978 20952 19984 21004
rect 20036 20992 20042 21004
rect 20073 20995 20131 21001
rect 20073 20992 20085 20995
rect 20036 20964 20085 20992
rect 20036 20952 20042 20964
rect 20073 20961 20085 20964
rect 20119 20961 20131 20995
rect 20073 20955 20131 20961
rect 20165 20995 20223 21001
rect 20165 20961 20177 20995
rect 20211 20992 20223 20995
rect 21174 20992 21180 21004
rect 20211 20964 21180 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 28442 20992 28448 21004
rect 22066 20964 28448 20992
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20893 10655 20927
rect 10597 20887 10655 20893
rect 10686 20884 10692 20936
rect 10744 20884 10750 20936
rect 13446 20884 13452 20936
rect 13504 20924 13510 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13504 20896 13553 20924
rect 13504 20884 13510 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 14516 20896 14565 20924
rect 14516 20884 14522 20896
rect 14553 20893 14565 20896
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20924 17463 20927
rect 18322 20924 18328 20936
rect 17451 20896 18328 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 14752 20856 14780 20887
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19705 20927 19763 20933
rect 19705 20924 19717 20927
rect 19208 20896 19717 20924
rect 19208 20884 19214 20896
rect 19705 20893 19717 20896
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 22066 20924 22094 20964
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 33045 20995 33103 21001
rect 33045 20992 33057 20995
rect 31680 20964 33057 20992
rect 19843 20896 22094 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 22554 20884 22560 20936
rect 22612 20884 22618 20936
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23308 20896 23765 20924
rect 14752 20828 19564 20856
rect 3142 20748 3148 20800
rect 3200 20788 3206 20800
rect 3329 20791 3387 20797
rect 3329 20788 3341 20791
rect 3200 20760 3341 20788
rect 3200 20748 3206 20760
rect 3329 20757 3341 20760
rect 3375 20757 3387 20791
rect 3329 20751 3387 20757
rect 7374 20748 7380 20800
rect 7432 20748 7438 20800
rect 10226 20748 10232 20800
rect 10284 20748 10290 20800
rect 14366 20748 14372 20800
rect 14424 20748 14430 20800
rect 19536 20797 19564 20828
rect 21358 20816 21364 20868
rect 21416 20856 21422 20868
rect 21634 20856 21640 20868
rect 21416 20828 21640 20856
rect 21416 20816 21422 20828
rect 21634 20816 21640 20828
rect 21692 20856 21698 20868
rect 23308 20856 23336 20896
rect 23753 20893 23765 20896
rect 23799 20924 23811 20927
rect 23842 20924 23848 20936
rect 23799 20896 23848 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 23934 20884 23940 20936
rect 23992 20884 23998 20936
rect 24026 20884 24032 20936
rect 24084 20884 24090 20936
rect 24765 20927 24823 20933
rect 24765 20923 24777 20927
rect 24688 20895 24777 20923
rect 21692 20828 23336 20856
rect 21692 20816 21698 20828
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 23440 20828 24593 20856
rect 23440 20816 23446 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24581 20819 24639 20825
rect 24688 20856 24716 20895
rect 24765 20893 24777 20895
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24946 20884 24952 20936
rect 25004 20924 25010 20936
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 25004 20896 25053 20924
rect 25004 20884 25010 20896
rect 25041 20893 25053 20896
rect 25087 20924 25099 20927
rect 25130 20924 25136 20936
rect 25087 20896 25136 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25130 20884 25136 20896
rect 25188 20924 25194 20936
rect 25498 20924 25504 20936
rect 25188 20896 25504 20924
rect 25188 20884 25194 20896
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 31680 20933 31708 20964
rect 33045 20961 33057 20964
rect 33091 20961 33103 20995
rect 33045 20955 33103 20961
rect 31572 20927 31630 20933
rect 31572 20893 31584 20927
rect 31618 20893 31630 20927
rect 31572 20887 31630 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 30926 20856 30932 20868
rect 24688 20828 30932 20856
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 21082 20748 21088 20800
rect 21140 20788 21146 20800
rect 24688 20788 24716 20828
rect 30926 20816 30932 20828
rect 30984 20816 30990 20868
rect 31588 20856 31616 20887
rect 32122 20884 32128 20936
rect 32180 20924 32186 20936
rect 32217 20927 32275 20933
rect 32217 20924 32229 20927
rect 32180 20896 32229 20924
rect 32180 20884 32186 20896
rect 32217 20893 32229 20896
rect 32263 20893 32275 20927
rect 32217 20887 32275 20893
rect 32306 20884 32312 20936
rect 32364 20924 32370 20936
rect 32401 20927 32459 20933
rect 32401 20924 32413 20927
rect 32364 20896 32413 20924
rect 32364 20884 32370 20896
rect 32401 20893 32413 20896
rect 32447 20893 32459 20927
rect 32401 20887 32459 20893
rect 32950 20884 32956 20936
rect 33008 20884 33014 20936
rect 33137 20927 33195 20933
rect 33137 20924 33149 20927
rect 33060 20896 33149 20924
rect 33060 20868 33088 20896
rect 33137 20893 33149 20896
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 32766 20856 32772 20868
rect 31588 20828 32772 20856
rect 32766 20816 32772 20828
rect 32824 20816 32830 20868
rect 33042 20816 33048 20868
rect 33100 20816 33106 20868
rect 21140 20760 24716 20788
rect 21140 20748 21146 20760
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 7834 20544 7840 20596
rect 7892 20544 7898 20596
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20553 8447 20587
rect 14182 20584 14188 20596
rect 8389 20547 8447 20553
rect 13372 20556 14188 20584
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 3418 20516 3424 20528
rect 3108 20488 3424 20516
rect 3108 20476 3114 20488
rect 3418 20476 3424 20488
rect 3476 20516 3482 20528
rect 3513 20519 3571 20525
rect 3513 20516 3525 20519
rect 3476 20488 3525 20516
rect 3476 20476 3482 20488
rect 3513 20485 3525 20488
rect 3559 20485 3571 20519
rect 3513 20479 3571 20485
rect 3602 20476 3608 20528
rect 3660 20476 3666 20528
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 7742 20516 7748 20528
rect 7515 20488 7748 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 7742 20476 7748 20488
rect 7800 20516 7806 20528
rect 8404 20516 8432 20547
rect 7800 20488 8432 20516
rect 7800 20476 7806 20488
rect 3142 20408 3148 20460
rect 3200 20408 3206 20460
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3970 20448 3976 20460
rect 3283 20420 3976 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 5074 20448 5080 20460
rect 4479 20420 5080 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7340 20420 7389 20448
rect 7340 20408 7346 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 8018 20448 8024 20460
rect 7699 20420 8024 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20349 4399 20383
rect 8312 20380 8340 20411
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 8481 20451 8539 20457
rect 8481 20448 8493 20451
rect 8444 20420 8493 20448
rect 8444 20408 8450 20420
rect 8481 20417 8493 20420
rect 8527 20417 8539 20451
rect 8481 20411 8539 20417
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 10226 20448 10232 20460
rect 8619 20420 10232 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13372 20448 13400 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 19521 20587 19579 20593
rect 19521 20553 19533 20587
rect 19567 20584 19579 20587
rect 19886 20584 19892 20596
rect 19567 20556 19892 20584
rect 19567 20553 19579 20556
rect 19521 20547 19579 20553
rect 19886 20544 19892 20556
rect 19944 20584 19950 20596
rect 20898 20584 20904 20596
rect 19944 20556 20904 20584
rect 19944 20544 19950 20556
rect 20898 20544 20904 20556
rect 20956 20544 20962 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 24854 20584 24860 20596
rect 21131 20556 24860 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 31570 20544 31576 20596
rect 31628 20544 31634 20596
rect 32582 20544 32588 20596
rect 32640 20544 32646 20596
rect 14366 20516 14372 20528
rect 13464 20488 14372 20516
rect 13464 20457 13492 20488
rect 14366 20476 14372 20488
rect 14424 20476 14430 20528
rect 15562 20516 15568 20528
rect 14476 20488 15568 20516
rect 13311 20420 13400 20448
rect 13449 20451 13507 20457
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13449 20411 13507 20417
rect 13556 20420 13829 20448
rect 9030 20380 9036 20392
rect 8312 20352 9036 20380
rect 4341 20343 4399 20349
rect 2406 20272 2412 20324
rect 2464 20312 2470 20324
rect 4356 20312 4384 20343
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 10410 20340 10416 20392
rect 10468 20340 10474 20392
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13556 20380 13584 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 14476 20448 14504 20488
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 21358 20516 21364 20528
rect 19352 20488 21364 20516
rect 14047 20420 14504 20448
rect 15105 20451 15163 20457
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15151 20420 15608 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 13412 20352 13584 20380
rect 13412 20340 13418 20352
rect 2464 20284 4384 20312
rect 2464 20272 2470 20284
rect 12802 20272 12808 20324
rect 12860 20312 12866 20324
rect 14016 20312 14044 20411
rect 14182 20340 14188 20392
rect 14240 20380 14246 20392
rect 14829 20383 14887 20389
rect 14829 20380 14841 20383
rect 14240 20352 14841 20380
rect 14240 20340 14246 20352
rect 14829 20349 14841 20352
rect 14875 20380 14887 20383
rect 14918 20380 14924 20392
rect 14875 20352 14924 20380
rect 14875 20349 14887 20352
rect 14829 20343 14887 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 12860 20284 14044 20312
rect 12860 20272 12866 20284
rect 14090 20272 14096 20324
rect 14148 20312 14154 20324
rect 15120 20312 15148 20411
rect 14148 20284 15148 20312
rect 15580 20312 15608 20420
rect 15654 20408 15660 20460
rect 15712 20408 15718 20460
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 19352 20457 19380 20488
rect 21358 20476 21364 20488
rect 21416 20476 21422 20528
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 23201 20519 23259 20525
rect 23201 20516 23213 20519
rect 22428 20488 23213 20516
rect 22428 20476 22434 20488
rect 23201 20485 23213 20488
rect 23247 20485 23259 20519
rect 23201 20479 23259 20485
rect 29086 20476 29092 20528
rect 29144 20516 29150 20528
rect 32122 20516 32128 20528
rect 29144 20488 32128 20516
rect 29144 20476 29150 20488
rect 32122 20476 32128 20488
rect 32180 20476 32186 20528
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20417 19395 20451
rect 19337 20411 19395 20417
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 20070 20448 20076 20460
rect 19659 20420 20076 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 20548 20380 20576 20411
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 20717 20451 20775 20457
rect 20717 20448 20729 20451
rect 20680 20420 20729 20448
rect 20680 20408 20686 20420
rect 20717 20417 20729 20420
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21266 20448 21272 20460
rect 20947 20420 21272 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 19306 20352 20576 20380
rect 20824 20380 20852 20411
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 27890 20408 27896 20460
rect 27948 20408 27954 20460
rect 27982 20408 27988 20460
rect 28040 20408 28046 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 32490 20448 32496 20460
rect 31803 20420 32496 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 20990 20380 20996 20392
rect 20824 20352 20996 20380
rect 18782 20312 18788 20324
rect 15580 20284 18788 20312
rect 14148 20272 14154 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19306 20312 19334 20352
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 31588 20380 31616 20411
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 32766 20408 32772 20460
rect 32824 20408 32830 20460
rect 33042 20408 33048 20460
rect 33100 20408 33106 20460
rect 31938 20380 31944 20392
rect 31588 20352 31944 20380
rect 31938 20340 31944 20352
rect 31996 20340 32002 20392
rect 18892 20284 19334 20312
rect 2958 20204 2964 20256
rect 3016 20204 3022 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7834 20244 7840 20256
rect 6972 20216 7840 20244
rect 6972 20204 6978 20216
rect 7834 20204 7840 20216
rect 7892 20244 7898 20256
rect 13081 20247 13139 20253
rect 13081 20244 13093 20247
rect 7892 20216 13093 20244
rect 7892 20204 7898 20216
rect 13081 20213 13093 20216
rect 13127 20213 13139 20247
rect 13081 20207 13139 20213
rect 15841 20247 15899 20253
rect 15841 20213 15853 20247
rect 15887 20244 15899 20247
rect 16850 20244 16856 20256
rect 15887 20216 16856 20244
rect 15887 20213 15899 20216
rect 15841 20207 15899 20213
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 18892 20244 18920 20284
rect 20806 20272 20812 20324
rect 20864 20312 20870 20324
rect 20864 20284 21312 20312
rect 20864 20272 20870 20284
rect 18288 20216 18920 20244
rect 19153 20247 19211 20253
rect 18288 20204 18294 20216
rect 19153 20213 19165 20247
rect 19199 20244 19211 20247
rect 19702 20244 19708 20256
rect 19199 20216 19708 20244
rect 19199 20213 19211 20216
rect 19153 20207 19211 20213
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 21284 20244 21312 20284
rect 27614 20272 27620 20324
rect 27672 20272 27678 20324
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32950 20312 32956 20324
rect 32364 20284 32956 20312
rect 32364 20272 32370 20284
rect 32950 20272 32956 20284
rect 33008 20272 33014 20324
rect 24489 20247 24547 20253
rect 24489 20244 24501 20247
rect 21284 20216 24501 20244
rect 24489 20213 24501 20216
rect 24535 20213 24547 20247
rect 24489 20207 24547 20213
rect 27985 20247 28043 20253
rect 27985 20213 27997 20247
rect 28031 20244 28043 20247
rect 28258 20244 28264 20256
rect 28031 20216 28264 20244
rect 28031 20213 28043 20216
rect 27985 20207 28043 20213
rect 28258 20204 28264 20216
rect 28316 20204 28322 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 3970 20000 3976 20052
rect 4028 20000 4034 20052
rect 7561 20043 7619 20049
rect 4172 20012 5396 20040
rect 2406 19904 2412 19916
rect 1688 19876 2412 19904
rect 1688 19845 1716 19876
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 3234 19864 3240 19916
rect 3292 19904 3298 19916
rect 4172 19904 4200 20012
rect 5077 19975 5135 19981
rect 5077 19941 5089 19975
rect 5123 19941 5135 19975
rect 5077 19935 5135 19941
rect 5368 19972 5396 20012
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7650 20040 7656 20052
rect 7607 20012 7656 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 6914 19972 6920 19984
rect 5368 19944 6920 19972
rect 3292 19876 4200 19904
rect 3292 19864 3298 19876
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 1854 19796 1860 19848
rect 1912 19796 1918 19848
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3510 19836 3516 19848
rect 3191 19808 3516 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3510 19796 3516 19808
rect 3568 19836 3574 19848
rect 4172 19845 4200 19876
rect 4157 19839 4215 19845
rect 3568 19808 4108 19836
rect 3568 19796 3574 19808
rect 1765 19771 1823 19777
rect 1765 19737 1777 19771
rect 1811 19768 1823 19771
rect 3326 19768 3332 19780
rect 1811 19740 3332 19768
rect 1811 19737 1823 19740
rect 1765 19731 1823 19737
rect 3326 19728 3332 19740
rect 3384 19728 3390 19780
rect 4080 19700 4108 19808
rect 4157 19805 4169 19839
rect 4203 19805 4215 19839
rect 4157 19799 4215 19805
rect 4522 19796 4528 19848
rect 4580 19796 4586 19848
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 5092 19836 5120 19935
rect 5368 19845 5396 19944
rect 6914 19932 6920 19944
rect 6972 19932 6978 19984
rect 7098 19932 7104 19984
rect 7156 19932 7162 19984
rect 7576 19904 7604 20003
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20040 14519 20043
rect 15654 20040 15660 20052
rect 14507 20012 15660 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 19242 20040 19248 20052
rect 18831 20012 19248 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 19794 20040 19800 20052
rect 19720 20012 19800 20040
rect 7742 19932 7748 19984
rect 7800 19932 7806 19984
rect 9125 19975 9183 19981
rect 9125 19941 9137 19975
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 9140 19904 9168 19935
rect 9214 19932 9220 19984
rect 9272 19972 9278 19984
rect 9272 19944 14412 19972
rect 9272 19932 9278 19944
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 6932 19876 7604 19904
rect 8312 19876 9168 19904
rect 9416 19876 10517 19904
rect 6932 19845 6960 19876
rect 4663 19808 5120 19836
rect 5353 19839 5411 19845
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 4246 19728 4252 19780
rect 4304 19728 4310 19780
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 4890 19768 4896 19780
rect 4387 19740 4896 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 4890 19728 4896 19740
rect 4948 19728 4954 19780
rect 5074 19728 5080 19780
rect 5132 19728 5138 19780
rect 6840 19768 6868 19799
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 8312 19836 8340 19876
rect 8076 19808 8340 19836
rect 8076 19796 8082 19808
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 9416 19845 9444 19876
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 11882 19904 11888 19916
rect 10505 19867 10563 19873
rect 10796 19876 11888 19904
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8444 19808 9413 19836
rect 8444 19796 8450 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 10410 19796 10416 19848
rect 10468 19796 10474 19848
rect 10796 19845 10824 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 14090 19904 14096 19916
rect 13771 19876 14096 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11103 19808 11713 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 7282 19768 7288 19780
rect 6840 19740 7288 19768
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 9030 19728 9036 19780
rect 9088 19768 9094 19780
rect 9125 19771 9183 19777
rect 9125 19768 9137 19771
rect 9088 19740 9137 19768
rect 9088 19728 9094 19740
rect 9125 19737 9137 19740
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9766 19768 9772 19780
rect 9355 19740 9772 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9766 19728 9772 19740
rect 9824 19768 9830 19780
rect 10226 19768 10232 19780
rect 9824 19740 10232 19768
rect 9824 19728 9830 19740
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 11072 19768 11100 19799
rect 13354 19796 13360 19848
rect 13412 19796 13418 19848
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 14384 19845 14412 19944
rect 19610 19904 19616 19916
rect 15120 19876 19616 19904
rect 15120 19848 15148 19876
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13504 19808 13553 19836
rect 13504 19796 13510 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 15102 19796 15108 19848
rect 15160 19796 15166 19848
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 18509 19839 18567 19845
rect 18509 19836 18521 19839
rect 16908 19808 18521 19836
rect 16908 19796 16914 19808
rect 18509 19805 18521 19808
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19518 19796 19524 19848
rect 19576 19796 19582 19848
rect 19720 19845 19748 20012
rect 19794 20000 19800 20012
rect 19852 20040 19858 20052
rect 20073 20043 20131 20049
rect 19852 20012 20024 20040
rect 19852 20000 19858 20012
rect 19886 19972 19892 19984
rect 19812 19944 19892 19972
rect 19812 19845 19840 19944
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 19996 19972 20024 20012
rect 20073 20009 20085 20043
rect 20119 20040 20131 20043
rect 24762 20040 24768 20052
rect 20119 20012 24768 20040
rect 20119 20009 20131 20012
rect 20073 20003 20131 20009
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 20622 19972 20628 19984
rect 19996 19944 20628 19972
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 32306 19932 32312 19984
rect 32364 19932 32370 19984
rect 21266 19904 21272 19916
rect 20640 19876 21272 19904
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 19886 19796 19892 19848
rect 19944 19845 19950 19848
rect 19944 19836 19952 19845
rect 20640 19836 20668 19876
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 23198 19904 23204 19916
rect 22603 19876 23204 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 32122 19864 32128 19916
rect 32180 19904 32186 19916
rect 32180 19876 32444 19904
rect 32180 19864 32186 19876
rect 32416 19848 32444 19876
rect 19944 19808 20668 19836
rect 19944 19799 19952 19808
rect 19944 19796 19950 19799
rect 31938 19796 31944 19848
rect 31996 19796 32002 19848
rect 32214 19796 32220 19848
rect 32272 19796 32278 19848
rect 32398 19796 32404 19848
rect 32456 19796 32462 19848
rect 32490 19796 32496 19848
rect 32548 19836 32554 19848
rect 32585 19839 32643 19845
rect 32585 19836 32597 19839
rect 32548 19808 32597 19836
rect 32548 19796 32554 19808
rect 32585 19805 32597 19808
rect 32631 19805 32643 19839
rect 32585 19799 32643 19805
rect 10744 19740 11100 19768
rect 10744 19728 10750 19740
rect 15654 19728 15660 19780
rect 15712 19728 15718 19780
rect 16022 19728 16028 19780
rect 16080 19768 16086 19780
rect 16301 19771 16359 19777
rect 16301 19768 16313 19771
rect 16080 19740 16313 19768
rect 16080 19728 16086 19740
rect 16301 19737 16313 19740
rect 16347 19768 16359 19771
rect 16347 19740 19748 19768
rect 16347 19737 16359 19740
rect 16301 19731 16359 19737
rect 4706 19700 4712 19712
rect 4080 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19700 4770 19712
rect 4982 19700 4988 19712
rect 4764 19672 4988 19700
rect 4764 19660 4770 19672
rect 4982 19660 4988 19672
rect 5040 19700 5046 19712
rect 5261 19703 5319 19709
rect 5261 19700 5273 19703
rect 5040 19672 5273 19700
rect 5040 19660 5046 19672
rect 5261 19669 5273 19672
rect 5307 19669 5319 19703
rect 5261 19663 5319 19669
rect 11514 19660 11520 19712
rect 11572 19660 11578 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19610 19700 19616 19712
rect 19484 19672 19616 19700
rect 19484 19660 19490 19672
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 19720 19700 19748 19740
rect 20806 19728 20812 19780
rect 20864 19728 20870 19780
rect 24670 19700 24676 19712
rect 19720 19672 24676 19700
rect 24670 19660 24676 19672
rect 24728 19660 24734 19712
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 1854 19456 1860 19508
rect 1912 19496 1918 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 1912 19468 4445 19496
rect 1912 19456 1918 19468
rect 4433 19465 4445 19468
rect 4479 19496 4491 19499
rect 5074 19496 5080 19508
rect 4479 19468 5080 19496
rect 4479 19465 4491 19468
rect 4433 19459 4491 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 17221 19499 17279 19505
rect 17221 19496 17233 19499
rect 16347 19468 17233 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 17221 19465 17233 19468
rect 17267 19496 17279 19499
rect 19518 19496 19524 19508
rect 17267 19468 19524 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 20349 19499 20407 19505
rect 20349 19465 20361 19499
rect 20395 19496 20407 19499
rect 20990 19496 20996 19508
rect 20395 19468 20996 19496
rect 20395 19465 20407 19468
rect 20349 19459 20407 19465
rect 20990 19456 20996 19468
rect 21048 19496 21054 19508
rect 21177 19499 21235 19505
rect 21177 19496 21189 19499
rect 21048 19468 21189 19496
rect 21048 19456 21054 19468
rect 21177 19465 21189 19468
rect 21223 19465 21235 19499
rect 29178 19496 29184 19508
rect 21177 19459 21235 19465
rect 24964 19468 29184 19496
rect 24964 19440 24992 19468
rect 29178 19456 29184 19468
rect 29236 19456 29242 19508
rect 32490 19456 32496 19508
rect 32548 19496 32554 19508
rect 32585 19499 32643 19505
rect 32585 19496 32597 19499
rect 32548 19468 32597 19496
rect 32548 19456 32554 19468
rect 32585 19465 32597 19468
rect 32631 19465 32643 19499
rect 32585 19459 32643 19465
rect 32861 19499 32919 19505
rect 32861 19465 32873 19499
rect 32907 19496 32919 19499
rect 33042 19496 33048 19508
rect 32907 19468 33048 19496
rect 32907 19465 32919 19468
rect 32861 19459 32919 19465
rect 33042 19456 33048 19468
rect 33100 19456 33106 19508
rect 2768 19431 2826 19437
rect 2768 19397 2780 19431
rect 2814 19428 2826 19431
rect 2958 19428 2964 19440
rect 2814 19400 2964 19428
rect 2814 19397 2826 19400
rect 2768 19391 2826 19397
rect 2958 19388 2964 19400
rect 3016 19388 3022 19440
rect 4540 19400 6776 19428
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 3510 19360 3516 19372
rect 2547 19332 3516 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 3510 19320 3516 19332
rect 3568 19360 3574 19372
rect 4540 19360 4568 19400
rect 6748 19372 6776 19400
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 15838 19428 15844 19440
rect 12492 19400 15844 19428
rect 12492 19388 12498 19400
rect 15838 19388 15844 19400
rect 15896 19388 15902 19440
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 19426 19428 19432 19440
rect 16080 19400 17080 19428
rect 16080 19388 16086 19400
rect 3568 19332 4568 19360
rect 3568 19320 3574 19332
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 6638 19360 6644 19372
rect 4672 19332 6644 19360
rect 4672 19320 4678 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 7101 19363 7159 19369
rect 7101 19360 7113 19363
rect 6788 19332 7113 19360
rect 6788 19320 6794 19332
rect 7101 19329 7113 19332
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7368 19363 7426 19369
rect 7368 19329 7380 19363
rect 7414 19360 7426 19363
rect 7650 19360 7656 19372
rect 7414 19332 7656 19360
rect 7414 19329 7426 19332
rect 7368 19323 7426 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9766 19360 9772 19372
rect 9263 19332 9772 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10376 19332 10701 19360
rect 10376 19320 10382 19332
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10689 19323 10747 19329
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 17052 19369 17080 19400
rect 18984 19400 19432 19428
rect 15188 19363 15246 19369
rect 15188 19329 15200 19363
rect 15234 19360 15246 19363
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15234 19332 16865 19360
rect 15234 19329 15246 19332
rect 15188 19323 15246 19329
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17678 19360 17684 19372
rect 17359 19332 17684 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 18984 19369 19012 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 24765 19431 24823 19437
rect 20128 19400 21312 19428
rect 20128 19388 20134 19400
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19236 19363 19294 19369
rect 19236 19329 19248 19363
rect 19282 19360 19294 19363
rect 20993 19363 21051 19369
rect 19282 19332 20024 19360
rect 19282 19329 19294 19332
rect 19236 19323 19294 19329
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19292 4859 19295
rect 7006 19292 7012 19304
rect 4847 19264 7012 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 3881 19227 3939 19233
rect 3881 19193 3893 19227
rect 3927 19224 3939 19227
rect 4246 19224 4252 19236
rect 3927 19196 4252 19224
rect 3927 19193 3939 19196
rect 3881 19187 3939 19193
rect 4246 19184 4252 19196
rect 4304 19224 4310 19236
rect 4816 19224 4844 19255
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 11054 19292 11060 19304
rect 10459 19264 11060 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 11514 19292 11520 19304
rect 11112 19264 11520 19292
rect 11112 19252 11118 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14792 19264 14933 19292
rect 14792 19252 14798 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 19996 19292 20024 19332
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21082 19360 21088 19372
rect 21039 19332 21088 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21174 19320 21180 19372
rect 21232 19360 21238 19372
rect 21284 19369 21312 19400
rect 24765 19397 24777 19431
rect 24811 19428 24823 19431
rect 24946 19428 24952 19440
rect 24811 19400 24952 19428
rect 24811 19397 24823 19400
rect 24765 19391 24823 19397
rect 24946 19388 24952 19400
rect 25004 19388 25010 19440
rect 28166 19388 28172 19440
rect 28224 19428 28230 19440
rect 28353 19431 28411 19437
rect 28353 19428 28365 19431
rect 28224 19400 28365 19428
rect 28224 19388 28230 19400
rect 28353 19397 28365 19400
rect 28399 19397 28411 19431
rect 29196 19428 29224 19456
rect 29196 19400 31754 19428
rect 28353 19391 28411 19397
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21232 19332 21281 19360
rect 21232 19320 21238 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23198 19360 23204 19372
rect 23155 19332 23204 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 27154 19320 27160 19372
rect 27212 19320 27218 19372
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 27890 19360 27896 19372
rect 27387 19332 27896 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 28994 19320 29000 19372
rect 29052 19320 29058 19372
rect 29362 19320 29368 19372
rect 29420 19320 29426 19372
rect 31220 19369 31248 19400
rect 31205 19363 31263 19369
rect 31205 19329 31217 19363
rect 31251 19329 31263 19363
rect 31205 19323 31263 19329
rect 31294 19320 31300 19372
rect 31352 19360 31358 19372
rect 31389 19363 31447 19369
rect 31389 19360 31401 19363
rect 31352 19332 31401 19360
rect 31352 19320 31358 19332
rect 31389 19329 31401 19332
rect 31435 19329 31447 19363
rect 31726 19360 31754 19400
rect 32214 19388 32220 19440
rect 32272 19428 32278 19440
rect 32677 19431 32735 19437
rect 32677 19428 32689 19431
rect 32272 19400 32689 19428
rect 32272 19388 32278 19400
rect 32677 19397 32689 19400
rect 32723 19397 32735 19431
rect 32677 19391 32735 19397
rect 31938 19360 31944 19372
rect 31726 19332 31944 19360
rect 31389 19323 31447 19329
rect 31938 19320 31944 19332
rect 31996 19360 32002 19372
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 31996 19332 32321 19360
rect 31996 19320 32002 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 32493 19363 32551 19369
rect 32493 19360 32505 19363
rect 32456 19332 32505 19360
rect 32456 19320 32462 19332
rect 32493 19329 32505 19332
rect 32539 19329 32551 19363
rect 32493 19323 32551 19329
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 19996 19264 20821 19292
rect 14921 19255 14979 19261
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 23382 19252 23388 19304
rect 23440 19252 23446 19304
rect 28534 19252 28540 19304
rect 28592 19292 28598 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28592 19264 28825 19292
rect 28592 19252 28598 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 29270 19252 29276 19304
rect 29328 19292 29334 19304
rect 29328 19264 31432 19292
rect 29328 19252 29334 19264
rect 31404 19236 31432 19264
rect 4304 19196 4844 19224
rect 4304 19184 4310 19196
rect 31386 19184 31392 19236
rect 31444 19184 31450 19236
rect 8481 19159 8539 19165
rect 8481 19125 8493 19159
rect 8527 19156 8539 19159
rect 8570 19156 8576 19168
rect 8527 19128 8576 19156
rect 8527 19125 8539 19128
rect 8481 19119 8539 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9122 19116 9128 19168
rect 9180 19116 9186 19168
rect 10134 19116 10140 19168
rect 10192 19116 10198 19168
rect 10594 19116 10600 19168
rect 10652 19116 10658 19168
rect 14918 19116 14924 19168
rect 14976 19156 14982 19168
rect 19334 19156 19340 19168
rect 14976 19128 19340 19156
rect 14976 19116 14982 19128
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 7650 18912 7656 18964
rect 7708 18912 7714 18964
rect 14553 18955 14611 18961
rect 14553 18921 14565 18955
rect 14599 18952 14611 18955
rect 14918 18952 14924 18964
rect 14599 18924 14924 18952
rect 14599 18921 14611 18924
rect 14553 18915 14611 18921
rect 14918 18912 14924 18924
rect 14976 18912 14982 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16264 18924 16681 18952
rect 16264 18912 16270 18924
rect 16669 18921 16681 18924
rect 16715 18952 16727 18955
rect 18230 18952 18236 18964
rect 16715 18924 18236 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18693 18955 18751 18961
rect 18693 18921 18705 18955
rect 18739 18952 18751 18955
rect 19334 18952 19340 18964
rect 18739 18924 19340 18952
rect 18739 18921 18751 18924
rect 18693 18915 18751 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 19794 18952 19800 18964
rect 19444 18924 19800 18952
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3145 18887 3203 18893
rect 3145 18884 3157 18887
rect 3016 18856 3157 18884
rect 3016 18844 3022 18856
rect 3145 18853 3157 18856
rect 3191 18853 3203 18887
rect 8386 18884 8392 18896
rect 3145 18847 3203 18853
rect 7944 18856 8392 18884
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7944 18825 7972 18856
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 19444 18884 19472 18924
rect 19794 18912 19800 18924
rect 19852 18912 19858 18964
rect 20809 18955 20867 18961
rect 20809 18921 20821 18955
rect 20855 18952 20867 18955
rect 20898 18952 20904 18964
rect 20855 18924 20904 18952
rect 20855 18921 20867 18924
rect 20809 18915 20867 18921
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 25866 18912 25872 18964
rect 25924 18912 25930 18964
rect 33137 18955 33195 18961
rect 33137 18921 33149 18955
rect 33183 18952 33195 18955
rect 33318 18952 33324 18964
rect 33183 18924 33324 18952
rect 33183 18921 33195 18924
rect 33137 18915 33195 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 27706 18884 27712 18896
rect 19352 18856 19472 18884
rect 26068 18856 27712 18884
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7156 18788 7849 18816
rect 7156 18776 7162 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 9122 18816 9128 18828
rect 8251 18788 9128 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18816 12403 18819
rect 12391 18788 15424 18816
rect 12391 18785 12403 18788
rect 12345 18779 12403 18785
rect 15396 18760 15424 18788
rect 3326 18708 3332 18760
rect 3384 18708 3390 18760
rect 3418 18708 3424 18760
rect 3476 18708 3482 18760
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 10134 18748 10140 18760
rect 8343 18720 10140 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10594 18748 10600 18760
rect 10551 18720 10600 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3234 18680 3240 18692
rect 3191 18652 3240 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3234 18640 3240 18652
rect 3292 18680 3298 18692
rect 7190 18680 7196 18692
rect 3292 18652 7196 18680
rect 3292 18640 3298 18652
rect 7190 18640 7196 18652
rect 7248 18680 7254 18692
rect 7248 18652 8064 18680
rect 7248 18640 7254 18652
rect 8036 18621 8064 18652
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 10428 18680 10456 18711
rect 10594 18708 10600 18720
rect 10652 18748 10658 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 10652 18720 11989 18748
rect 10652 18708 10658 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12434 18748 12440 18760
rect 12299 18720 12440 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14792 18720 15301 18748
rect 14792 18708 14798 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15378 18708 15384 18760
rect 15436 18708 15442 18760
rect 16942 18748 16948 18760
rect 15488 18720 16948 18748
rect 9824 18652 10456 18680
rect 9824 18640 9830 18652
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 12124 18652 14381 18680
rect 12124 18640 12130 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14553 18683 14611 18689
rect 14553 18649 14565 18683
rect 14599 18680 14611 18683
rect 15488 18680 15516 18720
rect 16942 18708 16948 18720
rect 17000 18748 17006 18760
rect 19352 18748 19380 18856
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 21876 18788 24808 18816
rect 21876 18776 21882 18788
rect 17000 18720 19380 18748
rect 17000 18708 17006 18720
rect 19426 18708 19432 18760
rect 19484 18708 19490 18760
rect 20714 18748 20720 18760
rect 19628 18720 20720 18748
rect 14599 18652 15516 18680
rect 15556 18683 15614 18689
rect 14599 18649 14611 18652
rect 14553 18643 14611 18649
rect 15556 18649 15568 18683
rect 15602 18680 15614 18683
rect 15746 18680 15752 18692
rect 15602 18652 15752 18680
rect 15602 18649 15614 18652
rect 15556 18643 15614 18649
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 18877 18683 18935 18689
rect 18877 18649 18889 18683
rect 18923 18680 18935 18683
rect 19518 18680 19524 18692
rect 18923 18652 19524 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 19518 18640 19524 18652
rect 19576 18680 19582 18692
rect 19628 18680 19656 18720
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 23750 18708 23756 18760
rect 23808 18708 23814 18760
rect 24780 18757 24808 18788
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18717 24087 18751
rect 24029 18711 24087 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 25130 18748 25136 18760
rect 25087 18720 25136 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 19702 18689 19708 18692
rect 19576 18652 19656 18680
rect 19576 18640 19582 18652
rect 19696 18643 19708 18689
rect 19760 18680 19766 18692
rect 24044 18680 24072 18711
rect 25056 18680 25084 18711
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 26068 18757 26096 18856
rect 27706 18844 27712 18856
rect 27764 18844 27770 18896
rect 26145 18819 26203 18825
rect 26145 18785 26157 18819
rect 26191 18816 26203 18819
rect 27246 18816 27252 18828
rect 26191 18788 27252 18816
rect 26191 18785 26203 18788
rect 26145 18779 26203 18785
rect 27246 18776 27252 18788
rect 27304 18776 27310 18828
rect 29086 18776 29092 18828
rect 29144 18816 29150 18828
rect 31849 18819 31907 18825
rect 29144 18788 30052 18816
rect 29144 18776 29150 18788
rect 26053 18751 26111 18757
rect 26053 18717 26065 18751
rect 26099 18717 26111 18751
rect 26053 18711 26111 18717
rect 26234 18708 26240 18760
rect 26292 18708 26298 18760
rect 26329 18751 26387 18757
rect 26329 18717 26341 18751
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 19760 18652 19796 18680
rect 24044 18652 25084 18680
rect 19702 18640 19708 18643
rect 19760 18640 19766 18652
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 14737 18615 14795 18621
rect 14737 18581 14749 18615
rect 14783 18612 14795 18615
rect 15194 18612 15200 18624
rect 14783 18584 15200 18612
rect 14783 18581 14795 18584
rect 14737 18575 14795 18581
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 18506 18572 18512 18624
rect 18564 18572 18570 18624
rect 18690 18572 18696 18624
rect 18748 18612 18754 18624
rect 19886 18612 19892 18624
rect 18748 18584 19892 18612
rect 18748 18572 18754 18584
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 23566 18572 23572 18624
rect 23624 18572 23630 18624
rect 23937 18615 23995 18621
rect 23937 18581 23949 18615
rect 23983 18612 23995 18615
rect 24486 18612 24492 18624
rect 23983 18584 24492 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 25056 18612 25084 18652
rect 25682 18640 25688 18692
rect 25740 18680 25746 18692
rect 26344 18680 26372 18711
rect 27154 18708 27160 18760
rect 27212 18748 27218 18760
rect 27522 18748 27528 18760
rect 27212 18720 27528 18748
rect 27212 18708 27218 18720
rect 27522 18708 27528 18720
rect 27580 18748 27586 18760
rect 27709 18751 27767 18757
rect 27709 18748 27721 18751
rect 27580 18720 27721 18748
rect 27580 18708 27586 18720
rect 27709 18717 27721 18720
rect 27755 18717 27767 18751
rect 27709 18711 27767 18717
rect 27890 18708 27896 18760
rect 27948 18708 27954 18760
rect 28534 18708 28540 18760
rect 28592 18708 28598 18760
rect 28626 18708 28632 18760
rect 28684 18748 28690 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28684 18720 28825 18748
rect 28684 18708 28690 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29270 18748 29276 18760
rect 29043 18720 29276 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 25740 18652 26372 18680
rect 25740 18640 25746 18652
rect 27338 18640 27344 18692
rect 27396 18640 27402 18692
rect 28828 18680 28856 18711
rect 29270 18708 29276 18720
rect 29328 18708 29334 18760
rect 29822 18708 29828 18760
rect 29880 18708 29886 18760
rect 30024 18757 30052 18788
rect 31849 18785 31861 18819
rect 31895 18816 31907 18819
rect 32490 18816 32496 18828
rect 31895 18788 32496 18816
rect 31895 18785 31907 18788
rect 31849 18779 31907 18785
rect 32490 18776 32496 18788
rect 32548 18776 32554 18828
rect 32582 18776 32588 18828
rect 32640 18816 32646 18828
rect 32769 18819 32827 18825
rect 32769 18816 32781 18819
rect 32640 18788 32781 18816
rect 32640 18776 32646 18788
rect 32769 18785 32781 18788
rect 32815 18785 32827 18819
rect 32769 18779 32827 18785
rect 30009 18751 30067 18757
rect 30009 18717 30021 18751
rect 30055 18717 30067 18751
rect 30009 18711 30067 18717
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 32217 18751 32275 18757
rect 32217 18717 32229 18751
rect 32263 18748 32275 18751
rect 32677 18751 32735 18757
rect 32677 18748 32689 18751
rect 32263 18720 32689 18748
rect 32263 18717 32275 18720
rect 32217 18711 32275 18717
rect 32677 18717 32689 18720
rect 32723 18717 32735 18751
rect 32677 18711 32735 18717
rect 29362 18680 29368 18692
rect 28828 18652 29368 18680
rect 29362 18640 29368 18652
rect 29420 18680 29426 18692
rect 29733 18683 29791 18689
rect 29733 18680 29745 18683
rect 29420 18652 29745 18680
rect 29420 18640 29426 18652
rect 29733 18649 29745 18652
rect 29779 18649 29791 18683
rect 32048 18680 32076 18711
rect 32858 18708 32864 18760
rect 32916 18748 32922 18760
rect 32953 18751 33011 18757
rect 32953 18748 32965 18751
rect 32916 18720 32965 18748
rect 32916 18708 32922 18720
rect 32953 18717 32965 18720
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 32398 18680 32404 18692
rect 32048 18652 32404 18680
rect 29733 18643 29791 18649
rect 32398 18640 32404 18652
rect 32456 18640 32462 18692
rect 26142 18612 26148 18624
rect 25056 18584 26148 18612
rect 26142 18572 26148 18584
rect 26200 18572 26206 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 27356 18612 27384 18640
rect 26292 18584 27384 18612
rect 26292 18572 26298 18584
rect 28350 18572 28356 18624
rect 28408 18572 28414 18624
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 9030 18408 9036 18420
rect 8251 18380 9036 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 15746 18368 15752 18420
rect 15804 18368 15810 18420
rect 16117 18411 16175 18417
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16206 18408 16212 18420
rect 16163 18380 16212 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 19426 18368 19432 18420
rect 19484 18408 19490 18420
rect 19794 18408 19800 18420
rect 19484 18380 19800 18408
rect 19484 18368 19490 18380
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 25682 18368 25688 18420
rect 25740 18368 25746 18420
rect 32769 18411 32827 18417
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 32858 18408 32864 18420
rect 32815 18380 32864 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 32858 18368 32864 18380
rect 32916 18368 32922 18420
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 6825 18343 6883 18349
rect 6825 18340 6837 18343
rect 6512 18312 6837 18340
rect 6512 18300 6518 18312
rect 6825 18309 6837 18312
rect 6871 18309 6883 18343
rect 6825 18303 6883 18309
rect 12066 18300 12072 18352
rect 12124 18340 12130 18352
rect 12124 18312 12480 18340
rect 12124 18300 12130 18312
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 6696 18244 8033 18272
rect 6696 18232 6702 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8021 18235 8079 18241
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8570 18272 8576 18284
rect 8251 18244 8576 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8570 18232 8576 18244
rect 8628 18272 8634 18284
rect 9766 18272 9772 18284
rect 8628 18244 9772 18272
rect 8628 18232 8634 18244
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 11054 18272 11060 18284
rect 10367 18244 11060 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11848 18244 12265 18272
rect 11848 18232 11854 18244
rect 12253 18241 12265 18244
rect 12299 18272 12311 18275
rect 12342 18272 12348 18284
rect 12299 18244 12348 18272
rect 12299 18241 12311 18244
rect 12253 18235 12311 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12452 18281 12480 18312
rect 14734 18300 14740 18352
rect 14792 18300 14798 18352
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 15896 18312 16252 18340
rect 15896 18300 15902 18312
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 16224 18281 16252 18312
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 19245 18343 19303 18349
rect 19245 18340 19257 18343
rect 18564 18312 19257 18340
rect 18564 18300 18570 18312
rect 19245 18309 19257 18312
rect 19291 18309 19303 18343
rect 19245 18303 19303 18309
rect 24857 18343 24915 18349
rect 24857 18309 24869 18343
rect 24903 18340 24915 18343
rect 24946 18340 24952 18352
rect 24903 18312 24952 18340
rect 24903 18309 24915 18312
rect 24857 18303 24915 18309
rect 24946 18300 24952 18312
rect 25004 18340 25010 18352
rect 28442 18340 28448 18352
rect 25004 18312 28448 18340
rect 25004 18300 25010 18312
rect 28442 18300 28448 18312
rect 28500 18300 28506 18352
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15712 18244 15945 18272
rect 15712 18232 15718 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 16209 18275 16267 18281
rect 16209 18241 16221 18275
rect 16255 18241 16267 18275
rect 16209 18235 16267 18241
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18272 23535 18275
rect 24578 18272 24584 18284
rect 23523 18244 24584 18272
rect 23523 18241 23535 18244
rect 23477 18235 23535 18241
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 6914 18164 6920 18216
rect 6972 18164 6978 18216
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 15948 18204 15976 18235
rect 24578 18232 24584 18244
rect 24636 18232 24642 18284
rect 25314 18232 25320 18284
rect 25372 18232 25378 18284
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18272 27951 18275
rect 28350 18272 28356 18284
rect 27939 18244 28356 18272
rect 27939 18241 27951 18244
rect 27893 18235 27951 18241
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28718 18232 28724 18284
rect 28776 18232 28782 18284
rect 29086 18232 29092 18284
rect 29144 18232 29150 18284
rect 29178 18232 29184 18284
rect 29236 18272 29242 18284
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 29236 18244 29377 18272
rect 29236 18232 29242 18244
rect 29365 18241 29377 18244
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 29730 18232 29736 18284
rect 29788 18232 29794 18284
rect 32490 18232 32496 18284
rect 32548 18232 32554 18284
rect 17126 18204 17132 18216
rect 15948 18176 17132 18204
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 23106 18164 23112 18216
rect 23164 18204 23170 18216
rect 23201 18207 23259 18213
rect 23201 18204 23213 18207
rect 23164 18176 23213 18204
rect 23164 18164 23170 18176
rect 23201 18173 23213 18176
rect 23247 18173 23259 18207
rect 23201 18167 23259 18173
rect 25406 18164 25412 18216
rect 25464 18164 25470 18216
rect 27522 18164 27528 18216
rect 27580 18164 27586 18216
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18204 28043 18207
rect 28994 18204 29000 18216
rect 28031 18176 29000 18204
rect 28031 18173 28043 18176
rect 27985 18167 28043 18173
rect 28994 18164 29000 18176
rect 29052 18164 29058 18216
rect 32306 18164 32312 18216
rect 32364 18164 32370 18216
rect 32858 18164 32864 18216
rect 32916 18164 32922 18216
rect 34333 18207 34391 18213
rect 34333 18173 34345 18207
rect 34379 18204 34391 18207
rect 35066 18204 35072 18216
rect 34379 18176 35072 18204
rect 34379 18173 34391 18176
rect 34333 18167 34391 18173
rect 35066 18164 35072 18176
rect 35124 18164 35130 18216
rect 7282 18096 7288 18148
rect 7340 18096 7346 18148
rect 28534 18096 28540 18148
rect 28592 18136 28598 18148
rect 28629 18139 28687 18145
rect 28629 18136 28641 18139
rect 28592 18108 28641 18136
rect 28592 18096 28598 18108
rect 28629 18105 28641 18108
rect 28675 18105 28687 18139
rect 28629 18099 28687 18105
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 18230 18028 18236 18080
rect 18288 18068 18294 18080
rect 20533 18071 20591 18077
rect 20533 18068 20545 18071
rect 18288 18040 20545 18068
rect 18288 18028 18294 18040
rect 20533 18037 20545 18040
rect 20579 18037 20591 18071
rect 20533 18031 20591 18037
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 25280 18040 25329 18068
rect 25280 18028 25286 18040
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 25317 18031 25375 18037
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 6730 17864 6736 17876
rect 6503 17836 6736 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 21637 17867 21695 17873
rect 15436 17836 21404 17864
rect 15436 17824 15442 17836
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 3510 17796 3516 17808
rect 3467 17768 3516 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 11664 17700 13093 17728
rect 11664 17688 11670 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 18708 17700 19564 17728
rect 3234 17620 3240 17672
rect 3292 17620 3298 17672
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 6549 17663 6607 17669
rect 6549 17629 6561 17663
rect 6595 17660 6607 17663
rect 7098 17660 7104 17672
rect 6595 17632 7104 17660
rect 6595 17629 6607 17632
rect 6549 17623 6607 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 15194 17620 15200 17672
rect 15252 17620 15258 17672
rect 17402 17620 17408 17672
rect 17460 17660 17466 17672
rect 18708 17669 18736 17700
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 17460 17632 17601 17660
rect 17460 17620 17466 17632
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17660 17923 17663
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 17911 17632 18429 17660
rect 17911 17629 17923 17632
rect 17865 17623 17923 17629
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 2869 17595 2927 17601
rect 2869 17592 2881 17595
rect 2740 17564 2881 17592
rect 2740 17552 2746 17564
rect 2869 17561 2881 17564
rect 2915 17561 2927 17595
rect 2869 17555 2927 17561
rect 12158 17552 12164 17604
rect 12216 17552 12222 17604
rect 12802 17552 12808 17604
rect 12860 17552 12866 17604
rect 16206 17552 16212 17604
rect 16264 17592 16270 17604
rect 17880 17592 17908 17623
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19300 17632 19441 17660
rect 19300 17620 19306 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19536 17660 19564 17700
rect 21376 17669 21404 17836
rect 21637 17833 21649 17867
rect 21683 17864 21695 17867
rect 21818 17864 21824 17876
rect 21683 17836 21824 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 21361 17663 21419 17669
rect 19536 17632 21036 17660
rect 19429 17623 19487 17629
rect 16264 17564 17908 17592
rect 18877 17595 18935 17601
rect 16264 17552 16270 17564
rect 18877 17561 18889 17595
rect 18923 17592 18935 17595
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 18923 17564 19686 17592
rect 18923 17561 18935 17564
rect 18877 17555 18935 17561
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 21008 17592 21036 17632
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21652 17592 21680 17827
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 27982 17824 27988 17876
rect 28040 17824 28046 17876
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 32677 17867 32735 17873
rect 32677 17864 32689 17867
rect 29052 17836 32689 17864
rect 29052 17824 29058 17836
rect 32677 17833 32689 17836
rect 32723 17833 32735 17867
rect 32677 17827 32735 17833
rect 23750 17756 23756 17808
rect 23808 17796 23814 17808
rect 32306 17796 32312 17808
rect 23808 17768 30880 17796
rect 23808 17756 23814 17768
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 25774 17728 25780 17740
rect 24728 17700 25780 17728
rect 24728 17688 24734 17700
rect 24780 17669 24808 17700
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 27617 17731 27675 17737
rect 27617 17697 27629 17731
rect 27663 17728 27675 17731
rect 27890 17728 27896 17740
rect 27663 17700 27896 17728
rect 27663 17697 27675 17700
rect 27617 17691 27675 17697
rect 27890 17688 27896 17700
rect 27948 17728 27954 17740
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 27948 17700 28457 17728
rect 27948 17688 27954 17700
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 28445 17691 28503 17697
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17629 24823 17663
rect 24765 17623 24823 17629
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 21008 17564 21680 17592
rect 25056 17592 25084 17623
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 25740 17632 27537 17660
rect 25740 17620 25746 17632
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27525 17623 27583 17629
rect 27706 17620 27712 17672
rect 27764 17620 27770 17672
rect 27798 17620 27804 17672
rect 27856 17620 27862 17672
rect 28534 17620 28540 17672
rect 28592 17660 28598 17672
rect 28629 17663 28687 17669
rect 28629 17660 28641 17663
rect 28592 17632 28641 17660
rect 28592 17620 28598 17632
rect 28629 17629 28641 17632
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 28902 17620 28908 17672
rect 28960 17660 28966 17672
rect 30745 17663 30803 17669
rect 30745 17660 30757 17663
rect 28960 17632 30757 17660
rect 28960 17620 28966 17632
rect 30745 17629 30757 17632
rect 30791 17629 30803 17663
rect 30745 17623 30803 17629
rect 26602 17592 26608 17604
rect 25056 17564 26608 17592
rect 19674 17555 19732 17561
rect 26602 17552 26608 17564
rect 26660 17552 26666 17604
rect 3050 17484 3056 17536
rect 3108 17484 3114 17536
rect 3142 17484 3148 17536
rect 3200 17484 3206 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11333 17527 11391 17533
rect 11333 17524 11345 17527
rect 11020 17496 11345 17524
rect 11020 17484 11026 17496
rect 11333 17493 11345 17496
rect 11379 17493 11391 17527
rect 11333 17487 11391 17493
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 13044 17496 16497 17524
rect 13044 17484 13050 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 16632 17496 17417 17524
rect 16632 17484 16638 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 17405 17487 17463 17493
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17773 17527 17831 17533
rect 17773 17524 17785 17527
rect 17552 17496 17785 17524
rect 17552 17484 17558 17496
rect 17773 17493 17785 17496
rect 17819 17493 17831 17527
rect 17773 17487 17831 17493
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 20809 17527 20867 17533
rect 20809 17524 20821 17527
rect 18555 17496 20821 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 20809 17493 20821 17496
rect 20855 17524 20867 17527
rect 20898 17524 20904 17536
rect 20855 17496 20904 17524
rect 20855 17493 20867 17496
rect 20809 17487 20867 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 24581 17527 24639 17533
rect 24581 17493 24593 17527
rect 24627 17524 24639 17527
rect 24854 17524 24860 17536
rect 24627 17496 24860 17524
rect 24627 17493 24639 17496
rect 24581 17487 24639 17493
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 24949 17527 25007 17533
rect 24949 17493 24961 17527
rect 24995 17524 25007 17527
rect 25958 17524 25964 17536
rect 24995 17496 25964 17524
rect 24995 17493 25007 17496
rect 24949 17487 25007 17493
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 28810 17484 28816 17536
rect 28868 17484 28874 17536
rect 30852 17524 30880 17768
rect 31772 17768 32312 17796
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 31772 17669 31800 17768
rect 32306 17756 32312 17768
rect 32364 17796 32370 17808
rect 32364 17768 33640 17796
rect 32364 17756 32370 17768
rect 33612 17737 33640 17768
rect 33597 17731 33655 17737
rect 31956 17700 33456 17728
rect 31956 17669 31984 17700
rect 33428 17672 33456 17700
rect 33597 17697 33609 17731
rect 33643 17697 33655 17731
rect 33597 17691 33655 17697
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 30984 17632 31769 17660
rect 30984 17620 30990 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 31757 17623 31815 17629
rect 31941 17663 31999 17669
rect 31941 17629 31953 17663
rect 31987 17629 31999 17663
rect 31941 17623 31999 17629
rect 32582 17620 32588 17672
rect 32640 17660 32646 17672
rect 33229 17663 33287 17669
rect 33229 17660 33241 17663
rect 32640 17632 33241 17660
rect 32640 17620 32646 17632
rect 33229 17629 33241 17632
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 33410 17620 33416 17672
rect 33468 17620 33474 17672
rect 31110 17552 31116 17604
rect 31168 17552 31174 17604
rect 31849 17595 31907 17601
rect 31849 17561 31861 17595
rect 31895 17592 31907 17595
rect 32401 17595 32459 17601
rect 32401 17592 32413 17595
rect 31895 17564 32413 17592
rect 31895 17561 31907 17564
rect 31849 17555 31907 17561
rect 32401 17561 32413 17564
rect 32447 17561 32459 17595
rect 32401 17555 32459 17561
rect 31938 17524 31944 17536
rect 30852 17496 31944 17524
rect 31938 17484 31944 17496
rect 31996 17484 32002 17536
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 6914 17320 6920 17332
rect 4479 17292 6920 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 19628 17292 22094 17320
rect 2958 17212 2964 17264
rect 3016 17212 3022 17264
rect 6932 17252 6960 17280
rect 6932 17224 8248 17252
rect 4246 17184 4252 17196
rect 4094 17156 4252 17184
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 6638 17144 6644 17196
rect 6696 17144 6702 17196
rect 6730 17144 6736 17196
rect 6788 17144 6794 17196
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6880 17156 7113 17184
rect 6880 17144 6886 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7524 17156 7573 17184
rect 7524 17144 7530 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8220 17193 8248 17224
rect 9214 17212 9220 17264
rect 9272 17252 9278 17264
rect 9585 17255 9643 17261
rect 9585 17252 9597 17255
rect 9272 17224 9597 17252
rect 9272 17212 9278 17224
rect 9585 17221 9597 17224
rect 9631 17252 9643 17255
rect 10318 17252 10324 17264
rect 9631 17224 10324 17252
rect 9631 17221 9643 17224
rect 9585 17215 9643 17221
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 13170 17212 13176 17264
rect 13228 17252 13234 17264
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 13228 17224 13277 17252
rect 13228 17212 13234 17224
rect 13265 17221 13277 17224
rect 13311 17221 13323 17255
rect 13265 17215 13323 17221
rect 18230 17212 18236 17264
rect 18288 17212 18294 17264
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 15436 17156 16221 17184
rect 15436 17144 15442 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16724 17156 16865 17184
rect 16724 17144 16730 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17218 17184 17224 17196
rect 17175 17156 17224 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17218 17144 17224 17156
rect 17276 17184 17282 17196
rect 19628 17184 19656 17292
rect 19794 17212 19800 17264
rect 19852 17212 19858 17264
rect 20809 17255 20867 17261
rect 20809 17221 20821 17255
rect 20855 17252 20867 17255
rect 21174 17252 21180 17264
rect 20855 17224 21180 17252
rect 20855 17221 20867 17224
rect 20809 17215 20867 17221
rect 21174 17212 21180 17224
rect 21232 17212 21238 17264
rect 17276 17156 19656 17184
rect 20625 17187 20683 17193
rect 17276 17144 17282 17156
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 21082 17184 21088 17196
rect 20947 17156 21088 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 2682 17076 2688 17128
rect 2740 17076 2746 17128
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 7064 17088 9781 17116
rect 7064 17076 7070 17088
rect 9769 17085 9781 17088
rect 9815 17116 9827 17119
rect 10594 17116 10600 17128
rect 9815 17088 10600 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 11664 17088 13553 17116
rect 11664 17076 11670 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 15930 17076 15936 17128
rect 15988 17076 15994 17128
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 20640 17116 20668 17147
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 22066 17184 22094 17292
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 22796 17292 25360 17320
rect 22796 17280 22802 17292
rect 23376 17255 23434 17261
rect 23376 17221 23388 17255
rect 23422 17252 23434 17255
rect 23566 17252 23572 17264
rect 23422 17224 23572 17252
rect 23422 17221 23434 17224
rect 23376 17215 23434 17221
rect 23566 17212 23572 17224
rect 23624 17212 23630 17264
rect 23750 17184 23756 17196
rect 22066 17156 23756 17184
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 25038 17144 25044 17196
rect 25096 17144 25102 17196
rect 25332 17193 25360 17292
rect 25682 17280 25688 17332
rect 25740 17280 25746 17332
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 28537 17323 28595 17329
rect 28537 17320 28549 17323
rect 27856 17292 28549 17320
rect 27856 17280 27862 17292
rect 28537 17289 28549 17292
rect 28583 17289 28595 17323
rect 28537 17283 28595 17289
rect 28810 17280 28816 17332
rect 28868 17280 28874 17332
rect 30006 17280 30012 17332
rect 30064 17320 30070 17332
rect 30745 17323 30803 17329
rect 30745 17320 30757 17323
rect 30064 17292 30757 17320
rect 30064 17280 30070 17292
rect 30745 17289 30757 17292
rect 30791 17289 30803 17323
rect 30745 17283 30803 17289
rect 30926 17280 30932 17332
rect 30984 17280 30990 17332
rect 32214 17320 32220 17332
rect 31496 17292 32220 17320
rect 25409 17255 25467 17261
rect 25409 17221 25421 17255
rect 25455 17252 25467 17255
rect 25958 17252 25964 17264
rect 25455 17224 25964 17252
rect 25455 17221 25467 17224
rect 25409 17215 25467 17221
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 28629 17255 28687 17261
rect 28629 17221 28641 17255
rect 28675 17252 28687 17255
rect 28828 17252 28856 17280
rect 31496 17261 31524 17292
rect 32214 17280 32220 17292
rect 32272 17320 32278 17332
rect 32509 17323 32567 17329
rect 32509 17320 32521 17323
rect 32272 17292 32521 17320
rect 32272 17280 32278 17292
rect 32509 17289 32521 17292
rect 32555 17289 32567 17323
rect 32509 17283 32567 17289
rect 32677 17323 32735 17329
rect 32677 17289 32689 17323
rect 32723 17320 32735 17323
rect 32858 17320 32864 17332
rect 32723 17292 32864 17320
rect 32723 17289 32735 17292
rect 32677 17283 32735 17289
rect 32858 17280 32864 17292
rect 32916 17280 32922 17332
rect 33229 17323 33287 17329
rect 33229 17289 33241 17323
rect 33275 17320 33287 17323
rect 33410 17320 33416 17332
rect 33275 17292 33416 17320
rect 33275 17289 33287 17292
rect 33229 17283 33287 17289
rect 33410 17280 33416 17292
rect 33468 17280 33474 17332
rect 29825 17255 29883 17261
rect 29825 17252 29837 17255
rect 28675 17224 29837 17252
rect 28675 17221 28687 17224
rect 28629 17215 28687 17221
rect 29825 17221 29837 17224
rect 29871 17221 29883 17255
rect 30837 17255 30895 17261
rect 30837 17252 30849 17255
rect 29825 17215 29883 17221
rect 29932 17224 30849 17252
rect 25134 17187 25192 17193
rect 25134 17153 25146 17187
rect 25180 17153 25192 17187
rect 25134 17147 25192 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25506 17187 25564 17193
rect 25506 17184 25518 17187
rect 25317 17147 25375 17153
rect 25424 17156 25518 17184
rect 17460 17088 20668 17116
rect 17460 17076 17466 17088
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23106 17116 23112 17128
rect 22612 17088 23112 17116
rect 22612 17076 22618 17088
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 6454 17008 6460 17060
rect 6512 17048 6518 17060
rect 10410 17048 10416 17060
rect 6512 17020 10416 17048
rect 6512 17008 6518 17020
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 25148 17048 25176 17147
rect 24044 17020 25176 17048
rect 8202 16940 8208 16992
rect 8260 16940 8266 16992
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 10042 16940 10048 16992
rect 10100 16940 10106 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11204 16952 11805 16980
rect 11204 16940 11210 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19518 16980 19524 16992
rect 19392 16952 19524 16980
rect 19392 16940 19398 16952
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 20438 16940 20444 16992
rect 20496 16940 20502 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 24044 16980 24072 17020
rect 22520 16952 24072 16980
rect 22520 16940 22526 16952
rect 24486 16940 24492 16992
rect 24544 16940 24550 16992
rect 24762 16940 24768 16992
rect 24820 16980 24826 16992
rect 25424 16980 25452 17156
rect 25506 17153 25518 17156
rect 25552 17153 25564 17187
rect 25506 17147 25564 17153
rect 26142 17144 26148 17196
rect 26200 17144 26206 17196
rect 28534 17144 28540 17196
rect 28592 17144 28598 17196
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17184 28871 17187
rect 28902 17184 28908 17196
rect 28859 17156 28908 17184
rect 28859 17153 28871 17156
rect 28813 17147 28871 17153
rect 28902 17144 28908 17156
rect 28960 17144 28966 17196
rect 29932 17193 29960 17224
rect 30837 17221 30849 17224
rect 30883 17252 30895 17255
rect 31481 17255 31539 17261
rect 31481 17252 31493 17255
rect 30883 17224 31493 17252
rect 30883 17221 30895 17224
rect 30837 17215 30895 17221
rect 31481 17221 31493 17224
rect 31527 17221 31539 17255
rect 32309 17255 32367 17261
rect 32309 17252 32321 17255
rect 31481 17215 31539 17221
rect 31680 17224 32321 17252
rect 29733 17187 29791 17193
rect 29733 17153 29745 17187
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 30613 17187 30671 17193
rect 30613 17153 30625 17187
rect 30659 17184 30671 17187
rect 31294 17184 31300 17196
rect 30659 17156 31300 17184
rect 30659 17153 30671 17156
rect 30613 17147 30671 17153
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 26602 17116 26608 17128
rect 26467 17088 26608 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 26602 17076 26608 17088
rect 26660 17076 26666 17128
rect 29748 17116 29776 17147
rect 30282 17116 30288 17128
rect 29748 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17116 30346 17128
rect 30484 17116 30512 17147
rect 31294 17144 31300 17156
rect 31352 17144 31358 17196
rect 31386 17144 31392 17196
rect 31444 17184 31450 17196
rect 31680 17193 31708 17224
rect 32309 17221 32321 17224
rect 32355 17221 32367 17255
rect 32309 17215 32367 17221
rect 31665 17187 31723 17193
rect 31665 17184 31677 17187
rect 31444 17156 31677 17184
rect 31444 17144 31450 17156
rect 31665 17153 31677 17156
rect 31711 17153 31723 17187
rect 31665 17147 31723 17153
rect 31757 17187 31815 17193
rect 31757 17153 31769 17187
rect 31803 17184 31815 17187
rect 32582 17184 32588 17196
rect 31803 17156 32588 17184
rect 31803 17153 31815 17156
rect 31757 17147 31815 17153
rect 32582 17144 32588 17156
rect 32640 17144 32646 17196
rect 32876 17184 32904 17280
rect 33137 17187 33195 17193
rect 33137 17184 33149 17187
rect 32876 17156 33149 17184
rect 33137 17153 33149 17156
rect 33183 17153 33195 17187
rect 33137 17147 33195 17153
rect 33321 17187 33379 17193
rect 33321 17153 33333 17187
rect 33367 17153 33379 17187
rect 33321 17147 33379 17153
rect 33336 17116 33364 17147
rect 30340 17088 30512 17116
rect 31726 17088 33364 17116
rect 30340 17076 30346 17088
rect 31481 17051 31539 17057
rect 31481 17017 31493 17051
rect 31527 17048 31539 17051
rect 31726 17048 31754 17088
rect 31527 17020 31754 17048
rect 31527 17017 31539 17020
rect 31481 17011 31539 17017
rect 24820 16952 25452 16980
rect 32493 16983 32551 16989
rect 24820 16940 24826 16952
rect 32493 16949 32505 16983
rect 32539 16980 32551 16983
rect 32582 16980 32588 16992
rect 32539 16952 32588 16980
rect 32539 16949 32551 16952
rect 32493 16943 32551 16949
rect 32582 16940 32588 16952
rect 32640 16940 32646 16992
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 2682 16736 2688 16788
rect 2740 16776 2746 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2740 16748 3065 16776
rect 2740 16736 2746 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 3053 16739 3111 16745
rect 3234 16736 3240 16788
rect 3292 16736 3298 16788
rect 4246 16736 4252 16788
rect 4304 16736 4310 16788
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 6825 16779 6883 16785
rect 6825 16776 6837 16779
rect 6696 16748 6837 16776
rect 6696 16736 6702 16748
rect 6825 16745 6837 16748
rect 6871 16745 6883 16779
rect 6825 16739 6883 16745
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 8260 16748 9781 16776
rect 8260 16736 8266 16748
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 9769 16739 9827 16745
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10962 16776 10968 16788
rect 9916 16748 10968 16776
rect 9916 16736 9922 16748
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 12250 16736 12256 16788
rect 12308 16736 12314 16788
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 21361 16779 21419 16785
rect 21361 16776 21373 16779
rect 21140 16748 21373 16776
rect 21140 16736 21146 16748
rect 21361 16745 21373 16748
rect 21407 16745 21419 16779
rect 21361 16739 21419 16745
rect 25958 16736 25964 16788
rect 26016 16736 26022 16788
rect 31110 16736 31116 16788
rect 31168 16776 31174 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 31168 16748 31217 16776
rect 31168 16736 31174 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 31205 16739 31263 16745
rect 32214 16736 32220 16788
rect 32272 16736 32278 16788
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16677 5963 16711
rect 5905 16671 5963 16677
rect 2590 16600 2596 16652
rect 2648 16640 2654 16652
rect 5920 16640 5948 16671
rect 6454 16668 6460 16720
rect 6512 16708 6518 16720
rect 7193 16711 7251 16717
rect 7193 16708 7205 16711
rect 6512 16680 7205 16708
rect 6512 16668 6518 16680
rect 7193 16677 7205 16680
rect 7239 16677 7251 16711
rect 7193 16671 7251 16677
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 12066 16708 12072 16720
rect 8352 16680 12072 16708
rect 8352 16668 8358 16680
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 14829 16711 14887 16717
rect 14829 16677 14841 16711
rect 14875 16708 14887 16711
rect 15194 16708 15200 16720
rect 14875 16680 15200 16708
rect 14875 16677 14887 16680
rect 14829 16671 14887 16677
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 16669 16711 16727 16717
rect 16669 16677 16681 16711
rect 16715 16708 16727 16711
rect 17494 16708 17500 16720
rect 16715 16680 17500 16708
rect 16715 16677 16727 16680
rect 16669 16671 16727 16677
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 31294 16708 31300 16720
rect 29932 16680 31300 16708
rect 2648 16612 4292 16640
rect 5920 16612 6684 16640
rect 2648 16600 2654 16612
rect 4264 16581 4292 16612
rect 6656 16584 6684 16612
rect 7098 16600 7104 16652
rect 7156 16600 7162 16652
rect 7322 16643 7380 16649
rect 7322 16640 7334 16643
rect 7208 16612 7334 16640
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3108 16476 3433 16504
rect 3108 16464 3114 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 4080 16504 4108 16535
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 7208 16572 7236 16612
rect 7322 16609 7334 16612
rect 7368 16640 7380 16643
rect 9858 16640 9864 16652
rect 7368 16612 9864 16640
rect 7368 16609 7380 16612
rect 7322 16603 7380 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10410 16640 10416 16652
rect 9968 16612 10416 16640
rect 6696 16544 7236 16572
rect 6696 16532 6702 16544
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 9968 16581 9996 16612
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 12084 16640 12112 16668
rect 12084 16612 12204 16640
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16541 10011 16575
rect 9953 16535 10011 16541
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 12176 16581 12204 16612
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 14792 16612 15301 16640
rect 14792 16600 14798 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 26142 16600 26148 16652
rect 26200 16640 26206 16652
rect 28902 16640 28908 16652
rect 26200 16612 26556 16640
rect 26200 16600 26206 16612
rect 12161 16575 12219 16581
rect 10100 16544 10143 16572
rect 10100 16532 10106 16544
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16566 12403 16575
rect 12452 16566 12480 16600
rect 12391 16541 12480 16566
rect 12345 16538 12480 16541
rect 12345 16535 12403 16538
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 15378 16572 15384 16584
rect 14691 16544 15384 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15556 16575 15614 16581
rect 15556 16541 15568 16575
rect 15602 16572 15614 16575
rect 16574 16572 16580 16584
rect 15602 16544 16580 16572
rect 15602 16541 15614 16544
rect 15556 16535 15614 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 17328 16544 18337 16572
rect 5074 16504 5080 16516
rect 4080 16476 5080 16504
rect 3421 16467 3479 16473
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 6546 16504 6552 16516
rect 5583 16476 6552 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 6546 16464 6552 16476
rect 6604 16504 6610 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 6604 16476 7481 16504
rect 6604 16464 6610 16476
rect 7469 16473 7481 16476
rect 7515 16504 7527 16507
rect 11146 16504 11152 16516
rect 7515 16476 11152 16504
rect 7515 16473 7527 16476
rect 7469 16467 7527 16473
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16504 14519 16507
rect 17034 16504 17040 16516
rect 14507 16476 17040 16504
rect 14507 16473 14519 16476
rect 14461 16467 14519 16473
rect 17034 16464 17040 16476
rect 17092 16464 17098 16516
rect 3221 16439 3279 16445
rect 3221 16405 3233 16439
rect 3267 16436 3279 16439
rect 5997 16439 6055 16445
rect 5997 16436 6009 16439
rect 3267 16408 6009 16436
rect 3267 16405 3279 16408
rect 3221 16399 3279 16405
rect 5997 16405 6009 16408
rect 6043 16436 6055 16439
rect 6362 16436 6368 16448
rect 6043 16408 6368 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7650 16436 7656 16448
rect 7156 16408 7656 16436
rect 7156 16396 7162 16408
rect 7650 16396 7656 16408
rect 7708 16436 7714 16448
rect 9674 16436 9680 16448
rect 7708 16408 9680 16436
rect 7708 16396 7714 16408
rect 9674 16396 9680 16408
rect 9732 16436 9738 16448
rect 10134 16436 10140 16448
rect 9732 16408 10140 16436
rect 9732 16396 9738 16408
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10229 16439 10287 16445
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10410 16436 10416 16448
rect 10275 16408 10416 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15930 16436 15936 16448
rect 15436 16408 15936 16436
rect 15436 16396 15442 16408
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 16114 16396 16120 16448
rect 16172 16436 16178 16448
rect 17328 16436 17356 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16572 19487 16575
rect 19518 16572 19524 16584
rect 19475 16544 19524 16572
rect 19475 16541 19487 16544
rect 19429 16535 19487 16541
rect 17402 16464 17408 16516
rect 17460 16504 17466 16516
rect 17589 16507 17647 16513
rect 17589 16504 17601 16507
rect 17460 16476 17601 16504
rect 17460 16464 17466 16476
rect 17589 16473 17601 16476
rect 17635 16473 17647 16507
rect 18524 16504 18552 16535
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 19696 16575 19754 16581
rect 19696 16541 19708 16575
rect 19742 16572 19754 16575
rect 20438 16572 20444 16584
rect 19742 16544 20444 16572
rect 19742 16541 19754 16544
rect 19696 16535 19754 16541
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16572 21603 16575
rect 23290 16572 23296 16584
rect 21591 16544 23296 16572
rect 21591 16541 21603 16544
rect 21545 16535 21603 16541
rect 17589 16467 17647 16473
rect 17880 16476 18552 16504
rect 16172 16408 17356 16436
rect 16172 16396 16178 16408
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 17880 16436 17908 16476
rect 18690 16464 18696 16516
rect 18748 16464 18754 16516
rect 19242 16464 19248 16516
rect 19300 16504 19306 16516
rect 21560 16504 21588 16535
rect 23290 16532 23296 16544
rect 23348 16572 23354 16584
rect 23348 16544 23980 16572
rect 23348 16532 23354 16544
rect 19300 16476 21588 16504
rect 19300 16464 19306 16476
rect 21634 16464 21640 16516
rect 21692 16504 21698 16516
rect 23952 16504 23980 16544
rect 24578 16532 24584 16584
rect 24636 16532 24642 16584
rect 24854 16581 24860 16584
rect 24848 16572 24860 16581
rect 24815 16544 24860 16572
rect 24848 16535 24860 16544
rect 24854 16532 24860 16535
rect 24912 16532 24918 16584
rect 26421 16575 26479 16581
rect 26421 16541 26433 16575
rect 26467 16541 26479 16575
rect 26528 16572 26556 16612
rect 28736 16612 28908 16640
rect 26697 16575 26755 16581
rect 26697 16572 26709 16575
rect 26528 16544 26709 16572
rect 26421 16535 26479 16541
rect 26697 16541 26709 16544
rect 26743 16572 26755 16575
rect 28736 16572 28764 16612
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 29086 16600 29092 16652
rect 29144 16640 29150 16652
rect 29730 16640 29736 16652
rect 29144 16612 29736 16640
rect 29144 16600 29150 16612
rect 29730 16600 29736 16612
rect 29788 16600 29794 16652
rect 29932 16581 29960 16680
rect 31294 16668 31300 16680
rect 31352 16668 31358 16720
rect 30006 16600 30012 16652
rect 30064 16640 30070 16652
rect 31386 16640 31392 16652
rect 30064 16612 31392 16640
rect 30064 16600 30070 16612
rect 31386 16600 31392 16612
rect 31444 16640 31450 16652
rect 31444 16612 31524 16640
rect 31444 16600 31450 16612
rect 26743 16544 28764 16572
rect 29917 16575 29975 16581
rect 26743 16541 26755 16544
rect 26697 16535 26755 16541
rect 29917 16541 29929 16575
rect 29963 16541 29975 16575
rect 29917 16535 29975 16541
rect 31205 16575 31263 16581
rect 31205 16541 31217 16575
rect 31251 16572 31263 16575
rect 31294 16572 31300 16584
rect 31251 16544 31300 16572
rect 31251 16541 31263 16544
rect 31205 16535 31263 16541
rect 26436 16504 26464 16535
rect 28350 16504 28356 16516
rect 21692 16476 22094 16504
rect 23952 16476 26464 16504
rect 27540 16476 28356 16504
rect 21692 16464 21698 16476
rect 17736 16408 17908 16436
rect 20809 16439 20867 16445
rect 17736 16396 17742 16408
rect 20809 16405 20821 16439
rect 20855 16436 20867 16439
rect 21174 16436 21180 16448
rect 20855 16408 21180 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 22066 16436 22094 16476
rect 26142 16436 26148 16448
rect 22066 16408 26148 16436
rect 26142 16396 26148 16408
rect 26200 16436 26206 16448
rect 27540 16436 27568 16476
rect 28350 16464 28356 16476
rect 28408 16464 28414 16516
rect 28718 16464 28724 16516
rect 28776 16504 28782 16516
rect 29932 16504 29960 16535
rect 31294 16532 31300 16544
rect 31352 16532 31358 16584
rect 31496 16581 31524 16612
rect 32306 16600 32312 16652
rect 32364 16640 32370 16652
rect 32585 16643 32643 16649
rect 32585 16640 32597 16643
rect 32364 16612 32597 16640
rect 32364 16600 32370 16612
rect 32585 16609 32597 16612
rect 32631 16640 32643 16643
rect 32766 16640 32772 16652
rect 32631 16612 32772 16640
rect 32631 16609 32643 16612
rect 32585 16603 32643 16609
rect 32766 16600 32772 16612
rect 32824 16600 32830 16652
rect 31481 16575 31539 16581
rect 31481 16541 31493 16575
rect 31527 16541 31539 16575
rect 31481 16535 31539 16541
rect 31609 16575 31667 16581
rect 31609 16541 31621 16575
rect 31655 16572 31667 16575
rect 32324 16572 32352 16600
rect 31655 16544 32352 16572
rect 31655 16541 31667 16544
rect 31609 16535 31667 16541
rect 32398 16532 32404 16584
rect 32456 16532 32462 16584
rect 31389 16507 31447 16513
rect 31389 16504 31401 16507
rect 28776 16476 29960 16504
rect 30116 16476 31401 16504
rect 28776 16464 28782 16476
rect 30116 16448 30144 16476
rect 31389 16473 31401 16476
rect 31435 16473 31447 16507
rect 31389 16467 31447 16473
rect 26200 16408 27568 16436
rect 26200 16396 26206 16408
rect 27798 16396 27804 16448
rect 27856 16436 27862 16448
rect 28442 16436 28448 16448
rect 27856 16408 28448 16436
rect 27856 16396 27862 16408
rect 28442 16396 28448 16408
rect 28500 16436 28506 16448
rect 30006 16436 30012 16448
rect 28500 16408 30012 16436
rect 28500 16396 28506 16408
rect 30006 16396 30012 16408
rect 30064 16396 30070 16448
rect 30098 16396 30104 16448
rect 30156 16396 30162 16448
rect 30282 16396 30288 16448
rect 30340 16396 30346 16448
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 6730 16192 6736 16244
rect 6788 16192 6794 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 12768 16204 13461 16232
rect 12768 16192 12774 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 19242 16232 19248 16244
rect 13449 16195 13507 16201
rect 14016 16204 19248 16232
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 6822 16164 6828 16176
rect 5776 16136 6828 16164
rect 5776 16124 5782 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 6454 16096 6460 16108
rect 5583 16068 6460 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 6696 16068 6745 16096
rect 6696 16056 6702 16068
rect 6733 16065 6745 16068
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9585 16099 9643 16105
rect 9585 16096 9597 16099
rect 9364 16068 9597 16096
rect 9364 16056 9370 16068
rect 9585 16065 9597 16068
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13464 16096 13492 16195
rect 14016 16105 14044 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19518 16192 19524 16244
rect 19576 16192 19582 16244
rect 20441 16235 20499 16241
rect 20441 16201 20453 16235
rect 20487 16232 20499 16235
rect 20530 16232 20536 16244
rect 20487 16204 20536 16232
rect 20487 16201 20499 16204
rect 20441 16195 20499 16201
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20824 16204 22324 16232
rect 15194 16173 15200 16176
rect 15188 16164 15200 16173
rect 15155 16136 15200 16164
rect 15188 16127 15200 16136
rect 15194 16124 15200 16127
rect 15252 16124 15258 16176
rect 18230 16124 18236 16176
rect 18288 16124 18294 16176
rect 18690 16124 18696 16176
rect 18748 16164 18754 16176
rect 20824 16173 20852 16204
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 18748 16136 20821 16164
rect 18748 16124 18754 16136
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 22296 16173 22324 16204
rect 22646 16192 22652 16244
rect 22704 16192 22710 16244
rect 24486 16192 24492 16244
rect 24544 16232 24550 16244
rect 28718 16232 28724 16244
rect 24544 16204 28396 16232
rect 24544 16192 24550 16204
rect 22281 16167 22339 16173
rect 21232 16136 22140 16164
rect 21232 16124 21238 16136
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13464 16068 14013 16096
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14366 16096 14372 16108
rect 14323 16068 14372 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14366 16056 14372 16068
rect 14424 16096 14430 16108
rect 16206 16096 16212 16108
rect 14424 16068 16212 16096
rect 14424 16056 14430 16068
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 7098 16028 7104 16040
rect 5399 16000 7104 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 5552 15972 5580 16000
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14792 16000 14933 16028
rect 14792 15988 14798 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 17052 16028 17080 16059
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20579 16099 20637 16105
rect 20579 16096 20591 16099
rect 20312 16068 20591 16096
rect 20312 16056 20318 16068
rect 20579 16065 20591 16068
rect 20625 16065 20637 16099
rect 20579 16059 20637 16065
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 16448 16000 17080 16028
rect 17405 16031 17463 16037
rect 16448 15988 16454 16000
rect 17405 15997 17417 16031
rect 17451 16028 17463 16031
rect 20162 16028 20168 16040
rect 17451 16000 20168 16028
rect 17451 15997 17463 16000
rect 17405 15991 17463 15997
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 5534 15920 5540 15972
rect 5592 15920 5598 15972
rect 15930 15920 15936 15972
rect 15988 15960 15994 15972
rect 20732 15960 20760 16059
rect 20898 16056 20904 16108
rect 20956 16105 20962 16108
rect 20956 16099 20995 16105
rect 20983 16065 20995 16099
rect 20956 16059 20995 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16096 21143 16099
rect 21818 16096 21824 16108
rect 21131 16068 21824 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 20956 16056 20962 16059
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 22112 16105 22140 16136
rect 22281 16133 22293 16167
rect 22327 16133 22339 16167
rect 22281 16127 22339 16133
rect 26050 16124 26056 16176
rect 26108 16164 26114 16176
rect 26513 16167 26571 16173
rect 26513 16164 26525 16167
rect 26108 16136 26525 16164
rect 26108 16124 26114 16136
rect 26513 16133 26525 16136
rect 26559 16133 26571 16167
rect 26513 16127 26571 16133
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22098 16099 22156 16105
rect 22098 16065 22110 16099
rect 22144 16065 22156 16099
rect 22098 16059 22156 16065
rect 22020 16028 22048 16059
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22511 16099 22569 16105
rect 22511 16065 22523 16099
rect 22557 16096 22569 16099
rect 22830 16096 22836 16108
rect 22557 16068 22836 16096
rect 22557 16065 22569 16068
rect 22511 16059 22569 16065
rect 22830 16056 22836 16068
rect 22888 16056 22894 16108
rect 25130 16056 25136 16108
rect 25188 16056 25194 16108
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 26329 16099 26387 16105
rect 26329 16096 26341 16099
rect 26200 16068 26341 16096
rect 26200 16056 26206 16068
rect 26329 16065 26341 16068
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26602 16056 26608 16108
rect 26660 16056 26666 16108
rect 27982 16028 27988 16040
rect 22020 16000 27988 16028
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 28368 16028 28396 16204
rect 28644 16204 28724 16232
rect 28644 16173 28672 16204
rect 28718 16192 28724 16204
rect 28776 16192 28782 16244
rect 32766 16192 32772 16244
rect 32824 16232 32830 16244
rect 33689 16235 33747 16241
rect 33689 16232 33701 16235
rect 32824 16204 33701 16232
rect 32824 16192 32830 16204
rect 33689 16201 33701 16204
rect 33735 16201 33747 16235
rect 33689 16195 33747 16201
rect 28629 16167 28687 16173
rect 28629 16133 28641 16167
rect 28675 16133 28687 16167
rect 30098 16164 30104 16176
rect 28629 16127 28687 16133
rect 28736 16136 30104 16164
rect 28442 16056 28448 16108
rect 28500 16096 28506 16108
rect 28736 16105 28764 16136
rect 30098 16124 30104 16136
rect 30156 16164 30162 16176
rect 30156 16136 31754 16164
rect 30156 16124 30162 16136
rect 28537 16099 28595 16105
rect 28537 16096 28549 16099
rect 28500 16068 28549 16096
rect 28500 16056 28506 16068
rect 28537 16065 28549 16068
rect 28583 16065 28595 16099
rect 28537 16059 28595 16065
rect 28721 16099 28779 16105
rect 28721 16065 28733 16099
rect 28767 16065 28779 16099
rect 28721 16059 28779 16065
rect 28736 16028 28764 16059
rect 28902 16056 28908 16108
rect 28960 16096 28966 16108
rect 29086 16096 29092 16108
rect 28960 16068 29092 16096
rect 28960 16056 28966 16068
rect 29086 16056 29092 16068
rect 29144 16056 29150 16108
rect 29549 16099 29607 16105
rect 29549 16065 29561 16099
rect 29595 16096 29607 16099
rect 30282 16096 30288 16108
rect 29595 16068 30288 16096
rect 29595 16065 29607 16068
rect 29549 16059 29607 16065
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 28368 16000 28764 16028
rect 31726 16028 31754 16136
rect 32398 16096 32404 16108
rect 32232 16068 32404 16096
rect 32232 16028 32260 16068
rect 32398 16056 32404 16068
rect 32456 16056 32462 16108
rect 32576 16099 32634 16105
rect 32576 16065 32588 16099
rect 32622 16096 32634 16099
rect 33870 16096 33876 16108
rect 32622 16068 33876 16096
rect 32622 16065 32634 16068
rect 32576 16059 32634 16065
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 31726 16000 32260 16028
rect 32306 15988 32312 16040
rect 32364 15988 32370 16040
rect 26050 15960 26056 15972
rect 15988 15932 19472 15960
rect 20732 15932 26056 15960
rect 15988 15920 15994 15932
rect 19444 15904 19472 15932
rect 26050 15920 26056 15932
rect 26108 15920 26114 15972
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 17034 15892 17040 15904
rect 16347 15864 17040 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 21634 15892 21640 15904
rect 19484 15864 21640 15892
rect 19484 15852 19490 15864
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 24578 15892 24584 15904
rect 23891 15864 24584 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 26142 15852 26148 15904
rect 26200 15852 26206 15904
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 28224 15864 28365 15892
rect 28224 15852 28230 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 28353 15855 28411 15861
rect 29454 15852 29460 15904
rect 29512 15852 29518 15904
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 4982 15648 4988 15700
rect 5040 15688 5046 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 5040 15660 5273 15688
rect 5040 15648 5046 15660
rect 5261 15657 5273 15660
rect 5307 15688 5319 15691
rect 7742 15688 7748 15700
rect 5307 15660 7748 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 11606 15688 11612 15700
rect 9263 15660 11612 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 23753 15691 23811 15697
rect 23753 15657 23765 15691
rect 23799 15688 23811 15691
rect 23842 15688 23848 15700
rect 23799 15660 23848 15688
rect 23799 15657 23811 15660
rect 23753 15651 23811 15657
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 26050 15688 26056 15700
rect 25188 15660 26056 15688
rect 25188 15648 25194 15660
rect 26050 15648 26056 15660
rect 26108 15688 26114 15700
rect 26513 15691 26571 15697
rect 26513 15688 26525 15691
rect 26108 15660 26525 15688
rect 26108 15648 26114 15660
rect 26513 15657 26525 15660
rect 26559 15657 26571 15691
rect 26513 15651 26571 15657
rect 27982 15648 27988 15700
rect 28040 15648 28046 15700
rect 31665 15691 31723 15697
rect 31665 15657 31677 15691
rect 31711 15688 31723 15691
rect 31754 15688 31760 15700
rect 31711 15660 31760 15688
rect 31711 15657 31723 15660
rect 31665 15651 31723 15657
rect 31754 15648 31760 15660
rect 31812 15688 31818 15700
rect 32306 15688 32312 15700
rect 31812 15660 32312 15688
rect 31812 15648 31818 15660
rect 32306 15648 32312 15660
rect 32364 15648 32370 15700
rect 33870 15648 33876 15700
rect 33928 15648 33934 15700
rect 7929 15623 7987 15629
rect 7929 15589 7941 15623
rect 7975 15620 7987 15623
rect 13262 15620 13268 15632
rect 7975 15592 13268 15620
rect 7975 15589 7987 15592
rect 7929 15583 7987 15589
rect 13262 15580 13268 15592
rect 13320 15580 13326 15632
rect 13633 15623 13691 15629
rect 13633 15589 13645 15623
rect 13679 15620 13691 15623
rect 15102 15620 15108 15632
rect 13679 15592 15108 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 32674 15620 32680 15632
rect 22428 15592 32680 15620
rect 22428 15580 22434 15592
rect 32674 15580 32680 15592
rect 32732 15580 32738 15632
rect 6638 15552 6644 15564
rect 6104 15524 6644 15552
rect 2590 15444 2596 15496
rect 2648 15444 2654 15496
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 5074 15484 5080 15496
rect 2915 15456 5080 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6104 15493 6132 15524
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 7650 15512 7656 15564
rect 7708 15512 7714 15564
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 10652 15524 12434 15552
rect 10652 15512 10658 15524
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5868 15456 6101 15484
rect 5868 15444 5874 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6546 15484 6552 15496
rect 6319 15456 6552 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 6730 15444 6736 15496
rect 6788 15444 6794 15496
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 2958 15376 2964 15428
rect 3016 15376 3022 15428
rect 5445 15419 5503 15425
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 5534 15416 5540 15428
rect 5491 15388 5540 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 7392 15416 7420 15447
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 7524 15456 9137 15484
rect 7524 15444 7530 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 11146 15444 11152 15496
rect 11204 15444 11210 15496
rect 12406 15484 12434 15524
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 13504 15524 14933 15552
rect 13504 15512 13510 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 16390 15552 16396 15564
rect 14921 15515 14979 15521
rect 15672 15524 16396 15552
rect 15672 15496 15700 15524
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 12406 15456 12541 15484
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12667 15456 13369 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 14366 15484 14372 15496
rect 13679 15456 14372 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14608 15456 15025 15484
rect 14608 15444 14614 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15484 15347 15487
rect 15654 15484 15660 15496
rect 15335 15456 15660 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 16316 15493 16344 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 19150 15552 19156 15564
rect 18279 15524 19156 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 22554 15512 22560 15564
rect 22612 15512 22618 15564
rect 25774 15552 25780 15564
rect 22664 15524 25780 15552
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 17678 15444 17684 15496
rect 17736 15444 17742 15496
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 6196 15388 7420 15416
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 4488 15320 5089 15348
rect 4488 15308 4494 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 5245 15351 5303 15357
rect 5245 15317 5257 15351
rect 5291 15348 5303 15351
rect 6086 15348 6092 15360
rect 5291 15320 6092 15348
rect 5291 15317 5303 15320
rect 5245 15311 5303 15317
rect 6086 15308 6092 15320
rect 6144 15348 6150 15360
rect 6196 15357 6224 15388
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 17880 15416 17908 15447
rect 20806 15444 20812 15496
rect 20864 15444 20870 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22664 15484 22692 15524
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 28166 15512 28172 15564
rect 28224 15512 28230 15564
rect 28353 15555 28411 15561
rect 28353 15521 28365 15555
rect 28399 15552 28411 15555
rect 29454 15552 29460 15564
rect 28399 15524 29460 15552
rect 28399 15521 28411 15524
rect 28353 15515 28411 15521
rect 29454 15512 29460 15524
rect 29512 15512 29518 15564
rect 31726 15524 33732 15552
rect 22244 15456 22692 15484
rect 24029 15487 24087 15493
rect 22244 15444 22250 15456
rect 24029 15453 24041 15487
rect 24075 15484 24087 15487
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24075 15456 25237 15484
rect 24075 15453 24087 15456
rect 24029 15447 24087 15453
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 27706 15484 27712 15496
rect 25225 15447 25283 15453
rect 25700 15456 27712 15484
rect 17644 15388 17908 15416
rect 17644 15376 17650 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 21910 15416 21916 15428
rect 19392 15388 21916 15416
rect 19392 15376 19398 15388
rect 21910 15376 21916 15388
rect 21968 15416 21974 15428
rect 23569 15419 23627 15425
rect 23569 15416 23581 15419
rect 21968 15388 23581 15416
rect 21968 15376 21974 15388
rect 23569 15385 23581 15388
rect 23615 15385 23627 15419
rect 23569 15379 23627 15385
rect 24394 15376 24400 15428
rect 24452 15416 24458 15428
rect 25700 15416 25728 15456
rect 27706 15444 27712 15456
rect 27764 15484 27770 15496
rect 28074 15484 28080 15496
rect 27764 15456 28080 15484
rect 27764 15444 27770 15456
rect 28074 15444 28080 15456
rect 28132 15484 28138 15496
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 28132 15456 28273 15484
rect 28132 15444 28138 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28442 15444 28448 15496
rect 28500 15444 28506 15496
rect 24452 15388 25728 15416
rect 24452 15376 24458 15388
rect 25774 15376 25780 15428
rect 25832 15416 25838 15428
rect 29546 15416 29552 15428
rect 25832 15388 29552 15416
rect 25832 15376 25838 15388
rect 29546 15376 29552 15388
rect 29604 15416 29610 15428
rect 31726 15416 31754 15524
rect 32858 15444 32864 15496
rect 32916 15484 32922 15496
rect 33704 15493 33732 15524
rect 33413 15487 33471 15493
rect 33413 15484 33425 15487
rect 32916 15456 33425 15484
rect 32916 15444 32922 15456
rect 33413 15453 33425 15456
rect 33459 15453 33471 15487
rect 33413 15447 33471 15453
rect 33689 15487 33747 15493
rect 33689 15453 33701 15487
rect 33735 15453 33747 15487
rect 33689 15447 33747 15453
rect 29604 15388 31754 15416
rect 29604 15376 29610 15388
rect 32950 15376 32956 15428
rect 33008 15376 33014 15428
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 6144 15320 6193 15348
rect 6144 15308 6150 15320
rect 6181 15317 6193 15320
rect 6227 15317 6239 15351
rect 6181 15311 6239 15317
rect 6822 15308 6828 15360
rect 6880 15308 6886 15360
rect 10965 15351 11023 15357
rect 10965 15317 10977 15351
rect 11011 15348 11023 15351
rect 12526 15348 12532 15360
rect 11011 15320 12532 15348
rect 11011 15317 11023 15320
rect 10965 15311 11023 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 16298 15308 16304 15360
rect 16356 15308 16362 15360
rect 23750 15308 23756 15360
rect 23808 15348 23814 15360
rect 24762 15348 24768 15360
rect 23808 15320 24768 15348
rect 23808 15308 23814 15320
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 32766 15308 32772 15360
rect 32824 15348 32830 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 32824 15320 33517 15348
rect 32824 15308 32830 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33505 15311 33563 15317
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 5436 15147 5494 15153
rect 5436 15113 5448 15147
rect 5482 15144 5494 15147
rect 5718 15144 5724 15156
rect 5482 15116 5724 15144
rect 5482 15113 5494 15116
rect 5436 15107 5494 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 9125 15147 9183 15153
rect 9125 15144 9137 15147
rect 8536 15116 9137 15144
rect 8536 15104 8542 15116
rect 9125 15113 9137 15116
rect 9171 15113 9183 15147
rect 9125 15107 9183 15113
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 16025 15147 16083 15153
rect 10008 15116 12434 15144
rect 10008 15104 10014 15116
rect 2958 15036 2964 15088
rect 3016 15036 3022 15088
rect 5810 15036 5816 15088
rect 5868 15036 5874 15088
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 12406 15076 12434 15116
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16482 15144 16488 15156
rect 16071 15116 16488 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 22373 15147 22431 15153
rect 17184 15116 18368 15144
rect 17184 15104 17190 15116
rect 12710 15076 12716 15088
rect 9079 15048 10732 15076
rect 12406 15048 12716 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 10704 15020 10732 15048
rect 12710 15036 12716 15048
rect 12768 15036 12774 15088
rect 17678 15076 17684 15088
rect 17328 15048 17684 15076
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4522 15008 4528 15020
rect 4203 14980 4528 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2682 14940 2688 14952
rect 1995 14912 2688 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2682 14900 2688 14912
rect 2740 14940 2746 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 2740 14912 4077 14940
rect 2740 14900 2746 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 3234 14832 3240 14884
rect 3292 14872 3298 14884
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3292 14844 3433 14872
rect 3292 14832 3298 14844
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 4172 14872 4200 14971
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 9950 15008 9956 15020
rect 9355 14980 9956 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 10376 14980 10425 15008
rect 10376 14968 10382 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 3467 14844 4200 14872
rect 10428 14872 10456 14971
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15712 14980 16129 15008
rect 15712 14968 15718 14980
rect 16117 14977 16129 14980
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16850 15008 16856 15020
rect 16347 14980 16856 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 17328 15017 17356 15048
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 12066 14940 12072 14952
rect 11195 14912 12072 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 17512 14940 17540 14971
rect 18230 14968 18236 15020
rect 18288 14968 18294 15020
rect 18340 15008 18368 15116
rect 22373 15113 22385 15147
rect 22419 15144 22431 15147
rect 22462 15144 22468 15156
rect 22419 15116 22468 15144
rect 22419 15113 22431 15116
rect 22373 15107 22431 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 32950 15104 32956 15156
rect 33008 15144 33014 15156
rect 33597 15147 33655 15153
rect 33597 15144 33609 15147
rect 33008 15116 33609 15144
rect 33008 15104 33014 15116
rect 33597 15113 33609 15116
rect 33643 15113 33655 15147
rect 33597 15107 33655 15113
rect 23934 15076 23940 15088
rect 20640 15048 23940 15076
rect 20640 15017 20668 15048
rect 23934 15036 23940 15048
rect 23992 15076 23998 15088
rect 24762 15076 24768 15088
rect 23992 15048 24768 15076
rect 23992 15036 23998 15048
rect 24762 15036 24768 15048
rect 24820 15076 24826 15088
rect 30834 15076 30840 15088
rect 24820 15048 30840 15076
rect 24820 15036 24826 15048
rect 30834 15036 30840 15048
rect 30892 15036 30898 15088
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 18340 14980 20637 15008
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20806 14968 20812 15020
rect 20864 14968 20870 15020
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 22186 14968 22192 15020
rect 22244 14968 22250 15020
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 22296 14980 22477 15008
rect 16632 14912 17540 14940
rect 17773 14943 17831 14949
rect 16632 14900 16638 14912
rect 17773 14909 17785 14943
rect 17819 14909 17831 14943
rect 20916 14940 20944 14968
rect 22296 14940 22324 14980
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 25130 14968 25136 15020
rect 25188 15017 25194 15020
rect 25188 14971 25200 15017
rect 25188 14968 25194 14971
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 29825 15011 29883 15017
rect 29825 15008 29837 15011
rect 29052 14980 29837 15008
rect 29052 14968 29058 14980
rect 29825 14977 29837 14980
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 29914 14968 29920 15020
rect 29972 15008 29978 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 29972 14980 32321 15008
rect 29972 14968 29978 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 20916 14912 22324 14940
rect 25409 14943 25467 14949
rect 17773 14903 17831 14909
rect 25409 14909 25421 14943
rect 25455 14940 25467 14943
rect 26418 14940 26424 14952
rect 25455 14912 26424 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 13262 14872 13268 14884
rect 10428 14844 13268 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 17788 14872 17816 14903
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 24394 14872 24400 14884
rect 17788 14844 24400 14872
rect 24394 14832 24400 14844
rect 24452 14832 24458 14884
rect 29638 14832 29644 14884
rect 29696 14832 29702 14884
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 4304 14776 5273 14804
rect 4304 14764 4310 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 6546 14804 6552 14816
rect 5491 14776 6552 14804
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14804 9643 14807
rect 11974 14804 11980 14816
rect 9631 14776 11980 14804
rect 9631 14773 9643 14776
rect 9585 14767 9643 14773
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 19702 14764 19708 14816
rect 19760 14764 19766 14816
rect 20438 14764 20444 14816
rect 20496 14764 20502 14816
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 21048 14776 22017 14804
rect 21048 14764 21054 14776
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 22005 14767 22063 14773
rect 24026 14764 24032 14816
rect 24084 14764 24090 14816
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6822 14600 6828 14612
rect 6227 14572 6828 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 9122 14600 9128 14612
rect 7423 14572 9128 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 6086 14492 6092 14544
rect 6144 14532 6150 14544
rect 7208 14532 7236 14563
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 19886 14600 19892 14612
rect 19659 14572 19892 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 22097 14603 22155 14609
rect 20272 14572 21680 14600
rect 20272 14544 20300 14572
rect 6144 14504 7236 14532
rect 6144 14492 6150 14504
rect 8478 14492 8484 14544
rect 8536 14492 8542 14544
rect 8846 14492 8852 14544
rect 8904 14532 8910 14544
rect 9217 14535 9275 14541
rect 9217 14532 9229 14535
rect 8904 14504 9229 14532
rect 8904 14492 8910 14504
rect 9217 14501 9229 14504
rect 9263 14501 9275 14535
rect 9217 14495 9275 14501
rect 9306 14492 9312 14544
rect 9364 14532 9370 14544
rect 18049 14535 18107 14541
rect 9364 14504 17356 14532
rect 9364 14492 9370 14504
rect 1762 14424 1768 14476
rect 1820 14464 1826 14476
rect 17328 14473 17356 14504
rect 18049 14501 18061 14535
rect 18095 14532 18107 14535
rect 20254 14532 20260 14544
rect 18095 14504 20260 14532
rect 18095 14501 18107 14504
rect 18049 14495 18107 14501
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 21652 14532 21680 14572
rect 22097 14569 22109 14603
rect 22143 14600 22155 14603
rect 22462 14600 22468 14612
rect 22143 14572 22468 14600
rect 22143 14569 22155 14572
rect 22097 14563 22155 14569
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 25958 14560 25964 14612
rect 26016 14560 26022 14612
rect 22186 14532 22192 14544
rect 21652 14504 22192 14532
rect 22186 14492 22192 14504
rect 22244 14532 22250 14544
rect 23750 14532 23756 14544
rect 22244 14504 23756 14532
rect 22244 14492 22250 14504
rect 23750 14492 23756 14504
rect 23808 14492 23814 14544
rect 17313 14467 17371 14473
rect 1820 14436 7236 14464
rect 1820 14424 1826 14436
rect 2682 14356 2688 14408
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3050 14396 3056 14408
rect 2915 14368 3056 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 7208 14396 7236 14436
rect 7484 14436 15608 14464
rect 7484 14396 7512 14436
rect 7208 14368 7512 14396
rect 6365 14359 6423 14365
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14297 3019 14331
rect 2961 14291 3019 14297
rect 2976 14260 3004 14291
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 6380 14328 6408 14359
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8168 14368 9076 14396
rect 8168 14356 8174 14368
rect 6454 14328 6460 14340
rect 5776 14300 6460 14328
rect 5776 14288 5782 14300
rect 6454 14288 6460 14300
rect 6512 14328 6518 14340
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6512 14300 7021 14328
rect 6512 14288 6518 14300
rect 7009 14297 7021 14300
rect 7055 14297 7067 14331
rect 7009 14291 7067 14297
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 7225 14331 7283 14337
rect 7225 14328 7237 14331
rect 7156 14300 7237 14328
rect 7156 14288 7162 14300
rect 7225 14297 7237 14300
rect 7271 14328 7283 14331
rect 7466 14328 7472 14340
rect 7271 14300 7472 14328
rect 7271 14297 7283 14300
rect 7225 14291 7283 14297
rect 7466 14288 7472 14300
rect 7524 14288 7530 14340
rect 7926 14288 7932 14340
rect 7984 14328 7990 14340
rect 8205 14331 8263 14337
rect 7984 14300 8156 14328
rect 7984 14288 7990 14300
rect 3786 14260 3792 14272
rect 2976 14232 3792 14260
rect 3786 14220 3792 14232
rect 3844 14260 3850 14272
rect 5810 14260 5816 14272
rect 3844 14232 5816 14260
rect 3844 14220 3850 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 6914 14260 6920 14272
rect 6595 14232 6920 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7892 14232 8033 14260
rect 7892 14220 7898 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8128 14260 8156 14300
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8570 14328 8576 14340
rect 8251 14300 8576 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 9048 14328 9076 14368
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 12802 14396 12808 14408
rect 9272 14368 12808 14396
rect 9272 14356 9278 14368
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13722 14396 13728 14408
rect 12943 14368 13728 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 9490 14328 9496 14340
rect 9048 14300 9496 14328
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 9769 14331 9827 14337
rect 9769 14328 9781 14331
rect 9600 14300 9781 14328
rect 9600 14260 9628 14300
rect 9769 14297 9781 14300
rect 9815 14328 9827 14331
rect 10686 14328 10692 14340
rect 9815 14300 10692 14328
rect 9815 14297 9827 14300
rect 9769 14291 9827 14297
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12912 14328 12940 14359
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 15580 14405 15608 14436
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 20530 14464 20536 14476
rect 17359 14436 20536 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 24578 14424 24584 14476
rect 24636 14424 24642 14476
rect 31389 14467 31447 14473
rect 31389 14433 31401 14467
rect 31435 14464 31447 14467
rect 31754 14464 31760 14476
rect 31435 14436 31760 14464
rect 31435 14433 31447 14436
rect 31389 14427 31447 14433
rect 31754 14424 31760 14436
rect 31812 14424 31818 14476
rect 31849 14467 31907 14473
rect 31849 14433 31861 14467
rect 31895 14464 31907 14467
rect 32306 14464 32312 14476
rect 31895 14436 32312 14464
rect 31895 14433 31907 14436
rect 31849 14427 31907 14433
rect 32306 14424 32312 14436
rect 32364 14424 32370 14476
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17644 14368 17785 14396
rect 17644 14356 17650 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18414 14396 18420 14408
rect 18095 14368 18420 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20990 14405 20996 14408
rect 20717 14399 20775 14405
rect 20717 14396 20729 14399
rect 19760 14368 20729 14396
rect 19760 14356 19766 14368
rect 20717 14365 20729 14368
rect 20763 14365 20775 14399
rect 20984 14396 20996 14405
rect 20951 14368 20996 14396
rect 20717 14359 20775 14365
rect 20984 14359 20996 14368
rect 20990 14356 20996 14359
rect 21048 14356 21054 14408
rect 24848 14399 24906 14405
rect 24848 14365 24860 14399
rect 24894 14396 24906 14399
rect 26142 14396 26148 14408
rect 24894 14368 26148 14396
rect 24894 14365 24906 14368
rect 24848 14359 24906 14365
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 26418 14356 26424 14408
rect 26476 14396 26482 14408
rect 26970 14396 26976 14408
rect 26476 14368 26976 14396
rect 26476 14356 26482 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 28261 14399 28319 14405
rect 28261 14396 28273 14399
rect 27580 14368 28273 14396
rect 27580 14356 27586 14368
rect 28261 14365 28273 14368
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28534 14356 28540 14408
rect 28592 14356 28598 14408
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 31113 14399 31171 14405
rect 31113 14396 31125 14399
rect 30156 14368 31125 14396
rect 30156 14356 30162 14368
rect 31113 14365 31125 14368
rect 31159 14365 31171 14399
rect 31113 14359 31171 14365
rect 32122 14356 32128 14408
rect 32180 14356 32186 14408
rect 12492 14300 12940 14328
rect 12492 14288 12498 14300
rect 13078 14288 13084 14340
rect 13136 14288 13142 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 19392 14300 19441 14328
rect 19392 14288 19398 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 19518 14288 19524 14340
rect 19576 14328 19582 14340
rect 19613 14331 19671 14337
rect 19613 14328 19625 14331
rect 19576 14300 19625 14328
rect 19576 14288 19582 14300
rect 19613 14297 19625 14300
rect 19659 14328 19671 14331
rect 22738 14328 22744 14340
rect 19659 14300 22744 14328
rect 19659 14297 19671 14300
rect 19613 14291 19671 14297
rect 22738 14288 22744 14300
rect 22796 14288 22802 14340
rect 26688 14331 26746 14337
rect 26688 14297 26700 14331
rect 26734 14328 26746 14331
rect 28721 14331 28779 14337
rect 28721 14328 28733 14331
rect 26734 14300 28733 14328
rect 26734 14297 26746 14300
rect 26688 14291 26746 14297
rect 28721 14297 28733 14300
rect 28767 14297 28779 14331
rect 28721 14291 28779 14297
rect 29730 14288 29736 14340
rect 29788 14288 29794 14340
rect 8128 14232 9628 14260
rect 9677 14263 9735 14269
rect 8021 14223 8079 14229
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 10226 14260 10232 14272
rect 9723 14232 10232 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 19794 14220 19800 14272
rect 19852 14220 19858 14272
rect 19886 14220 19892 14272
rect 19944 14260 19950 14272
rect 23842 14260 23848 14272
rect 19944 14232 23848 14260
rect 19944 14220 19950 14232
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 27798 14220 27804 14272
rect 27856 14260 27862 14272
rect 28353 14263 28411 14269
rect 28353 14260 28365 14263
rect 27856 14232 28365 14260
rect 27856 14220 27862 14232
rect 28353 14229 28365 14232
rect 28399 14229 28411 14263
rect 28353 14223 28411 14229
rect 31294 14220 31300 14272
rect 31352 14260 31358 14272
rect 33226 14260 33232 14272
rect 31352 14232 33232 14260
rect 31352 14220 31358 14232
rect 33226 14220 33232 14232
rect 33284 14220 33290 14272
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 1728 14028 2605 14056
rect 1728 14016 1734 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 7926 14056 7932 14068
rect 5951 14028 7932 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 12434 14056 12440 14068
rect 9784 14028 12440 14056
rect 4430 13948 4436 14000
rect 4488 13948 4494 14000
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6512 13960 6561 13988
rect 6512 13948 6518 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 7098 13988 7104 14000
rect 6779 13960 7104 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3050 13920 3056 13932
rect 2731 13892 3056 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3050 13880 3056 13892
rect 3108 13920 3114 13932
rect 4062 13920 4068 13932
rect 3108 13892 4068 13920
rect 3108 13880 3114 13892
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5810 13880 5816 13932
rect 5868 13920 5874 13932
rect 6748 13920 6776 13951
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 9784 13988 9812 14028
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 12860 14028 14412 14056
rect 12860 14016 12866 14028
rect 7208 13960 9812 13988
rect 7208 13920 7236 13960
rect 5868 13892 6776 13920
rect 6840 13892 7236 13920
rect 5868 13880 5874 13892
rect 4154 13812 4160 13864
rect 4212 13812 4218 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 6840 13852 6868 13892
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9214 13920 9220 13932
rect 8352 13892 9220 13920
rect 8352 13880 8358 13892
rect 9214 13880 9220 13892
rect 9272 13920 9278 13932
rect 9784 13929 9812 13960
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12069 13991 12127 13997
rect 12069 13988 12081 13991
rect 12032 13960 12081 13988
rect 12032 13948 12038 13960
rect 12069 13957 12081 13960
rect 12115 13957 12127 13991
rect 12069 13951 12127 13957
rect 13078 13948 13084 14000
rect 13136 13948 13142 14000
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9272 13892 9505 13920
rect 9272 13880 9278 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14384 13929 14412 14028
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 19886 14056 19892 14068
rect 19076 14028 19892 14056
rect 16960 13988 16988 14016
rect 19076 14000 19104 14028
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 20864 14028 21097 14056
rect 20864 14016 20870 14028
rect 21085 14025 21097 14028
rect 21131 14025 21143 14059
rect 21085 14019 21143 14025
rect 16960 13960 19012 13988
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13780 13892 14197 13920
rect 13780 13880 13786 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 15378 13880 15384 13932
rect 15436 13880 15442 13932
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16301 13923 16359 13929
rect 16301 13920 16313 13923
rect 15988 13892 16313 13920
rect 15988 13880 15994 13892
rect 16301 13889 16313 13892
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 16850 13880 16856 13932
rect 16908 13880 16914 13932
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 17678 13920 17684 13932
rect 17451 13892 17684 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 8386 13852 8392 13864
rect 5132 13824 6868 13852
rect 6932 13824 8392 13852
rect 5132 13812 5138 13824
rect 6932 13793 6960 13824
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 6917 13787 6975 13793
rect 6917 13753 6929 13787
rect 6963 13753 6975 13787
rect 6917 13747 6975 13753
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 10318 13784 10324 13796
rect 8628 13756 10324 13784
rect 8628 13744 8634 13756
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 16025 13787 16083 13793
rect 16025 13753 16037 13787
rect 16071 13784 16083 13787
rect 17420 13784 17448 13883
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 18782 13880 18788 13932
rect 18840 13880 18846 13932
rect 18984 13852 19012 13960
rect 19058 13948 19064 14000
rect 19116 13948 19122 14000
rect 19972 13991 20030 13997
rect 19972 13957 19984 13991
rect 20018 13988 20030 13991
rect 20438 13988 20444 14000
rect 20018 13960 20444 13988
rect 20018 13957 20030 13960
rect 19972 13951 20030 13957
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 19702 13880 19708 13932
rect 19760 13880 19766 13932
rect 21100 13920 21128 14019
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 22005 14059 22063 14065
rect 22005 14056 22017 14059
rect 21232 14028 22017 14056
rect 21232 14016 21238 14028
rect 22005 14025 22017 14028
rect 22051 14025 22063 14059
rect 22005 14019 22063 14025
rect 22278 14016 22284 14068
rect 22336 14056 22342 14068
rect 24026 14056 24032 14068
rect 22336 14028 24032 14056
rect 22336 14016 22342 14028
rect 24026 14016 24032 14028
rect 24084 14056 24090 14068
rect 24673 14059 24731 14065
rect 24673 14056 24685 14059
rect 24084 14028 24685 14056
rect 24084 14016 24090 14028
rect 24673 14025 24685 14028
rect 24719 14025 24731 14059
rect 24673 14019 24731 14025
rect 25041 14059 25099 14065
rect 25041 14025 25053 14059
rect 25087 14056 25099 14059
rect 25130 14056 25136 14068
rect 25087 14028 25136 14056
rect 25087 14025 25099 14028
rect 25041 14019 25099 14025
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 26602 14056 26608 14068
rect 25608 14028 26608 14056
rect 25608 13988 25636 14028
rect 26602 14016 26608 14028
rect 26660 14056 26666 14068
rect 27522 14056 27528 14068
rect 26660 14028 27528 14056
rect 26660 14016 26666 14028
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 28074 14056 28080 14068
rect 27908 14028 28080 14056
rect 24596 13960 25636 13988
rect 24596 13932 24624 13960
rect 27706 13948 27712 14000
rect 27764 13948 27770 14000
rect 21100 13892 22094 13920
rect 22066 13852 22094 13892
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22278 13880 22284 13932
rect 22336 13880 22342 13932
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13920 22431 13923
rect 22462 13920 22468 13932
rect 22419 13892 22468 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22572 13852 22600 13883
rect 23290 13880 23296 13932
rect 23348 13880 23354 13932
rect 24578 13880 24584 13932
rect 24636 13880 24642 13932
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 24820 13892 24869 13920
rect 24820 13880 24826 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 26786 13880 26792 13932
rect 26844 13920 26850 13932
rect 27479 13923 27537 13929
rect 27479 13920 27491 13923
rect 26844 13892 27491 13920
rect 26844 13880 26850 13892
rect 27479 13889 27491 13892
rect 27525 13889 27537 13923
rect 27479 13883 27537 13889
rect 27614 13880 27620 13932
rect 27672 13880 27678 13932
rect 27801 13929 27859 13935
rect 27801 13895 27813 13929
rect 27847 13926 27859 13929
rect 27908 13926 27936 14028
rect 28074 14016 28080 14028
rect 28132 14056 28138 14068
rect 28905 14059 28963 14065
rect 28905 14056 28917 14059
rect 28132 14028 28917 14056
rect 28132 14016 28138 14028
rect 28905 14025 28917 14028
rect 28951 14025 28963 14059
rect 28905 14019 28963 14025
rect 29089 14059 29147 14065
rect 29089 14025 29101 14059
rect 29135 14056 29147 14059
rect 29914 14056 29920 14068
rect 29135 14028 29920 14056
rect 29135 14025 29147 14028
rect 29089 14019 29147 14025
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 30098 14016 30104 14068
rect 30156 14016 30162 14068
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 31294 14056 31300 14068
rect 30892 14028 31300 14056
rect 30892 14016 30898 14028
rect 31294 14016 31300 14028
rect 31352 14016 31358 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 32582 14056 32588 14068
rect 31435 14028 32588 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 32582 14016 32588 14028
rect 32640 14056 32646 14068
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 32640 14028 33701 14056
rect 32640 14016 32646 14028
rect 33689 14025 33701 14028
rect 33735 14025 33747 14059
rect 33689 14019 33747 14025
rect 27982 13948 27988 14000
rect 28040 13988 28046 14000
rect 28721 13991 28779 13997
rect 28721 13988 28733 13991
rect 28040 13960 28733 13988
rect 28040 13948 28046 13960
rect 28721 13957 28733 13960
rect 28767 13957 28779 13991
rect 28721 13951 28779 13957
rect 29656 13960 31340 13988
rect 29656 13932 29684 13960
rect 27847 13898 27936 13926
rect 27847 13895 27859 13898
rect 27801 13889 27859 13895
rect 28166 13880 28172 13932
rect 28224 13920 28230 13932
rect 28902 13920 28908 13932
rect 28224 13892 28908 13920
rect 28224 13880 28230 13892
rect 28902 13880 28908 13892
rect 28960 13920 28966 13932
rect 28960 13892 29592 13920
rect 28960 13880 28966 13892
rect 18984 13824 19748 13852
rect 22066 13824 22600 13852
rect 16071 13756 17448 13784
rect 16071 13753 16083 13756
rect 16025 13747 16083 13753
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 4246 13716 4252 13728
rect 3016 13688 4252 13716
rect 3016 13676 3022 13688
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 6733 13719 6791 13725
rect 6733 13685 6745 13719
rect 6779 13716 6791 13719
rect 6822 13716 6828 13728
rect 6779 13688 6828 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 13446 13676 13452 13728
rect 13504 13716 13510 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13504 13688 13553 13716
rect 13504 13676 13510 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 19720 13716 19748 13824
rect 23842 13812 23848 13864
rect 23900 13852 23906 13864
rect 25774 13852 25780 13864
rect 23900 13824 25780 13852
rect 23900 13812 23906 13824
rect 25774 13812 25780 13824
rect 25832 13812 25838 13864
rect 26878 13812 26884 13864
rect 26936 13852 26942 13864
rect 27341 13855 27399 13861
rect 27341 13852 27353 13855
rect 26936 13824 27353 13852
rect 26936 13812 26942 13824
rect 27341 13821 27353 13824
rect 27387 13821 27399 13855
rect 27341 13815 27399 13821
rect 27985 13855 28043 13861
rect 27985 13821 27997 13855
rect 28031 13852 28043 13855
rect 28626 13852 28632 13864
rect 28031 13824 28632 13852
rect 28031 13821 28043 13824
rect 27985 13815 28043 13821
rect 28626 13812 28632 13824
rect 28684 13812 28690 13864
rect 29564 13852 29592 13892
rect 29638 13880 29644 13932
rect 29696 13880 29702 13932
rect 29730 13880 29736 13932
rect 29788 13880 29794 13932
rect 31312 13929 31340 13960
rect 29917 13923 29975 13929
rect 29917 13889 29929 13923
rect 29963 13889 29975 13923
rect 29917 13883 29975 13889
rect 31297 13923 31355 13929
rect 31297 13889 31309 13923
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 29748 13852 29776 13880
rect 29564 13824 29776 13852
rect 27614 13744 27620 13796
rect 27672 13784 27678 13796
rect 28166 13784 28172 13796
rect 27672 13756 28172 13784
rect 27672 13744 27678 13756
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 28350 13744 28356 13796
rect 28408 13784 28414 13796
rect 29932 13784 29960 13883
rect 30374 13784 30380 13796
rect 28408 13756 30380 13784
rect 28408 13744 28414 13756
rect 30374 13744 30380 13756
rect 30432 13744 30438 13796
rect 19886 13716 19892 13728
rect 19720 13688 19892 13716
rect 13541 13679 13599 13685
rect 19886 13676 19892 13688
rect 19944 13676 19950 13728
rect 20898 13676 20904 13728
rect 20956 13716 20962 13728
rect 23109 13719 23167 13725
rect 23109 13716 23121 13719
rect 20956 13688 23121 13716
rect 20956 13676 20962 13688
rect 23109 13685 23121 13688
rect 23155 13685 23167 13719
rect 23109 13679 23167 13685
rect 28902 13676 28908 13728
rect 28960 13676 28966 13728
rect 31312 13716 31340 13883
rect 31386 13880 31392 13932
rect 31444 13920 31450 13932
rect 31573 13923 31631 13929
rect 31573 13920 31585 13923
rect 31444 13892 31585 13920
rect 31444 13880 31450 13892
rect 31573 13889 31585 13892
rect 31619 13889 31631 13923
rect 31573 13883 31631 13889
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13920 31815 13923
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 31803 13892 32597 13920
rect 31803 13889 31815 13892
rect 31757 13883 31815 13889
rect 32585 13889 32597 13892
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 32306 13812 32312 13864
rect 32364 13812 32370 13864
rect 32766 13716 32772 13728
rect 31312 13688 32772 13716
rect 32766 13676 32772 13688
rect 32824 13676 32830 13728
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4154 13512 4160 13524
rect 3467 13484 4160 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4540 13484 5488 13512
rect 2590 13404 2596 13456
rect 2648 13444 2654 13456
rect 2648 13416 2774 13444
rect 2648 13404 2654 13416
rect 2746 13376 2774 13416
rect 4540 13376 4568 13484
rect 5258 13376 5264 13388
rect 2746 13348 4568 13376
rect 4632 13348 5264 13376
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2958 13308 2964 13320
rect 2547 13280 2964 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2332 13240 2360 13271
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3878 13308 3884 13320
rect 3283 13280 3884 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3068 13240 3096 13271
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 4632 13317 4660 13348
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5460 13376 5488 13484
rect 5534 13472 5540 13524
rect 5592 13472 5598 13524
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 10870 13512 10876 13524
rect 5684 13484 10876 13512
rect 5684 13472 5690 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 15654 13472 15660 13524
rect 15712 13472 15718 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 27028 13484 27353 13512
rect 27028 13472 27034 13484
rect 27341 13481 27353 13484
rect 27387 13481 27399 13515
rect 27341 13475 27399 13481
rect 31665 13515 31723 13521
rect 31665 13481 31677 13515
rect 31711 13512 31723 13515
rect 32306 13512 32312 13524
rect 31711 13484 32312 13512
rect 31711 13481 31723 13484
rect 31665 13475 31723 13481
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 14550 13404 14556 13456
rect 14608 13444 14614 13456
rect 17586 13444 17592 13456
rect 14608 13416 17592 13444
rect 14608 13404 14614 13416
rect 17586 13404 17592 13416
rect 17644 13444 17650 13456
rect 17644 13416 17724 13444
rect 17644 13404 17650 13416
rect 5460 13348 5580 13376
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5552 13317 5580 13348
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 9030 13376 9036 13388
rect 8536 13348 9036 13376
rect 8536 13336 8542 13348
rect 9030 13336 9036 13348
rect 9088 13376 9094 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9088 13348 9413 13376
rect 9088 13336 9094 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 15378 13376 15384 13388
rect 9401 13339 9459 13345
rect 10888 13348 15384 13376
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5132 13280 5365 13308
rect 5132 13268 5138 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 8294 13308 8300 13320
rect 5583 13280 8300 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 3970 13240 3976 13252
rect 2332 13212 3976 13240
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4249 13243 4307 13249
rect 4249 13209 4261 13243
rect 4295 13240 4307 13243
rect 8404 13240 8432 13271
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 4295 13212 8432 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 2406 13132 2412 13184
rect 2464 13132 2470 13184
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 4264 13172 4292 13203
rect 8570 13200 8576 13252
rect 8628 13200 8634 13252
rect 9858 13200 9864 13252
rect 9916 13200 9922 13252
rect 3292 13144 4292 13172
rect 3292 13132 3298 13144
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 10888 13181 10916 13348
rect 15378 13336 15384 13348
rect 15436 13376 15442 13388
rect 16761 13379 16819 13385
rect 15436 13348 15516 13376
rect 15436 13336 15442 13348
rect 11790 13268 11796 13320
rect 11848 13268 11854 13320
rect 15488 13317 15516 13348
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 16850 13376 16856 13388
rect 16807 13348 16856 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14752 13280 15025 13308
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 14090 13240 14096 13252
rect 13294 13212 14096 13240
rect 14090 13200 14096 13212
rect 14148 13200 14154 13252
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 8996 13144 10885 13172
rect 8996 13132 9002 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13136 13144 13553 13172
rect 13136 13132 13142 13144
rect 13541 13141 13553 13144
rect 13587 13172 13599 13175
rect 14752 13172 14780 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 15746 13308 15752 13320
rect 15519 13280 15752 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 17696 13317 17724 13416
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 22830 13376 22836 13388
rect 19668 13348 22836 13376
rect 19668 13336 19674 13348
rect 22830 13336 22836 13348
rect 22888 13376 22894 13388
rect 28074 13376 28080 13388
rect 22888 13348 28080 13376
rect 22888 13336 22894 13348
rect 28074 13336 28080 13348
rect 28132 13336 28138 13388
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18322 13308 18328 13320
rect 18279 13280 18328 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 19852 13280 20269 13308
rect 19852 13268 19858 13280
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 26050 13268 26056 13320
rect 26108 13268 26114 13320
rect 32950 13268 32956 13320
rect 33008 13268 33014 13320
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15620 13212 16221 13240
rect 15620 13200 15626 13212
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 18417 13243 18475 13249
rect 18417 13209 18429 13243
rect 18463 13240 18475 13243
rect 20346 13240 20352 13252
rect 18463 13212 20352 13240
rect 18463 13209 18475 13212
rect 18417 13203 18475 13209
rect 20346 13200 20352 13212
rect 20404 13200 20410 13252
rect 15930 13172 15936 13184
rect 13587 13144 15936 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 18230 13132 18236 13184
rect 18288 13172 18294 13184
rect 21545 13175 21603 13181
rect 21545 13172 21557 13175
rect 18288 13144 21557 13172
rect 18288 13132 18294 13144
rect 21545 13141 21557 13144
rect 21591 13141 21603 13175
rect 21545 13135 21603 13141
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 2590 12928 2596 12980
rect 2648 12928 2654 12980
rect 3878 12928 3884 12980
rect 3936 12928 3942 12980
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 4028 12940 4353 12968
rect 4028 12928 4034 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 9122 12928 9128 12980
rect 9180 12928 9186 12980
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17552 12940 19564 12968
rect 17552 12928 17558 12940
rect 2608 12900 2636 12928
rect 2148 12872 2636 12900
rect 2148 12841 2176 12872
rect 3050 12860 3056 12912
rect 3108 12860 3114 12912
rect 8570 12860 8576 12912
rect 8628 12860 8634 12912
rect 9140 12900 9168 12928
rect 11790 12900 11796 12912
rect 9140 12872 11796 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4120 12804 4353 12832
rect 4120 12792 4126 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4522 12792 4528 12844
rect 4580 12792 4586 12844
rect 9600 12841 9628 12872
rect 11790 12860 11796 12872
rect 11848 12860 11854 12912
rect 12986 12860 12992 12912
rect 13044 12860 13050 12912
rect 14734 12860 14740 12912
rect 14792 12860 14798 12912
rect 18414 12900 18420 12912
rect 18064 12872 18420 12900
rect 18064 12844 18092 12872
rect 18414 12860 18420 12872
rect 18472 12900 18478 12912
rect 19153 12903 19211 12909
rect 18472 12872 19012 12900
rect 18472 12860 18478 12872
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15252 12804 15393 12832
rect 15252 12792 15258 12804
rect 15381 12801 15393 12804
rect 15427 12832 15439 12835
rect 15562 12832 15568 12844
rect 15427 12804 15568 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16390 12832 16396 12844
rect 16071 12804 16396 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 2406 12724 2412 12776
rect 2464 12724 2470 12776
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 8846 12764 8852 12776
rect 5868 12736 8852 12764
rect 5868 12724 5874 12736
rect 8846 12724 8852 12736
rect 8904 12764 8910 12776
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 8904 12736 9321 12764
rect 8904 12724 8910 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 16040 12764 16068 12795
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17586 12832 17592 12844
rect 17052 12804 17592 12832
rect 9309 12727 9367 12733
rect 14384 12736 16068 12764
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 12986 12696 12992 12708
rect 10928 12668 12992 12696
rect 10928 12656 10934 12668
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 14384 12640 14412 12736
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 17052 12764 17080 12804
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18984 12841 19012 12872
rect 19153 12869 19165 12903
rect 19199 12900 19211 12903
rect 19426 12900 19432 12912
rect 19199 12872 19432 12900
rect 19199 12869 19211 12872
rect 19153 12863 19211 12869
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 19536 12900 19564 12940
rect 19886 12928 19892 12980
rect 19944 12968 19950 12980
rect 19944 12940 22600 12968
rect 19944 12928 19950 12940
rect 22572 12909 22600 12940
rect 22922 12928 22928 12980
rect 22980 12928 22986 12980
rect 27798 12968 27804 12980
rect 27448 12940 27804 12968
rect 22557 12903 22615 12909
rect 19536 12872 22416 12900
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18156 12804 18797 12832
rect 16172 12736 17080 12764
rect 16172 12724 16178 12736
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 18156 12764 18184 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 19961 12835 20019 12841
rect 19961 12832 19973 12835
rect 19852 12804 19973 12832
rect 19852 12792 19858 12804
rect 19961 12801 19973 12804
rect 20007 12801 20019 12835
rect 19961 12795 20019 12801
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20404 12804 22094 12832
rect 20404 12792 20410 12804
rect 17276 12736 18184 12764
rect 18325 12767 18383 12773
rect 17276 12724 17282 12736
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 19610 12764 19616 12776
rect 18371 12736 19616 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7616 12600 7849 12628
rect 7616 12588 7622 12600
rect 7837 12597 7849 12600
rect 7883 12628 7895 12631
rect 14366 12628 14372 12640
rect 7883 12600 14372 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 19720 12628 19748 12727
rect 22066 12696 22094 12804
rect 22278 12792 22284 12844
rect 22336 12792 22342 12844
rect 22388 12841 22416 12872
rect 22557 12869 22569 12903
rect 22603 12869 22615 12903
rect 22557 12863 22615 12869
rect 22649 12903 22707 12909
rect 22649 12869 22661 12903
rect 22695 12900 22707 12903
rect 24762 12900 24768 12912
rect 22695 12872 24768 12900
rect 22695 12869 22707 12872
rect 22649 12863 22707 12869
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 22374 12835 22432 12841
rect 22374 12801 22386 12835
rect 22420 12801 22432 12835
rect 22374 12795 22432 12801
rect 22746 12835 22804 12841
rect 22746 12801 22758 12835
rect 22792 12801 22804 12835
rect 22746 12795 22804 12801
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 22756 12764 22784 12795
rect 26694 12792 26700 12844
rect 26752 12832 26758 12844
rect 27448 12841 27476 12940
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 27893 12971 27951 12977
rect 27893 12937 27905 12971
rect 27939 12968 27951 12971
rect 28442 12968 28448 12980
rect 27939 12940 28448 12968
rect 27939 12937 27951 12940
rect 27893 12931 27951 12937
rect 28442 12928 28448 12940
rect 28500 12928 28506 12980
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 32309 12971 32367 12977
rect 32309 12968 32321 12971
rect 32180 12940 32321 12968
rect 32180 12928 32186 12940
rect 32309 12937 32321 12940
rect 32355 12937 32367 12971
rect 32309 12931 32367 12937
rect 32677 12971 32735 12977
rect 32677 12937 32689 12971
rect 32723 12968 32735 12971
rect 33226 12968 33232 12980
rect 32723 12940 33232 12968
rect 32723 12937 32735 12940
rect 32677 12931 32735 12937
rect 33226 12928 33232 12940
rect 33284 12928 33290 12980
rect 27617 12903 27675 12909
rect 27617 12869 27629 12903
rect 27663 12900 27675 12903
rect 27982 12900 27988 12912
rect 27663 12872 27988 12900
rect 27663 12869 27675 12872
rect 27617 12863 27675 12869
rect 27982 12860 27988 12872
rect 28040 12860 28046 12912
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 26752 12804 27261 12832
rect 26752 12792 26758 12804
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27397 12835 27476 12841
rect 27397 12801 27409 12835
rect 27443 12804 27476 12835
rect 27525 12835 27583 12841
rect 27443 12801 27455 12804
rect 27397 12795 27455 12801
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27714 12835 27772 12841
rect 27714 12832 27726 12835
rect 27525 12795 27583 12801
rect 27632 12804 27726 12832
rect 22520 12736 22784 12764
rect 22520 12724 22526 12736
rect 23750 12724 23756 12776
rect 23808 12764 23814 12776
rect 27540 12764 27568 12795
rect 23808 12736 27568 12764
rect 23808 12724 23814 12736
rect 27632 12696 27660 12804
rect 27714 12801 27726 12804
rect 27760 12801 27772 12835
rect 27714 12795 27772 12801
rect 28350 12792 28356 12844
rect 28408 12832 28414 12844
rect 28537 12835 28595 12841
rect 28537 12832 28549 12835
rect 28408 12804 28549 12832
rect 28408 12792 28414 12804
rect 28537 12801 28549 12804
rect 28583 12801 28595 12835
rect 28537 12795 28595 12801
rect 28718 12792 28724 12844
rect 28776 12792 28782 12844
rect 28813 12835 28871 12841
rect 28813 12801 28825 12835
rect 28859 12801 28871 12835
rect 28813 12795 28871 12801
rect 28828 12764 28856 12795
rect 29638 12792 29644 12844
rect 29696 12832 29702 12844
rect 29733 12835 29791 12841
rect 29733 12832 29745 12835
rect 29696 12804 29745 12832
rect 29696 12792 29702 12804
rect 29733 12801 29745 12804
rect 29779 12801 29791 12835
rect 29733 12795 29791 12801
rect 31938 12792 31944 12844
rect 31996 12832 32002 12844
rect 32493 12835 32551 12841
rect 32493 12832 32505 12835
rect 31996 12804 32505 12832
rect 31996 12792 32002 12804
rect 32493 12801 32505 12804
rect 32539 12801 32551 12835
rect 32493 12795 32551 12801
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 32858 12832 32864 12844
rect 32815 12804 32864 12832
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 32858 12792 32864 12804
rect 32916 12792 32922 12844
rect 29549 12767 29607 12773
rect 29549 12764 29561 12767
rect 28828 12736 29561 12764
rect 29549 12733 29561 12736
rect 29595 12764 29607 12767
rect 30190 12764 30196 12776
rect 29595 12736 30196 12764
rect 29595 12733 29607 12736
rect 29549 12727 29607 12733
rect 30190 12724 30196 12736
rect 30248 12724 30254 12776
rect 27706 12696 27712 12708
rect 22066 12668 27712 12696
rect 27706 12656 27712 12668
rect 27764 12656 27770 12708
rect 28902 12696 28908 12708
rect 27816 12668 28908 12696
rect 19978 12628 19984 12640
rect 19720 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 21082 12588 21088 12640
rect 21140 12588 21146 12640
rect 25774 12588 25780 12640
rect 25832 12628 25838 12640
rect 27816 12628 27844 12668
rect 28902 12656 28908 12668
rect 28960 12656 28966 12708
rect 25832 12600 27844 12628
rect 25832 12588 25838 12600
rect 28350 12588 28356 12640
rect 28408 12588 28414 12640
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 3050 12384 3056 12436
rect 3108 12384 3114 12436
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19852 12396 19901 12424
rect 19852 12384 19858 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 19889 12387 19947 12393
rect 21910 12384 21916 12436
rect 21968 12424 21974 12436
rect 22097 12427 22155 12433
rect 22097 12424 22109 12427
rect 21968 12396 22109 12424
rect 21968 12384 21974 12396
rect 22097 12393 22109 12396
rect 22143 12424 22155 12427
rect 22554 12424 22560 12436
rect 22143 12396 22560 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 22554 12384 22560 12396
rect 22612 12424 22618 12436
rect 22612 12396 24624 12424
rect 22612 12384 22618 12396
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 15988 12328 16620 12356
rect 15988 12316 15994 12328
rect 3050 12180 3056 12232
rect 3108 12180 3114 12232
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14424 12192 14565 12220
rect 14424 12180 14430 12192
rect 14553 12189 14565 12192
rect 14599 12220 14611 12223
rect 14734 12220 14740 12232
rect 14599 12192 14740 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15804 12192 15945 12220
rect 15804 12180 15810 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 16592 12220 16620 12328
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19702 12356 19708 12368
rect 19392 12328 19708 12356
rect 19392 12316 19398 12328
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 21818 12316 21824 12368
rect 21876 12356 21882 12368
rect 23017 12359 23075 12365
rect 23017 12356 23029 12359
rect 21876 12328 23029 12356
rect 21876 12316 21882 12328
rect 23017 12325 23029 12328
rect 23063 12325 23075 12359
rect 24596 12356 24624 12396
rect 24670 12384 24676 12436
rect 24728 12424 24734 12436
rect 28534 12424 28540 12436
rect 24728 12396 28540 12424
rect 24728 12384 24734 12396
rect 28534 12384 28540 12396
rect 28592 12384 28598 12436
rect 25682 12356 25688 12368
rect 24596 12328 25688 12356
rect 23017 12319 23075 12325
rect 25682 12316 25688 12328
rect 25740 12356 25746 12368
rect 27890 12356 27896 12368
rect 25740 12328 27896 12356
rect 25740 12316 25746 12328
rect 27890 12316 27896 12328
rect 27948 12316 27954 12368
rect 27985 12359 28043 12365
rect 27985 12325 27997 12359
rect 28031 12325 28043 12359
rect 27985 12319 28043 12325
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 18046 12288 18052 12300
rect 16715 12260 18052 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16592 12192 16773 12220
rect 15933 12183 15991 12189
rect 16761 12189 16773 12192
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17494 12220 17500 12232
rect 16908 12192 17500 12220
rect 16908 12180 16914 12192
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17972 12229 18000 12260
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 21082 12288 21088 12300
rect 19536 12260 21088 12288
rect 19536 12229 19564 12260
rect 21082 12248 21088 12260
rect 21140 12288 21146 12300
rect 28000 12288 28028 12319
rect 28718 12288 28724 12300
rect 21140 12260 23336 12288
rect 21140 12248 21146 12260
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 15013 12155 15071 12161
rect 15013 12121 15025 12155
rect 15059 12152 15071 12155
rect 16574 12152 16580 12164
rect 15059 12124 16580 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 16574 12112 16580 12124
rect 16632 12152 16638 12164
rect 17218 12152 17224 12164
rect 16632 12124 17224 12152
rect 16632 12112 16638 12124
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 18233 12155 18291 12161
rect 18233 12121 18245 12155
rect 18279 12152 18291 12155
rect 18690 12152 18696 12164
rect 18279 12124 18696 12152
rect 18279 12121 18291 12124
rect 18233 12115 18291 12121
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 19444 12152 19472 12183
rect 19702 12180 19708 12232
rect 19760 12180 19766 12232
rect 20898 12220 20904 12232
rect 19812 12192 20904 12220
rect 19812 12152 19840 12192
rect 20898 12180 20904 12192
rect 20956 12220 20962 12232
rect 21542 12220 21548 12232
rect 20956 12192 21548 12220
rect 20956 12180 20962 12192
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 23308 12229 23336 12260
rect 23492 12260 28028 12288
rect 28552 12260 28724 12288
rect 23492 12229 23520 12260
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 22796 12192 23213 12220
rect 22796 12180 22802 12192
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23293 12223 23351 12229
rect 23293 12189 23305 12223
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 19444 12124 19840 12152
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 20809 12155 20867 12161
rect 20809 12152 20821 12155
rect 20588 12124 20821 12152
rect 20588 12112 20594 12124
rect 20809 12121 20821 12124
rect 20855 12121 20867 12155
rect 23584 12152 23612 12183
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 28166 12229 28172 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24728 12192 24777 12220
rect 24728 12180 24734 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12189 25099 12223
rect 28164 12220 28172 12229
rect 28127 12192 28172 12220
rect 25041 12183 25099 12189
rect 28164 12183 28172 12192
rect 20809 12115 20867 12121
rect 20916 12124 22094 12152
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 20916 12084 20944 12124
rect 20680 12056 20944 12084
rect 22066 12084 22094 12124
rect 22664 12124 23612 12152
rect 22664 12084 22692 12124
rect 24026 12112 24032 12164
rect 24084 12152 24090 12164
rect 24596 12152 24624 12180
rect 25056 12152 25084 12183
rect 28166 12180 28172 12183
rect 28224 12180 28230 12232
rect 28552 12229 28580 12260
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 28536 12223 28594 12229
rect 28536 12189 28548 12223
rect 28582 12189 28594 12223
rect 28536 12183 28594 12189
rect 28626 12180 28632 12232
rect 28684 12180 28690 12232
rect 24084 12124 25084 12152
rect 28261 12155 28319 12161
rect 24084 12112 24090 12124
rect 28261 12121 28273 12155
rect 28307 12121 28319 12155
rect 28261 12115 28319 12121
rect 28353 12155 28411 12161
rect 28353 12121 28365 12155
rect 28399 12152 28411 12155
rect 28442 12152 28448 12164
rect 28399 12124 28448 12152
rect 28399 12121 28411 12124
rect 28353 12115 28411 12121
rect 22066 12056 22692 12084
rect 20680 12044 20686 12056
rect 24578 12044 24584 12096
rect 24636 12044 24642 12096
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 24949 12087 25007 12093
rect 24949 12084 24961 12087
rect 24820 12056 24961 12084
rect 24820 12044 24826 12056
rect 24949 12053 24961 12056
rect 24995 12053 25007 12087
rect 28276 12084 28304 12115
rect 28442 12112 28448 12124
rect 28500 12112 28506 12164
rect 30374 12112 30380 12164
rect 30432 12152 30438 12164
rect 31386 12152 31392 12164
rect 30432 12124 31392 12152
rect 30432 12112 30438 12124
rect 31386 12112 31392 12124
rect 31444 12112 31450 12164
rect 31202 12084 31208 12096
rect 28276 12056 31208 12084
rect 24949 12047 25007 12053
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 22370 11840 22376 11892
rect 22428 11840 22434 11892
rect 22664 11852 24716 11880
rect 15194 11812 15200 11824
rect 14200 11784 15200 11812
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 14200 11753 14228 11784
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 15746 11772 15752 11824
rect 15804 11772 15810 11824
rect 16301 11815 16359 11821
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 22664 11812 22692 11852
rect 16347 11784 18092 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13504 11716 14197 11744
rect 13504 11704 13510 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14550 11704 14556 11756
rect 14608 11704 14614 11756
rect 14734 11704 14740 11756
rect 14792 11704 14798 11756
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 18064 11753 18092 11784
rect 19812 11784 22692 11812
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11744 18107 11747
rect 18322 11744 18328 11756
rect 18095 11716 18328 11744
rect 18095 11713 18107 11716
rect 18049 11707 18107 11713
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 19812 11688 19840 11784
rect 20340 11747 20398 11753
rect 20340 11713 20352 11747
rect 20386 11744 20398 11747
rect 20898 11744 20904 11756
rect 20386 11716 20904 11744
rect 20386 11713 20398 11716
rect 20340 11707 20398 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 22572 11753 22600 11784
rect 22738 11772 22744 11824
rect 22796 11772 22802 11824
rect 23474 11812 23480 11824
rect 22848 11784 23480 11812
rect 22557 11747 22615 11753
rect 22557 11713 22569 11747
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11744 22707 11747
rect 22848 11744 22876 11784
rect 23474 11772 23480 11784
rect 23532 11772 23538 11824
rect 24112 11815 24170 11821
rect 24112 11781 24124 11815
rect 24158 11812 24170 11815
rect 24578 11812 24584 11824
rect 24158 11784 24584 11812
rect 24158 11781 24170 11784
rect 24112 11775 24170 11781
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 24688 11812 24716 11852
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 25225 11883 25283 11889
rect 25225 11880 25237 11883
rect 24820 11852 25237 11880
rect 24820 11840 24826 11852
rect 25225 11849 25237 11852
rect 25271 11849 25283 11883
rect 25225 11843 25283 11849
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 25869 11883 25927 11889
rect 25869 11880 25881 11883
rect 25372 11852 25881 11880
rect 25372 11840 25378 11852
rect 25869 11849 25881 11852
rect 25915 11880 25927 11883
rect 28442 11880 28448 11892
rect 25915 11852 28448 11880
rect 25915 11849 25927 11852
rect 25869 11843 25927 11849
rect 28442 11840 28448 11852
rect 28500 11840 28506 11892
rect 28718 11840 28724 11892
rect 28776 11840 28782 11892
rect 31202 11840 31208 11892
rect 31260 11840 31266 11892
rect 32674 11840 32680 11892
rect 32732 11880 32738 11892
rect 33686 11880 33692 11892
rect 32732 11852 33692 11880
rect 32732 11840 32738 11852
rect 33686 11840 33692 11852
rect 33744 11840 33750 11892
rect 25130 11812 25136 11824
rect 24688 11784 25136 11812
rect 25130 11772 25136 11784
rect 25188 11772 25194 11824
rect 25682 11772 25688 11824
rect 25740 11772 25746 11824
rect 27608 11815 27666 11821
rect 27608 11781 27620 11815
rect 27654 11812 27666 11815
rect 28350 11812 28356 11824
rect 27654 11784 28356 11812
rect 27654 11781 27666 11784
rect 27608 11775 27666 11781
rect 28350 11772 28356 11784
rect 28408 11772 28414 11824
rect 31312 11784 32812 11812
rect 22695 11716 22876 11744
rect 22925 11747 22983 11753
rect 22695 11713 22707 11716
rect 22649 11707 22707 11713
rect 22925 11713 22937 11747
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 19794 11676 19800 11688
rect 18279 11648 19800 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 20036 11648 20085 11676
rect 20036 11636 20042 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 22940 11676 22968 11707
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 27890 11744 27896 11756
rect 23716 11716 27896 11744
rect 23716 11704 23722 11716
rect 27890 11704 27896 11716
rect 27948 11704 27954 11756
rect 30190 11704 30196 11756
rect 30248 11744 30254 11756
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 30248 11716 31125 11744
rect 30248 11704 30254 11716
rect 31113 11713 31125 11716
rect 31159 11744 31171 11747
rect 31312 11744 31340 11784
rect 31159 11716 31340 11744
rect 31159 11713 31171 11716
rect 31113 11707 31171 11713
rect 31386 11704 31392 11756
rect 31444 11704 31450 11756
rect 32784 11753 32812 11784
rect 32493 11747 32551 11753
rect 32493 11713 32505 11747
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11744 32827 11747
rect 33410 11744 33416 11756
rect 32815 11716 33416 11744
rect 32815 11713 32827 11716
rect 32769 11707 32827 11713
rect 20073 11639 20131 11645
rect 22066 11648 22968 11676
rect 21358 11568 21364 11620
rect 21416 11608 21422 11620
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 21416 11580 21465 11608
rect 21416 11568 21422 11580
rect 21453 11577 21465 11580
rect 21499 11608 21511 11611
rect 22066 11608 22094 11648
rect 23842 11636 23848 11688
rect 23900 11636 23906 11688
rect 27338 11636 27344 11688
rect 27396 11636 27402 11688
rect 28534 11636 28540 11688
rect 28592 11676 28598 11688
rect 32508 11676 32536 11707
rect 33410 11704 33416 11716
rect 33468 11704 33474 11756
rect 28592 11648 32536 11676
rect 28592 11636 28598 11648
rect 21499 11580 22094 11608
rect 31573 11611 31631 11617
rect 21499 11577 21511 11580
rect 21453 11571 21511 11577
rect 31573 11577 31585 11611
rect 31619 11608 31631 11611
rect 32490 11608 32496 11620
rect 31619 11580 32496 11608
rect 31619 11577 31631 11580
rect 31573 11571 31631 11577
rect 32490 11568 32496 11580
rect 32548 11568 32554 11620
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 22462 11540 22468 11552
rect 17920 11512 22468 11540
rect 17920 11500 17926 11512
rect 22462 11500 22468 11512
rect 22520 11540 22526 11552
rect 25314 11540 25320 11552
rect 22520 11512 25320 11540
rect 22520 11500 22526 11512
rect 25314 11500 25320 11512
rect 25372 11500 25378 11552
rect 25774 11500 25780 11552
rect 25832 11540 25838 11552
rect 25869 11543 25927 11549
rect 25869 11540 25881 11543
rect 25832 11512 25881 11540
rect 25832 11500 25838 11512
rect 25869 11509 25881 11512
rect 25915 11509 25927 11543
rect 25869 11503 25927 11509
rect 26050 11500 26056 11552
rect 26108 11500 26114 11552
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 32398 11540 32404 11552
rect 32355 11512 32404 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 32398 11500 32404 11512
rect 32456 11500 32462 11552
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 4522 11336 4528 11348
rect 4203 11308 4528 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 20533 11339 20591 11345
rect 20533 11305 20545 11339
rect 20579 11336 20591 11339
rect 20622 11336 20628 11348
rect 20579 11308 20628 11336
rect 20579 11305 20591 11308
rect 20533 11299 20591 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20956 11308 21005 11336
rect 20956 11296 20962 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 26786 11336 26792 11348
rect 21140 11308 26792 11336
rect 21140 11296 21146 11308
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 31202 11296 31208 11348
rect 31260 11336 31266 11348
rect 31389 11339 31447 11345
rect 31389 11336 31401 11339
rect 31260 11308 31401 11336
rect 31260 11296 31266 11308
rect 31389 11305 31401 11308
rect 31435 11305 31447 11339
rect 31389 11299 31447 11305
rect 17862 11228 17868 11280
rect 17920 11228 17926 11280
rect 19886 11228 19892 11280
rect 19944 11228 19950 11280
rect 23658 11268 23664 11280
rect 20272 11240 23664 11268
rect 12348 11212 12400 11218
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 19904 11200 19932 11228
rect 17092 11172 18460 11200
rect 19904 11172 20208 11200
rect 17092 11160 17098 11172
rect 12348 11154 12400 11160
rect 5074 11092 5080 11144
rect 5132 11132 5138 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5132 11104 5549 11132
rect 5132 11092 5138 11104
rect 5537 11101 5549 11104
rect 5583 11132 5595 11135
rect 7190 11132 7196 11144
rect 5583 11104 7196 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 7190 11092 7196 11104
rect 7248 11132 7254 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 7248 11104 10333 11132
rect 7248 11092 7254 11104
rect 10321 11101 10333 11104
rect 10367 11132 10379 11135
rect 11054 11132 11060 11144
rect 10367 11104 11060 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11974 11132 11980 11144
rect 11164 11104 11980 11132
rect 11164 11076 11192 11104
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12584 11104 12725 11132
rect 12584 11092 12590 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 12894 11132 12900 11144
rect 12759 11104 12900 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11092 13084 11144
rect 13136 11092 13142 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13463 11135 13521 11141
rect 13463 11132 13475 11135
rect 13320 11104 13475 11132
rect 13320 11092 13326 11104
rect 13463 11101 13475 11104
rect 13509 11101 13521 11135
rect 13463 11095 13521 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17218 11132 17224 11144
rect 17175 11104 17224 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 3970 11024 3976 11076
rect 4028 11024 4034 11076
rect 4246 11073 4252 11076
rect 4189 11067 4252 11073
rect 4189 11033 4201 11067
rect 4235 11033 4252 11067
rect 4189 11027 4252 11033
rect 4246 11024 4252 11027
rect 4304 11024 4310 11076
rect 5810 11073 5816 11076
rect 5804 11064 5816 11073
rect 5771 11036 5816 11064
rect 5804 11027 5816 11036
rect 5810 11024 5816 11027
rect 5868 11024 5874 11076
rect 10588 11067 10646 11073
rect 10588 11033 10600 11067
rect 10634 11064 10646 11067
rect 11146 11064 11152 11076
rect 10634 11036 11152 11064
rect 10634 11033 10646 11036
rect 10588 11027 10646 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 12434 11064 12440 11076
rect 11716 11036 12440 11064
rect 4338 10956 4344 11008
rect 4396 10956 4402 11008
rect 6914 10956 6920 11008
rect 6972 10956 6978 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 7834 10996 7840 11008
rect 7340 10968 7840 10996
rect 7340 10956 7346 10968
rect 7834 10956 7840 10968
rect 7892 10996 7898 11008
rect 9214 10996 9220 11008
rect 7892 10968 9220 10996
rect 7892 10956 7898 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 11716 11005 11744 11036
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 12618 11024 12624 11076
rect 12676 11024 12682 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13228 11036 13676 11064
rect 13228 11024 13234 11036
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 12345 10999 12403 11005
rect 12345 10965 12357 10999
rect 12391 10996 12403 10999
rect 12802 10996 12808 11008
rect 12391 10968 12808 10996
rect 12391 10965 12403 10968
rect 12345 10959 12403 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 12986 10956 12992 11008
rect 13044 10996 13050 11008
rect 13262 10996 13268 11008
rect 13044 10968 13268 10996
rect 13044 10956 13050 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 13648 11005 13676 11036
rect 16666 11024 16672 11076
rect 16724 11064 16730 11076
rect 16761 11067 16819 11073
rect 16761 11064 16773 11067
rect 16724 11036 16773 11064
rect 16724 11024 16730 11036
rect 16761 11033 16773 11036
rect 16807 11033 16819 11067
rect 16960 11064 16988 11095
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17586 11092 17592 11144
rect 17644 11092 17650 11144
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11132 17923 11135
rect 18322 11132 18328 11144
rect 17911 11104 18328 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 17880 11064 17908 11095
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 16960 11036 17908 11064
rect 18432 11064 18460 11172
rect 19886 11092 19892 11144
rect 19944 11092 19950 11144
rect 20180 11141 20208 11172
rect 20272 11141 20300 11240
rect 23658 11228 23664 11240
rect 23716 11228 23722 11280
rect 24670 11268 24676 11280
rect 23860 11240 24676 11268
rect 21910 11200 21916 11212
rect 21192 11172 21916 11200
rect 19982 11135 20040 11141
rect 19982 11101 19994 11135
rect 20028 11101 20040 11135
rect 19982 11095 20040 11101
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20257 11135 20315 11141
rect 20257 11101 20269 11135
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 19996 11064 20024 11095
rect 20346 11092 20352 11144
rect 20404 11141 20410 11144
rect 20404 11132 20412 11141
rect 20404 11104 20449 11132
rect 20404 11095 20412 11104
rect 20404 11092 20410 11095
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21192 11141 21220 11172
rect 21910 11160 21916 11172
rect 21968 11200 21974 11212
rect 23860 11200 23888 11240
rect 24670 11228 24676 11240
rect 24728 11228 24734 11280
rect 25958 11200 25964 11212
rect 21968 11172 23888 11200
rect 23952 11172 25964 11200
rect 21968 11160 21974 11172
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 20772 11104 21189 11132
rect 20772 11092 20778 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21358 11092 21364 11144
rect 21416 11092 21422 11144
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11132 21511 11135
rect 21542 11132 21548 11144
rect 21499 11104 21548 11132
rect 21499 11101 21511 11104
rect 21453 11095 21511 11101
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 23750 11092 23756 11144
rect 23808 11092 23814 11144
rect 23952 11141 23980 11172
rect 25958 11160 25964 11172
rect 26016 11160 26022 11212
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24026 11092 24032 11144
rect 24084 11092 24090 11144
rect 26050 11092 26056 11144
rect 26108 11092 26114 11144
rect 29546 11092 29552 11144
rect 29604 11132 29610 11144
rect 29822 11132 29828 11144
rect 29604 11104 29828 11132
rect 29604 11092 29610 11104
rect 29822 11092 29828 11104
rect 29880 11132 29886 11144
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 29880 11104 29929 11132
rect 29880 11092 29886 11104
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 29917 11095 29975 11101
rect 30190 11092 30196 11144
rect 30248 11092 30254 11144
rect 32769 11135 32827 11141
rect 32769 11132 32781 11135
rect 32324 11104 32781 11132
rect 32324 11076 32352 11104
rect 32769 11101 32781 11104
rect 32815 11101 32827 11135
rect 32769 11095 32827 11101
rect 18432 11036 20024 11064
rect 23569 11067 23627 11073
rect 16761 11027 16819 11033
rect 23569 11033 23581 11067
rect 23615 11064 23627 11067
rect 24854 11064 24860 11076
rect 23615 11036 24860 11064
rect 23615 11033 23627 11036
rect 23569 11027 23627 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 32306 11024 32312 11076
rect 32364 11024 32370 11076
rect 32490 11024 32496 11076
rect 32548 11073 32554 11076
rect 32548 11064 32560 11073
rect 32548 11036 32593 11064
rect 32548 11027 32560 11036
rect 32548 11024 32554 11027
rect 13633 10999 13691 11005
rect 13633 10965 13645 10999
rect 13679 10965 13691 10999
rect 13633 10959 13691 10965
rect 26602 10956 26608 11008
rect 26660 10996 26666 11008
rect 27341 10999 27399 11005
rect 27341 10996 27353 10999
rect 26660 10968 27353 10996
rect 26660 10956 26666 10968
rect 27341 10965 27353 10968
rect 27387 10965 27399 10999
rect 27341 10959 27399 10965
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 29733 10999 29791 11005
rect 29733 10996 29745 10999
rect 29052 10968 29745 10996
rect 29052 10956 29058 10968
rect 29733 10965 29745 10968
rect 29779 10965 29791 10999
rect 29733 10959 29791 10965
rect 30098 10956 30104 11008
rect 30156 10956 30162 11008
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7929 10795 7987 10801
rect 6696 10764 7880 10792
rect 6696 10752 6702 10764
rect 3326 10684 3332 10736
rect 3384 10724 3390 10736
rect 3384 10696 4200 10724
rect 3384 10684 3390 10696
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 2832 10628 3249 10656
rect 2832 10616 2838 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4172 10665 4200 10696
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6788 10696 6837 10724
rect 6788 10684 6794 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7101 10727 7159 10733
rect 7101 10724 7113 10727
rect 6972 10696 7113 10724
rect 6972 10684 6978 10696
rect 7101 10693 7113 10696
rect 7147 10693 7159 10727
rect 7101 10687 7159 10693
rect 7193 10727 7251 10733
rect 7193 10693 7205 10727
rect 7239 10724 7251 10727
rect 7282 10724 7288 10736
rect 7239 10696 7288 10724
rect 7239 10693 7251 10696
rect 7193 10687 7251 10693
rect 7282 10684 7288 10696
rect 7340 10684 7346 10736
rect 7558 10684 7564 10736
rect 7616 10684 7622 10736
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3844 10628 3985 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4246 10656 4252 10668
rect 4203 10628 4252 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 7852 10656 7880 10764
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8202 10792 8208 10804
rect 7975 10764 8208 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9953 10795 10011 10801
rect 8996 10764 9628 10792
rect 8996 10752 9002 10764
rect 8846 10684 8852 10736
rect 8904 10684 8910 10736
rect 9490 10724 9496 10736
rect 8956 10696 9496 10724
rect 8956 10656 8984 10696
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 9600 10733 9628 10764
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10318 10792 10324 10804
rect 9999 10764 10324 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 10612 10764 12664 10792
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10693 9643 10727
rect 10612 10724 10640 10764
rect 9585 10687 9643 10693
rect 9784 10696 10640 10724
rect 7852 10628 8984 10656
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 9784 10656 9812 10696
rect 12526 10684 12532 10736
rect 12584 10684 12590 10736
rect 12636 10724 12664 10764
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 12768 10764 13645 10792
rect 12768 10752 12774 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 25958 10752 25964 10804
rect 26016 10752 26022 10804
rect 28721 10795 28779 10801
rect 28721 10761 28733 10795
rect 28767 10792 28779 10795
rect 29086 10792 29092 10804
rect 28767 10764 29092 10792
rect 28767 10761 28779 10764
rect 28721 10755 28779 10761
rect 29086 10752 29092 10764
rect 29144 10792 29150 10804
rect 30098 10792 30104 10804
rect 29144 10764 30104 10792
rect 29144 10752 29150 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 33686 10752 33692 10804
rect 33744 10752 33750 10804
rect 12894 10724 12900 10736
rect 12636 10696 12900 10724
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 13265 10727 13323 10733
rect 13265 10693 13277 10727
rect 13311 10724 13323 10727
rect 13446 10724 13452 10736
rect 13311 10696 13452 10724
rect 13311 10693 13323 10696
rect 13265 10687 13323 10693
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 18230 10684 18236 10736
rect 18288 10684 18294 10736
rect 19978 10684 19984 10736
rect 20036 10684 20042 10736
rect 24854 10733 24860 10736
rect 24848 10724 24860 10733
rect 24815 10696 24860 10724
rect 24848 10687 24860 10696
rect 24854 10684 24860 10687
rect 24912 10684 24918 10736
rect 27608 10727 27666 10733
rect 27608 10693 27620 10727
rect 27654 10724 27666 10727
rect 28994 10724 29000 10736
rect 27654 10696 29000 10724
rect 27654 10693 27666 10696
rect 27608 10687 27666 10693
rect 28994 10684 29000 10696
rect 29052 10684 29058 10736
rect 29362 10684 29368 10736
rect 29420 10684 29426 10736
rect 29549 10727 29607 10733
rect 29549 10693 29561 10727
rect 29595 10693 29607 10727
rect 29549 10687 29607 10693
rect 9272 10628 9812 10656
rect 9272 10616 9278 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12492 10628 12817 10656
rect 12492 10616 12498 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 28166 10616 28172 10668
rect 28224 10656 28230 10668
rect 28718 10656 28724 10668
rect 28224 10628 28724 10656
rect 28224 10616 28230 10628
rect 28718 10616 28724 10628
rect 28776 10656 28782 10668
rect 29564 10656 29592 10687
rect 28776 10628 29592 10656
rect 28776 10616 28782 10628
rect 32398 10616 32404 10668
rect 32456 10656 32462 10668
rect 32565 10659 32623 10665
rect 32565 10656 32577 10659
rect 32456 10628 32577 10656
rect 32456 10616 32462 10628
rect 32565 10625 32577 10628
rect 32611 10625 32623 10659
rect 32565 10619 32623 10625
rect 6644 10600 6696 10606
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3068 10520 3096 10551
rect 3142 10548 3148 10600
rect 3200 10548 3206 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3418 10588 3424 10600
rect 3375 10560 3424 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3418 10548 3424 10560
rect 3476 10588 3482 10600
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 3476 10560 4077 10588
rect 3476 10548 3482 10560
rect 4065 10557 4077 10560
rect 4111 10557 4123 10591
rect 4065 10551 4123 10557
rect 6644 10542 6696 10548
rect 9864 10600 9916 10606
rect 12348 10600 12400 10606
rect 9916 10560 12348 10588
rect 9864 10542 9916 10548
rect 24578 10548 24584 10600
rect 24636 10548 24642 10600
rect 27338 10548 27344 10600
rect 27396 10548 27402 10600
rect 32306 10548 32312 10600
rect 32364 10548 32370 10600
rect 12348 10542 12400 10548
rect 3234 10520 3240 10532
rect 3068 10492 3240 10520
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 3513 10523 3571 10529
rect 3513 10489 3525 10523
rect 3559 10520 3571 10523
rect 4246 10520 4252 10532
rect 3559 10492 4252 10520
rect 3559 10489 3571 10492
rect 3513 10483 3571 10489
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 3252 10452 3280 10480
rect 3602 10452 3608 10464
rect 3252 10424 3608 10452
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 10134 10412 10140 10464
rect 10192 10412 10198 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 14458 10452 14464 10464
rect 13863 10424 14464 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 29178 10412 29184 10464
rect 29236 10452 29242 10464
rect 29549 10455 29607 10461
rect 29549 10452 29561 10455
rect 29236 10424 29561 10452
rect 29236 10412 29242 10424
rect 29549 10421 29561 10424
rect 29595 10421 29607 10455
rect 29549 10415 29607 10421
rect 29733 10455 29791 10461
rect 29733 10421 29745 10455
rect 29779 10452 29791 10455
rect 30834 10452 30840 10464
rect 29779 10424 30840 10452
rect 29779 10421 29791 10424
rect 29733 10415 29791 10421
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 2832 10220 4169 10248
rect 2832 10208 2838 10220
rect 4157 10217 4169 10220
rect 4203 10248 4215 10251
rect 4522 10248 4528 10260
rect 4203 10220 4528 10248
rect 4203 10217 4215 10220
rect 4157 10211 4215 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 6730 10208 6736 10260
rect 6788 10208 6794 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9122 10248 9128 10260
rect 8619 10220 9128 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 23842 10248 23848 10260
rect 21315 10220 23848 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 23842 10208 23848 10220
rect 23900 10248 23906 10260
rect 24578 10248 24584 10260
rect 23900 10220 24584 10248
rect 23900 10208 23906 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 24949 10251 25007 10257
rect 24949 10217 24961 10251
rect 24995 10248 25007 10251
rect 25406 10248 25412 10260
rect 24995 10220 25412 10248
rect 24995 10217 25007 10220
rect 24949 10211 25007 10217
rect 25406 10208 25412 10220
rect 25464 10208 25470 10260
rect 27338 10208 27344 10260
rect 27396 10208 27402 10260
rect 28258 10208 28264 10260
rect 28316 10208 28322 10260
rect 28442 10208 28448 10260
rect 28500 10248 28506 10260
rect 29914 10248 29920 10260
rect 28500 10220 29920 10248
rect 28500 10208 28506 10220
rect 29914 10208 29920 10220
rect 29972 10248 29978 10260
rect 29972 10220 30052 10248
rect 29972 10208 29978 10220
rect 2133 10183 2191 10189
rect 2133 10149 2145 10183
rect 2179 10180 2191 10183
rect 2958 10180 2964 10192
rect 2179 10152 2964 10180
rect 2179 10149 2191 10152
rect 2133 10143 2191 10149
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 29733 10183 29791 10189
rect 29733 10180 29745 10183
rect 25608 10152 29745 10180
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 4246 10112 4252 10124
rect 2915 10084 4252 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 7190 10072 7196 10124
rect 7248 10072 7254 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 11112 10084 11253 10112
rect 11112 10072 11118 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2271 10016 2697 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 2700 9908 2728 10007
rect 2976 9976 3004 10007
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5902 10044 5908 10056
rect 5399 10016 5908 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 3142 9976 3148 9988
rect 2976 9948 3148 9976
rect 3142 9936 3148 9948
rect 3200 9976 3206 9988
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 3200 9948 3985 9976
rect 3200 9936 3206 9948
rect 3973 9945 3985 9948
rect 4019 9976 4031 9979
rect 4062 9976 4068 9988
rect 4019 9948 4068 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4189 9979 4247 9985
rect 4189 9945 4201 9979
rect 4235 9976 4247 9979
rect 4356 9976 4384 10004
rect 4235 9948 4384 9976
rect 4235 9945 4247 9948
rect 4189 9939 4247 9945
rect 3053 9911 3111 9917
rect 3053 9908 3065 9911
rect 2700 9880 3065 9908
rect 3053 9877 3065 9880
rect 3099 9877 3111 9911
rect 3053 9871 3111 9877
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3786 9908 3792 9920
rect 3283 9880 3792 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 5368 9908 5396 10007
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 11508 10047 11566 10053
rect 11508 10013 11520 10047
rect 11554 10044 11566 10047
rect 12066 10044 12072 10056
rect 11554 10016 12072 10044
rect 11554 10013 11566 10016
rect 11508 10007 11566 10013
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 25130 10053 25136 10056
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 25128 10044 25136 10053
rect 25091 10016 25136 10044
rect 22557 10007 22615 10013
rect 25128 10007 25136 10016
rect 5620 9979 5678 9985
rect 5620 9945 5632 9979
rect 5666 9976 5678 9979
rect 5810 9976 5816 9988
rect 5666 9948 5816 9976
rect 5666 9945 5678 9948
rect 5620 9939 5678 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 7466 9985 7472 9988
rect 7460 9976 7472 9985
rect 7427 9948 7472 9976
rect 7460 9939 7472 9948
rect 7524 9976 7530 9988
rect 9030 9976 9036 9988
rect 7524 9948 9036 9976
rect 7466 9936 7472 9939
rect 7524 9936 7530 9948
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 4387 9880 5396 9908
rect 22572 9908 22600 10007
rect 25130 10004 25136 10007
rect 25188 10004 25194 10056
rect 25314 10004 25320 10056
rect 25372 10004 25378 10056
rect 25608 10053 25636 10152
rect 29733 10149 29745 10152
rect 29779 10149 29791 10183
rect 29733 10143 29791 10149
rect 28534 10072 28540 10124
rect 28592 10112 28598 10124
rect 29086 10112 29092 10124
rect 28592 10084 28672 10112
rect 28592 10072 28598 10084
rect 25500 10047 25558 10053
rect 25500 10013 25512 10047
rect 25546 10013 25558 10047
rect 25500 10007 25558 10013
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10013 25651 10047
rect 25593 10007 25651 10013
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10044 26111 10047
rect 26602 10044 26608 10056
rect 26099 10016 26608 10044
rect 26099 10013 26111 10016
rect 26053 10007 26111 10013
rect 25222 9936 25228 9988
rect 25280 9936 25286 9988
rect 25516 9976 25544 10007
rect 25958 9976 25964 9988
rect 25516 9948 25964 9976
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 26068 9908 26096 10007
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 27706 10004 27712 10056
rect 27764 10044 27770 10056
rect 28442 10053 28448 10056
rect 28399 10047 28448 10053
rect 28399 10044 28411 10047
rect 27764 10016 28411 10044
rect 27764 10004 27770 10016
rect 28399 10013 28411 10016
rect 28445 10013 28448 10047
rect 28399 10007 28448 10013
rect 28442 10004 28448 10007
rect 28500 10004 28506 10056
rect 28644 10053 28672 10084
rect 28828 10084 29092 10112
rect 28828 10053 28856 10084
rect 29086 10072 29092 10084
rect 29144 10072 29150 10124
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 28812 10047 28870 10053
rect 28812 10013 28824 10047
rect 28858 10013 28870 10047
rect 28812 10007 28870 10013
rect 28902 10004 28908 10056
rect 28960 10004 28966 10056
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 30024 10044 30052 10220
rect 32306 10208 32312 10260
rect 32364 10248 32370 10260
rect 32493 10251 32551 10257
rect 32493 10248 32505 10251
rect 32364 10220 32505 10248
rect 32364 10208 32370 10220
rect 32493 10217 32505 10220
rect 32539 10217 32551 10251
rect 32493 10211 32551 10217
rect 30374 10072 30380 10124
rect 30432 10112 30438 10124
rect 30926 10112 30932 10124
rect 30432 10084 30932 10112
rect 30432 10072 30438 10084
rect 30926 10072 30932 10084
rect 30984 10112 30990 10124
rect 30984 10084 33732 10112
rect 30984 10072 30990 10084
rect 30101 10047 30159 10053
rect 30101 10044 30113 10047
rect 30024 10016 30113 10044
rect 29917 10007 29975 10013
rect 30101 10013 30113 10016
rect 30147 10013 30159 10047
rect 30101 10007 30159 10013
rect 28537 9979 28595 9985
rect 28537 9945 28549 9979
rect 28583 9945 28595 9979
rect 28537 9939 28595 9945
rect 22572 9880 26096 9908
rect 28552 9908 28580 9939
rect 28718 9936 28724 9988
rect 28776 9976 28782 9988
rect 29932 9976 29960 10007
rect 30282 10004 30288 10056
rect 30340 10004 30346 10056
rect 33410 10004 33416 10056
rect 33468 10004 33474 10056
rect 33704 10053 33732 10084
rect 33689 10047 33747 10053
rect 33689 10013 33701 10047
rect 33735 10013 33747 10047
rect 33689 10007 33747 10013
rect 28776 9948 29960 9976
rect 30009 9979 30067 9985
rect 28776 9936 28782 9948
rect 30009 9945 30021 9979
rect 30055 9945 30067 9979
rect 30009 9939 30067 9945
rect 29086 9908 29092 9920
rect 28552 9880 29092 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 30024 9908 30052 9939
rect 31202 9936 31208 9988
rect 31260 9936 31266 9988
rect 33505 9911 33563 9917
rect 33505 9908 33517 9911
rect 30024 9880 33517 9908
rect 33505 9877 33517 9880
rect 33551 9908 33563 9911
rect 33686 9908 33692 9920
rect 33551 9880 33692 9908
rect 33551 9877 33563 9880
rect 33505 9871 33563 9877
rect 33686 9868 33692 9880
rect 33744 9868 33750 9920
rect 33870 9868 33876 9920
rect 33928 9868 33934 9920
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3016 9676 4200 9704
rect 3016 9664 3022 9676
rect 4172 9645 4200 9676
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 5185 9707 5243 9713
rect 5185 9704 5197 9707
rect 4396 9676 5197 9704
rect 4396 9664 4402 9676
rect 5185 9673 5197 9676
rect 5231 9673 5243 9707
rect 5185 9667 5243 9673
rect 8573 9707 8631 9713
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 8846 9704 8852 9716
rect 8619 9676 8852 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 27709 9707 27767 9713
rect 27709 9673 27721 9707
rect 27755 9704 27767 9707
rect 28902 9704 28908 9716
rect 27755 9676 28908 9704
rect 27755 9673 27767 9676
rect 27709 9667 27767 9673
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9636 2007 9639
rect 4157 9639 4215 9645
rect 1995 9608 4108 9636
rect 1995 9605 2007 9608
rect 1949 9599 2007 9605
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 3142 9568 3148 9580
rect 2455 9540 3148 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2148 9432 2176 9531
rect 2332 9500 2360 9531
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3510 9568 3516 9580
rect 3283 9540 3516 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3510 9528 3516 9540
rect 3568 9568 3574 9580
rect 4080 9577 4108 9608
rect 4157 9605 4169 9639
rect 4203 9605 4215 9639
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4157 9599 4215 9605
rect 4448 9608 4997 9636
rect 4065 9571 4123 9577
rect 3568 9540 4016 9568
rect 3568 9528 3574 9540
rect 2774 9500 2780 9512
rect 2332 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9500 2838 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2832 9472 3341 9500
rect 2832 9460 2838 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3418 9460 3424 9512
rect 3476 9460 3482 9512
rect 2682 9432 2688 9444
rect 2148 9404 2688 9432
rect 2682 9392 2688 9404
rect 2740 9432 2746 9444
rect 3234 9432 3240 9444
rect 2740 9404 3240 9432
rect 2740 9392 2746 9404
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 3988 9364 4016 9540
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 4304 9540 4353 9568
rect 4304 9528 4310 9540
rect 4341 9537 4353 9540
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4448 9432 4476 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 11968 9639 12026 9645
rect 5960 9608 10824 9636
rect 5960 9596 5966 9608
rect 4522 9528 4528 9580
rect 4580 9528 4586 9580
rect 7208 9577 7236 9608
rect 7466 9577 7472 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7460 9568 7472 9577
rect 7427 9540 7472 9568
rect 7193 9531 7251 9537
rect 7460 9531 7472 9540
rect 7466 9528 7472 9531
rect 7524 9528 7530 9580
rect 10796 9512 10824 9608
rect 11968 9605 11980 9639
rect 12014 9636 12026 9639
rect 12066 9636 12072 9648
rect 12014 9608 12072 9636
rect 12014 9605 12026 9608
rect 11968 9599 12026 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16264 9608 17172 9636
rect 16264 9596 16270 9608
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17144 9568 17172 9608
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 20993 9639 21051 9645
rect 17276 9608 20760 9636
rect 17276 9596 17282 9608
rect 17310 9568 17316 9580
rect 17144 9540 17316 9568
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 17828 9540 19441 9568
rect 17828 9528 17834 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 10836 9472 11713 9500
rect 10836 9460 10842 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 19628 9500 19656 9531
rect 17920 9472 19656 9500
rect 19720 9500 19748 9531
rect 19794 9528 19800 9580
rect 19852 9528 19858 9580
rect 20732 9577 20760 9608
rect 20993 9605 21005 9639
rect 21039 9636 21051 9639
rect 21266 9636 21272 9648
rect 21039 9608 21272 9636
rect 21039 9605 21051 9608
rect 20993 9599 21051 9605
rect 21266 9596 21272 9608
rect 21324 9636 21330 9648
rect 22373 9639 22431 9645
rect 22373 9636 22385 9639
rect 21324 9608 22385 9636
rect 21324 9596 21330 9608
rect 22373 9605 22385 9608
rect 22419 9605 22431 9639
rect 22373 9599 22431 9605
rect 25130 9596 25136 9648
rect 25188 9636 25194 9648
rect 27341 9639 27399 9645
rect 27341 9636 27353 9639
rect 25188 9608 27353 9636
rect 25188 9596 25194 9608
rect 27341 9605 27353 9608
rect 27387 9605 27399 9639
rect 27341 9599 27399 9605
rect 30834 9596 30840 9648
rect 30892 9636 30898 9648
rect 32401 9639 32459 9645
rect 32401 9636 32413 9639
rect 30892 9608 32413 9636
rect 30892 9596 30898 9608
rect 32401 9605 32413 9608
rect 32447 9605 32459 9639
rect 32401 9599 32459 9605
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 20718 9571 20776 9577
rect 20718 9537 20730 9571
rect 20764 9537 20776 9571
rect 20718 9531 20776 9537
rect 20640 9500 20668 9531
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20864 9540 20913 9568
rect 20864 9528 20870 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21082 9528 21088 9580
rect 21140 9577 21146 9580
rect 21140 9568 21148 9577
rect 22189 9571 22247 9577
rect 21140 9540 21185 9568
rect 21140 9531 21148 9540
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 21140 9528 21146 9531
rect 20990 9500 20996 9512
rect 19720 9472 20576 9500
rect 20640 9472 20996 9500
rect 17920 9460 17926 9472
rect 4120 9404 4476 9432
rect 4120 9392 4126 9404
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 5132 9404 5365 9432
rect 5132 9392 5138 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13081 9435 13139 9441
rect 13081 9432 13093 9435
rect 12860 9404 13093 9432
rect 12860 9392 12866 9404
rect 13081 9401 13093 9404
rect 13127 9401 13139 9435
rect 13081 9395 13139 9401
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 18598 9432 18604 9444
rect 16080 9404 18604 9432
rect 16080 9392 16086 9404
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 19886 9392 19892 9444
rect 19944 9432 19950 9444
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 19944 9404 19993 9432
rect 19944 9392 19950 9404
rect 19981 9401 19993 9404
rect 20027 9401 20039 9435
rect 20548 9432 20576 9472
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 21284 9472 22140 9500
rect 21174 9432 21180 9444
rect 20548 9404 21180 9432
rect 19981 9395 20039 9401
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 3988 9336 5181 9364
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 19334 9364 19340 9376
rect 17644 9336 19340 9364
rect 17644 9324 17650 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 21284 9373 21312 9472
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21416 9336 22017 9364
rect 21416 9324 21422 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22112 9364 22140 9472
rect 22204 9432 22232 9531
rect 22462 9528 22468 9580
rect 22520 9528 22526 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26016 9540 27169 9568
rect 26016 9528 26022 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9568 27583 9571
rect 28718 9568 28724 9580
rect 27571 9540 28724 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 27448 9500 27476 9531
rect 28718 9528 28724 9540
rect 28776 9528 28782 9580
rect 30190 9528 30196 9580
rect 30248 9568 30254 9580
rect 31294 9574 31300 9580
rect 31128 9568 31300 9574
rect 30248 9546 31300 9568
rect 30248 9540 31156 9546
rect 30248 9528 30254 9540
rect 31294 9528 31300 9546
rect 31352 9528 31358 9580
rect 31386 9528 31392 9580
rect 31444 9528 31450 9580
rect 31478 9528 31484 9580
rect 31536 9577 31542 9580
rect 31536 9571 31585 9577
rect 31536 9537 31539 9571
rect 31573 9537 31585 9571
rect 31536 9531 31585 9537
rect 31536 9528 31542 9531
rect 27448 9472 28994 9500
rect 23750 9432 23756 9444
rect 22204 9404 23756 9432
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 28966 9432 28994 9472
rect 31386 9432 31392 9444
rect 28966 9404 31392 9432
rect 31386 9392 31392 9404
rect 31444 9392 31450 9444
rect 31938 9392 31944 9444
rect 31996 9432 32002 9444
rect 33689 9435 33747 9441
rect 33689 9432 33701 9435
rect 31996 9404 33701 9432
rect 31996 9392 32002 9404
rect 33689 9401 33701 9404
rect 33735 9401 33747 9435
rect 33689 9395 33747 9401
rect 25038 9364 25044 9376
rect 22112 9336 25044 9364
rect 22005 9327 22063 9333
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 31754 9324 31760 9376
rect 31812 9324 31818 9376
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 2774 9120 2780 9172
rect 2832 9120 2838 9172
rect 2958 9120 2964 9172
rect 3016 9120 3022 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12526 9160 12532 9172
rect 12207 9132 12532 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 17218 9160 17224 9172
rect 15611 9132 17224 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 18877 9163 18935 9169
rect 17736 9132 18368 9160
rect 17736 9120 17742 9132
rect 2792 9024 2820 9120
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 17368 9064 17908 9092
rect 17368 9052 17374 9064
rect 3970 9024 3976 9036
rect 2792 8996 3976 9024
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8956 3387 8959
rect 3602 8956 3608 8968
rect 3375 8928 3608 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4338 8956 4344 8968
rect 4203 8928 4344 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 16689 8959 16747 8965
rect 16689 8925 16701 8959
rect 16735 8956 16747 8959
rect 16850 8956 16856 8968
rect 16735 8928 16856 8956
rect 16735 8925 16747 8928
rect 16689 8919 16747 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 16942 8916 16948 8968
rect 17000 8916 17006 8968
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 17770 8916 17776 8968
rect 17828 8916 17834 8968
rect 17880 8965 17908 9064
rect 18340 8965 18368 9132
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19610 9160 19616 9172
rect 18923 9132 19616 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 19904 9132 21220 9160
rect 19334 9052 19340 9104
rect 19392 9092 19398 9104
rect 19904 9092 19932 9132
rect 19392 9064 19932 9092
rect 21192 9092 21220 9132
rect 21266 9120 21272 9172
rect 21324 9120 21330 9172
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 22462 9160 22468 9172
rect 21600 9132 22468 9160
rect 21600 9120 21606 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 33686 9120 33692 9172
rect 33744 9120 33750 9172
rect 22738 9092 22744 9104
rect 21192 9064 22744 9092
rect 19392 9052 19398 9064
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 26694 9024 26700 9036
rect 22066 8996 26700 9024
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 2866 8848 2872 8900
rect 2924 8897 2930 8900
rect 2924 8891 2973 8897
rect 2924 8857 2927 8891
rect 2961 8857 2973 8891
rect 2924 8851 2973 8857
rect 11048 8891 11106 8897
rect 11048 8857 11060 8891
rect 11094 8888 11106 8891
rect 11146 8888 11152 8900
rect 11094 8860 11152 8888
rect 11094 8857 11106 8860
rect 11048 8851 11106 8857
rect 2924 8848 2930 8851
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 15378 8848 15384 8900
rect 15436 8888 15442 8900
rect 17788 8888 17816 8916
rect 15436 8860 17816 8888
rect 17880 8888 17908 8919
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 19889 8959 19947 8965
rect 18748 8928 19840 8956
rect 18748 8916 18754 8928
rect 18414 8888 18420 8900
rect 17880 8860 18420 8888
rect 15436 8848 15442 8860
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 18509 8891 18567 8897
rect 18509 8857 18521 8891
rect 18555 8857 18567 8891
rect 18509 8851 18567 8857
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8888 18659 8891
rect 18782 8888 18788 8900
rect 18647 8860 18788 8888
rect 18647 8857 18659 8860
rect 18601 8851 18659 8857
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17862 8820 17868 8832
rect 16724 8792 17868 8820
rect 16724 8780 16730 8792
rect 17862 8780 17868 8792
rect 17920 8820 17926 8832
rect 18524 8820 18552 8851
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 19812 8888 19840 8928
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 19978 8956 19984 8968
rect 19935 8928 19984 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20156 8959 20214 8965
rect 20156 8925 20168 8959
rect 20202 8956 20214 8959
rect 21358 8956 21364 8968
rect 20202 8928 21364 8956
rect 20202 8925 20214 8928
rect 20156 8919 20214 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 19812 8860 20760 8888
rect 20622 8820 20628 8832
rect 17920 8792 20628 8820
rect 17920 8780 17926 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20732 8820 20760 8860
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 22066 8888 22094 8996
rect 26694 8984 26700 8996
rect 26752 8984 26758 9036
rect 29822 9024 29828 9036
rect 28920 8996 29828 9024
rect 24026 8916 24032 8968
rect 24084 8956 24090 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24084 8928 24593 8956
rect 24084 8916 24090 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 21048 8860 22094 8888
rect 24596 8888 24624 8919
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 28920 8965 28948 8996
rect 29822 8984 29828 8996
rect 29880 8984 29886 9036
rect 28905 8959 28963 8965
rect 28905 8956 28917 8959
rect 27672 8928 28917 8956
rect 27672 8916 27678 8928
rect 28905 8925 28917 8928
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 28994 8916 29000 8968
rect 29052 8956 29058 8968
rect 29181 8959 29239 8965
rect 29181 8956 29193 8959
rect 29052 8928 29193 8956
rect 29052 8916 29058 8928
rect 29181 8925 29193 8928
rect 29227 8956 29239 8959
rect 30190 8956 30196 8968
rect 29227 8928 30196 8956
rect 29227 8925 29239 8928
rect 29181 8919 29239 8925
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 32306 8916 32312 8968
rect 32364 8916 32370 8968
rect 32576 8959 32634 8965
rect 32576 8925 32588 8959
rect 32622 8956 32634 8959
rect 33870 8956 33876 8968
rect 32622 8928 33876 8956
rect 32622 8925 32634 8928
rect 32576 8919 32634 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 26050 8888 26056 8900
rect 24596 8860 26056 8888
rect 21048 8848 21054 8860
rect 26050 8848 26056 8860
rect 26108 8848 26114 8900
rect 21082 8820 21088 8832
rect 20732 8792 21088 8820
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 23658 8780 23664 8832
rect 23716 8820 23722 8832
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 23716 8792 24685 8820
rect 23716 8780 23722 8792
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 25041 8823 25099 8829
rect 25041 8820 25053 8823
rect 25004 8792 25053 8820
rect 25004 8780 25010 8792
rect 25041 8789 25053 8792
rect 25087 8789 25099 8823
rect 25041 8783 25099 8789
rect 28718 8780 28724 8832
rect 28776 8780 28782 8832
rect 29086 8780 29092 8832
rect 29144 8820 29150 8832
rect 29730 8820 29736 8832
rect 29144 8792 29736 8820
rect 29144 8780 29150 8792
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3510 8616 3516 8628
rect 3467 8588 3516 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 16574 8616 16580 8628
rect 16255 8588 16580 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16574 8576 16580 8588
rect 16632 8616 16638 8628
rect 17678 8616 17684 8628
rect 16632 8588 17684 8616
rect 16632 8576 16638 8588
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18472 8588 20760 8616
rect 18472 8576 18478 8588
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 9364 8520 9597 8548
rect 9364 8508 9370 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 15197 8551 15255 8557
rect 15197 8517 15209 8551
rect 15243 8517 15255 8551
rect 15197 8511 15255 8517
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8548 15439 8551
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 15427 8520 18245 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 18233 8517 18245 8520
rect 18279 8548 18291 8551
rect 18322 8548 18328 8560
rect 18279 8520 18328 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 3292 8452 3525 8480
rect 3292 8440 3298 8452
rect 3513 8449 3525 8452
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3970 8440 3976 8492
rect 4028 8440 4034 8492
rect 15212 8412 15240 8511
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 16264 8452 16313 8480
rect 16264 8440 16270 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16666 8480 16672 8492
rect 16301 8443 16359 8449
rect 16408 8452 16672 8480
rect 16408 8412 16436 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8480 17831 8483
rect 18432 8480 18460 8576
rect 19981 8551 20039 8557
rect 19981 8517 19993 8551
rect 20027 8548 20039 8551
rect 20530 8548 20536 8560
rect 20027 8520 20536 8548
rect 20027 8517 20039 8520
rect 19981 8511 20039 8517
rect 20530 8508 20536 8520
rect 20588 8508 20594 8560
rect 20622 8508 20628 8560
rect 20680 8508 20686 8560
rect 20732 8548 20760 8588
rect 20990 8576 20996 8628
rect 21048 8576 21054 8628
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 23658 8616 23664 8628
rect 21232 8588 23664 8616
rect 21232 8576 21238 8588
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 23750 8576 23756 8628
rect 23808 8616 23814 8628
rect 23808 8588 25176 8616
rect 23808 8576 23814 8588
rect 22462 8548 22468 8560
rect 20732 8520 22468 8548
rect 22462 8508 22468 8520
rect 22520 8508 22526 8560
rect 22554 8508 22560 8560
rect 22612 8548 22618 8560
rect 22741 8551 22799 8557
rect 22741 8548 22753 8551
rect 22612 8520 22753 8548
rect 22612 8508 22618 8520
rect 22741 8517 22753 8520
rect 22787 8517 22799 8551
rect 22741 8511 22799 8517
rect 22925 8551 22983 8557
rect 22925 8517 22937 8551
rect 22971 8517 22983 8551
rect 22925 8511 22983 8517
rect 17819 8452 18460 8480
rect 20441 8483 20499 8489
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 20441 8449 20453 8483
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 15212 8384 16436 8412
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17696 8412 17724 8443
rect 20456 8412 20484 8443
rect 20714 8440 20720 8492
rect 20772 8440 20778 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 21082 8480 21088 8492
rect 20855 8452 21088 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 16540 8384 20484 8412
rect 16540 8372 16546 8384
rect 15013 8347 15071 8353
rect 15013 8313 15025 8347
rect 15059 8344 15071 8347
rect 15286 8344 15292 8356
rect 15059 8316 15292 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15838 8304 15844 8356
rect 15896 8304 15902 8356
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 16080 8316 17325 8344
rect 16080 8304 16086 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 19794 8304 19800 8356
rect 19852 8344 19858 8356
rect 22940 8344 22968 8511
rect 24670 8508 24676 8560
rect 24728 8548 24734 8560
rect 25148 8548 25176 8588
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25866 8616 25872 8628
rect 25280 8588 25872 8616
rect 25280 8576 25286 8588
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 31386 8576 31392 8628
rect 31444 8616 31450 8628
rect 33689 8619 33747 8625
rect 33689 8616 33701 8619
rect 31444 8588 33701 8616
rect 31444 8576 31450 8588
rect 33689 8585 33701 8588
rect 33735 8585 33747 8619
rect 33689 8579 33747 8585
rect 24728 8520 25084 8548
rect 25148 8520 25728 8548
rect 24728 8508 24734 8520
rect 24785 8483 24843 8489
rect 24785 8449 24797 8483
rect 24831 8480 24843 8483
rect 24946 8480 24952 8492
rect 24831 8452 24952 8480
rect 24831 8449 24843 8452
rect 24785 8443 24843 8449
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 25056 8489 25084 8520
rect 25700 8489 25728 8520
rect 30006 8508 30012 8560
rect 30064 8548 30070 8560
rect 30282 8548 30288 8560
rect 30064 8520 30288 8548
rect 30064 8508 30070 8520
rect 30282 8508 30288 8520
rect 30340 8548 30346 8560
rect 30561 8551 30619 8557
rect 30561 8548 30573 8551
rect 30340 8520 30573 8548
rect 30340 8508 30346 8520
rect 30561 8517 30573 8520
rect 30607 8517 30619 8551
rect 30561 8511 30619 8517
rect 31754 8508 31760 8560
rect 31812 8548 31818 8560
rect 32554 8551 32612 8557
rect 32554 8548 32566 8551
rect 31812 8520 32566 8548
rect 31812 8508 31818 8520
rect 32554 8517 32566 8520
rect 32600 8517 32612 8551
rect 32554 8511 32612 8517
rect 25041 8483 25099 8489
rect 25041 8449 25053 8483
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8480 26019 8483
rect 26050 8480 26056 8492
rect 26007 8452 26056 8480
rect 26007 8449 26019 8452
rect 25961 8443 26019 8449
rect 26050 8440 26056 8452
rect 26108 8440 26114 8492
rect 28166 8440 28172 8492
rect 28224 8480 28230 8492
rect 28609 8483 28667 8489
rect 28609 8480 28621 8483
rect 28224 8452 28621 8480
rect 28224 8440 28230 8452
rect 28609 8449 28621 8452
rect 28655 8449 28667 8483
rect 28609 8443 28667 8449
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 30193 8483 30251 8489
rect 30193 8480 30205 8483
rect 28960 8452 30205 8480
rect 28960 8440 28966 8452
rect 30193 8449 30205 8452
rect 30239 8449 30251 8483
rect 30193 8443 30251 8449
rect 30374 8440 30380 8492
rect 30432 8440 30438 8492
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8480 30711 8483
rect 31294 8480 31300 8492
rect 30699 8452 31300 8480
rect 30699 8449 30711 8452
rect 30653 8443 30711 8449
rect 31294 8440 31300 8452
rect 31352 8440 31358 8492
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 32306 8372 32312 8424
rect 32364 8372 32370 8424
rect 19852 8316 22968 8344
rect 23109 8347 23167 8353
rect 19852 8304 19858 8316
rect 23109 8313 23121 8347
rect 23155 8344 23167 8347
rect 24026 8344 24032 8356
rect 23155 8316 24032 8344
rect 23155 8313 23167 8316
rect 23109 8307 23167 8313
rect 24026 8304 24032 8316
rect 24084 8304 24090 8356
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 25188 8316 25513 8344
rect 25188 8304 25194 8316
rect 25501 8313 25513 8316
rect 25547 8313 25559 8347
rect 29733 8347 29791 8353
rect 29733 8344 29745 8347
rect 25501 8307 25559 8313
rect 29288 8316 29745 8344
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8294 8276 8300 8288
rect 8159 8248 8300 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8294 8236 8300 8248
rect 8352 8276 8358 8288
rect 9858 8276 9864 8288
rect 8352 8248 9864 8276
rect 8352 8236 8358 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 19058 8276 19064 8288
rect 15252 8248 19064 8276
rect 15252 8236 15258 8248
rect 19058 8236 19064 8248
rect 19116 8276 19122 8288
rect 20622 8276 20628 8288
rect 19116 8248 20628 8276
rect 19116 8236 19122 8248
rect 20622 8236 20628 8248
rect 20680 8276 20686 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 20680 8248 22937 8276
rect 20680 8236 20686 8248
rect 22925 8245 22937 8248
rect 22971 8245 22983 8279
rect 22925 8239 22983 8245
rect 27890 8236 27896 8288
rect 27948 8276 27954 8288
rect 29288 8276 29316 8316
rect 29733 8313 29745 8316
rect 29779 8313 29791 8347
rect 29733 8307 29791 8313
rect 27948 8248 29316 8276
rect 27948 8236 27954 8248
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 16942 8032 16948 8084
rect 17000 8032 17006 8084
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 23753 8075 23811 8081
rect 23753 8072 23765 8075
rect 22612 8044 23765 8072
rect 22612 8032 22618 8044
rect 23753 8041 23765 8044
rect 23799 8072 23811 8075
rect 26878 8072 26884 8084
rect 23799 8044 26884 8072
rect 23799 8041 23811 8044
rect 23753 8035 23811 8041
rect 26878 8032 26884 8044
rect 26936 8032 26942 8084
rect 29178 8032 29184 8084
rect 29236 8072 29242 8084
rect 29917 8075 29975 8081
rect 29917 8072 29929 8075
rect 29236 8044 29929 8072
rect 29236 8032 29242 8044
rect 29917 8041 29929 8044
rect 29963 8041 29975 8075
rect 29917 8035 29975 8041
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32493 8075 32551 8081
rect 32493 8072 32505 8075
rect 32364 8044 32505 8072
rect 32364 8032 32370 8044
rect 32493 8041 32505 8044
rect 32539 8041 32551 8075
rect 32493 8035 32551 8041
rect 23382 7964 23388 8016
rect 23440 8004 23446 8016
rect 25869 8007 25927 8013
rect 25869 8004 25881 8007
rect 23440 7976 25881 8004
rect 23440 7964 23446 7976
rect 25869 7973 25881 7976
rect 25915 7973 25927 8007
rect 25869 7967 25927 7973
rect 8294 7936 8300 7948
rect 7116 7908 8300 7936
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 7116 7877 7144 7908
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 21542 7936 21548 7948
rect 18892 7908 21548 7936
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 3108 7840 7113 7868
rect 3108 7828 3114 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 8202 7868 8208 7880
rect 7331 7840 8208 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 4062 7800 4068 7812
rect 3660 7772 4068 7800
rect 3660 7760 3666 7772
rect 4062 7760 4068 7772
rect 4120 7800 4126 7812
rect 7300 7800 7328 7831
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10594 7868 10600 7880
rect 10091 7840 10600 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 18892 7877 18920 7908
rect 21542 7896 21548 7908
rect 21600 7896 21606 7948
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7837 18935 7871
rect 18877 7831 18935 7837
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 20036 7840 22385 7868
rect 20036 7828 20042 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 24026 7828 24032 7880
rect 24084 7868 24090 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24084 7840 24593 7868
rect 24084 7828 24090 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 31202 7828 31208 7880
rect 31260 7828 31266 7880
rect 4120 7772 7328 7800
rect 4120 7760 4126 7772
rect 7374 7760 7380 7812
rect 7432 7760 7438 7812
rect 10137 7803 10195 7809
rect 10137 7769 10149 7803
rect 10183 7800 10195 7803
rect 10226 7800 10232 7812
rect 10183 7772 10232 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 15657 7803 15715 7809
rect 15657 7769 15669 7803
rect 15703 7800 15715 7803
rect 16298 7800 16304 7812
rect 15703 7772 16304 7800
rect 15703 7769 15715 7772
rect 15657 7763 15715 7769
rect 16298 7760 16304 7772
rect 16356 7760 16362 7812
rect 18417 7803 18475 7809
rect 18417 7769 18429 7803
rect 18463 7800 18475 7803
rect 19702 7800 19708 7812
rect 18463 7772 19708 7800
rect 18463 7769 18475 7772
rect 18417 7763 18475 7769
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 20165 7803 20223 7809
rect 20165 7769 20177 7803
rect 20211 7800 20223 7803
rect 20530 7800 20536 7812
rect 20211 7772 20536 7800
rect 20211 7769 20223 7772
rect 20165 7763 20223 7769
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 22640 7803 22698 7809
rect 22640 7769 22652 7803
rect 22686 7800 22698 7803
rect 22922 7800 22928 7812
rect 22686 7772 22928 7800
rect 22686 7769 22698 7772
rect 22640 7763 22698 7769
rect 22922 7760 22928 7772
rect 22980 7760 22986 7812
rect 28537 7803 28595 7809
rect 28537 7769 28549 7803
rect 28583 7800 28595 7803
rect 28810 7800 28816 7812
rect 28583 7772 28816 7800
rect 28583 7769 28595 7772
rect 28537 7763 28595 7769
rect 28810 7760 28816 7772
rect 28868 7760 28874 7812
rect 29362 7760 29368 7812
rect 29420 7800 29426 7812
rect 29733 7803 29791 7809
rect 29733 7800 29745 7803
rect 29420 7772 29745 7800
rect 29420 7760 29426 7772
rect 29733 7769 29745 7772
rect 29779 7769 29791 7803
rect 29733 7763 29791 7769
rect 29914 7760 29920 7812
rect 29972 7760 29978 7812
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 18932 7704 21465 7732
rect 18932 7692 18938 7704
rect 21453 7701 21465 7704
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 27249 7735 27307 7741
rect 27249 7701 27261 7735
rect 27295 7732 27307 7735
rect 28350 7732 28356 7744
rect 27295 7704 28356 7732
rect 27295 7701 27307 7704
rect 27249 7695 27307 7701
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 30101 7735 30159 7741
rect 30101 7701 30113 7735
rect 30147 7732 30159 7735
rect 30558 7732 30564 7744
rect 30147 7704 30564 7732
rect 30147 7701 30159 7704
rect 30101 7695 30159 7701
rect 30558 7692 30564 7704
rect 30616 7692 30622 7744
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15378 7528 15384 7540
rect 14967 7500 15384 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 16206 7528 16212 7540
rect 15948 7500 16212 7528
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 6822 7460 6828 7472
rect 5868 7432 6828 7460
rect 5868 7420 5874 7432
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 10226 7420 10232 7472
rect 10284 7420 10290 7472
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 11946 7463 12004 7469
rect 11946 7460 11958 7463
rect 11204 7432 11958 7460
rect 11204 7420 11210 7432
rect 11946 7429 11958 7432
rect 11992 7429 12004 7463
rect 15948 7460 15976 7500
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 21082 7528 21088 7540
rect 20763 7500 21088 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 25958 7488 25964 7540
rect 26016 7488 26022 7540
rect 27801 7531 27859 7537
rect 27801 7497 27813 7531
rect 27847 7528 27859 7531
rect 27890 7528 27896 7540
rect 27847 7500 27896 7528
rect 27847 7497 27859 7500
rect 27801 7491 27859 7497
rect 27890 7488 27896 7500
rect 27948 7488 27954 7540
rect 28166 7488 28172 7540
rect 28224 7488 28230 7540
rect 11946 7423 12004 7429
rect 13556 7432 15976 7460
rect 16056 7463 16114 7469
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 3878 7392 3884 7404
rect 2556 7364 3884 7392
rect 2556 7352 2562 7364
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 8386 7324 8392 7336
rect 6595 7296 8392 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 8386 7284 8392 7296
rect 8444 7324 8450 7336
rect 8938 7324 8944 7336
rect 8444 7296 8944 7324
rect 8444 7284 8450 7296
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 11164 7324 11192 7420
rect 13556 7401 13584 7432
rect 16056 7429 16068 7463
rect 16102 7460 16114 7463
rect 17402 7460 17408 7472
rect 16102 7432 17408 7460
rect 16102 7429 16114 7432
rect 16056 7423 16114 7429
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 18874 7460 18880 7472
rect 18288 7432 18880 7460
rect 18288 7420 18294 7432
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 19978 7420 19984 7472
rect 20036 7420 20042 7472
rect 20898 7420 20904 7472
rect 20956 7420 20962 7472
rect 23382 7420 23388 7472
rect 23440 7420 23446 7472
rect 24854 7420 24860 7472
rect 24912 7460 24918 7472
rect 24912 7432 28028 7460
rect 24912 7420 24918 7432
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 15194 7392 15200 7404
rect 13771 7364 15200 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16942 7392 16948 7404
rect 16347 7364 16948 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 22738 7352 22744 7404
rect 22796 7392 22802 7404
rect 24872 7392 24900 7420
rect 22796 7364 24900 7392
rect 25777 7395 25835 7401
rect 22796 7352 22802 7364
rect 25777 7361 25789 7395
rect 25823 7361 25835 7395
rect 25777 7355 25835 7361
rect 9263 7296 11192 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 11698 7284 11704 7336
rect 11756 7284 11762 7336
rect 25792 7324 25820 7355
rect 26050 7352 26056 7404
rect 26108 7352 26114 7404
rect 28000 7401 28028 7432
rect 30558 7420 30564 7472
rect 30616 7420 30622 7472
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7361 28043 7395
rect 28994 7392 29000 7404
rect 27985 7355 28043 7361
rect 28736 7364 29000 7392
rect 27614 7324 27620 7336
rect 25792 7296 27620 7324
rect 27614 7284 27620 7296
rect 27672 7284 27678 7336
rect 27724 7324 27752 7355
rect 28736 7324 28764 7364
rect 28994 7352 29000 7364
rect 29052 7352 29058 7404
rect 27724 7296 28764 7324
rect 28810 7284 28816 7336
rect 28868 7284 28874 7336
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 13541 7259 13599 7265
rect 13541 7256 13553 7259
rect 12952 7228 13553 7256
rect 12952 7216 12958 7228
rect 13541 7225 13553 7228
rect 13587 7225 13599 7259
rect 13541 7219 13599 7225
rect 2590 7148 2596 7200
rect 2648 7148 2654 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8386 7188 8392 7200
rect 8343 7160 8392 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 10778 7188 10784 7200
rect 10735 7160 10784 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 20622 7148 20628 7200
rect 20680 7188 20686 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 20680 7160 20729 7188
rect 20680 7148 20686 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 25590 7148 25596 7200
rect 25648 7148 25654 7200
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 2498 6984 2504 6996
rect 1719 6956 2504 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3157 6987 3215 6993
rect 3157 6984 3169 6987
rect 2648 6956 3169 6984
rect 2648 6944 2654 6956
rect 3157 6953 3169 6956
rect 3203 6953 3215 6987
rect 3157 6947 3215 6953
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 20898 6984 20904 6996
rect 18380 6956 20904 6984
rect 18380 6944 18386 6956
rect 20898 6944 20904 6956
rect 20956 6944 20962 6996
rect 26050 6984 26056 6996
rect 24596 6956 26056 6984
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 10594 6916 10600 6928
rect 8260 6888 10600 6916
rect 8260 6876 8266 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 12710 6916 12716 6928
rect 12268 6888 12716 6916
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6817 3479 6851
rect 3421 6811 3479 6817
rect 2682 6672 2688 6724
rect 2740 6672 2746 6724
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3436 6712 3464 6811
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 8444 6820 10149 6848
rect 8444 6808 8450 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10137 6811 10195 6817
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10686 6848 10692 6860
rect 10468 6820 10692 6848
rect 10468 6808 10474 6820
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 12268 6857 12296 6888
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12299 6820 12333 6848
rect 21468 6820 21956 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 5074 6780 5080 6792
rect 4396 6752 5080 6780
rect 4396 6740 4402 6752
rect 5074 6740 5080 6752
rect 5132 6780 5138 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5132 6752 5457 6780
rect 5132 6740 5138 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5712 6783 5770 6789
rect 5712 6749 5724 6783
rect 5758 6780 5770 6783
rect 6822 6780 6828 6792
rect 5758 6752 6828 6780
rect 5758 6749 5770 6752
rect 5712 6743 5770 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 8404 6780 8432 6808
rect 7699 6752 8432 6780
rect 10229 6783 10287 6789
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 3200 6684 3464 6712
rect 6840 6684 7757 6712
rect 3200 6672 3206 6684
rect 6840 6653 6868 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 10244 6712 10272 6743
rect 10502 6740 10508 6792
rect 10560 6789 10566 6792
rect 10560 6783 10609 6789
rect 10560 6749 10563 6783
rect 10597 6749 10609 6783
rect 10560 6743 10609 6749
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 13078 6780 13084 6792
rect 12391 6752 13084 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 10560 6740 10566 6743
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19518 6780 19524 6792
rect 19475 6752 19524 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19702 6789 19708 6792
rect 19696 6743 19708 6789
rect 19702 6740 19708 6743
rect 19760 6740 19766 6792
rect 21468 6789 21496 6820
rect 21928 6792 21956 6820
rect 23474 6808 23480 6860
rect 23532 6848 23538 6860
rect 24596 6848 24624 6956
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 27154 6944 27160 6996
rect 27212 6984 27218 6996
rect 29362 6984 29368 6996
rect 27212 6956 29368 6984
rect 27212 6944 27218 6956
rect 29362 6944 29368 6956
rect 29420 6944 29426 6996
rect 27801 6919 27859 6925
rect 27801 6885 27813 6919
rect 27847 6885 27859 6919
rect 27801 6879 27859 6885
rect 23532 6820 23980 6848
rect 23532 6808 23538 6820
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21600 6752 21741 6780
rect 21600 6740 21606 6752
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 23952 6789 23980 6820
rect 24044 6820 24624 6848
rect 27816 6848 27844 6879
rect 27982 6848 27988 6860
rect 27816 6820 27988 6848
rect 24044 6789 24072 6820
rect 27982 6808 27988 6820
rect 28040 6808 28046 6860
rect 29104 6820 30144 6848
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 21968 6752 23765 6780
rect 21968 6740 21974 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 23753 6743 23811 6749
rect 23937 6783 23995 6789
rect 23937 6749 23949 6783
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24670 6780 24676 6792
rect 24627 6752 24676 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 10778 6712 10784 6724
rect 10244 6684 10784 6712
rect 7745 6675 7803 6681
rect 10778 6672 10784 6684
rect 10836 6712 10842 6724
rect 12437 6715 12495 6721
rect 12437 6712 12449 6715
rect 10836 6684 12449 6712
rect 10836 6672 10842 6684
rect 12437 6681 12449 6684
rect 12483 6681 12495 6715
rect 13354 6712 13360 6724
rect 12437 6675 12495 6681
rect 12728 6684 13360 6712
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 12728 6644 12756 6684
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 21637 6715 21695 6721
rect 21637 6712 21649 6715
rect 20772 6684 21649 6712
rect 20772 6672 20778 6684
rect 21637 6681 21649 6684
rect 21683 6681 21695 6715
rect 23768 6712 23796 6743
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 24848 6783 24906 6789
rect 24848 6749 24860 6783
rect 24894 6780 24906 6783
rect 25130 6780 25136 6792
rect 24894 6752 25136 6780
rect 24894 6749 24906 6752
rect 24848 6743 24906 6749
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 28000 6780 28028 6808
rect 29104 6780 29132 6820
rect 28000 6752 29132 6780
rect 29178 6740 29184 6792
rect 29236 6740 29242 6792
rect 30116 6789 30144 6820
rect 29917 6783 29975 6789
rect 29917 6749 29929 6783
rect 29963 6749 29975 6783
rect 29917 6743 29975 6749
rect 30101 6783 30159 6789
rect 30101 6749 30113 6783
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 28936 6715 28994 6721
rect 23768 6684 26096 6712
rect 21637 6675 21695 6681
rect 11011 6616 12756 6644
rect 12805 6647 12863 6653
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 12986 6644 12992 6656
rect 12851 6616 12992 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 16298 6644 16304 6656
rect 15896 6616 16304 6644
rect 15896 6604 15902 6616
rect 16298 6604 16304 6616
rect 16356 6644 16362 6656
rect 16577 6647 16635 6653
rect 16577 6644 16589 6647
rect 16356 6616 16589 6644
rect 16356 6604 16362 6616
rect 16577 6613 16589 6616
rect 16623 6613 16635 6647
rect 16577 6607 16635 6613
rect 18782 6604 18788 6656
rect 18840 6644 18846 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 18840 6616 20821 6644
rect 18840 6604 18846 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 21266 6604 21272 6656
rect 21324 6604 21330 6656
rect 23566 6604 23572 6656
rect 23624 6604 23630 6656
rect 25866 6604 25872 6656
rect 25924 6644 25930 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25924 6616 25973 6644
rect 25924 6604 25930 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 26068 6644 26096 6684
rect 28936 6681 28948 6715
rect 28982 6712 28994 6715
rect 29733 6715 29791 6721
rect 29733 6712 29745 6715
rect 28982 6684 29745 6712
rect 28982 6681 28994 6684
rect 28936 6675 28994 6681
rect 29733 6681 29745 6684
rect 29779 6681 29791 6715
rect 29733 6675 29791 6681
rect 29932 6644 29960 6743
rect 30190 6740 30196 6792
rect 30248 6740 30254 6792
rect 26068 6616 29960 6644
rect 25961 6607 26019 6613
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6440 6975 6443
rect 7282 6440 7288 6452
rect 6963 6412 7288 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 12894 6400 12900 6452
rect 12952 6400 12958 6452
rect 12986 6400 12992 6452
rect 13044 6400 13050 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 16482 6440 16488 6452
rect 16347 6412 16488 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20772 6412 20913 6440
rect 20772 6400 20778 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 20901 6403 20959 6409
rect 30006 6400 30012 6452
rect 30064 6400 30070 6452
rect 2682 6332 2688 6384
rect 2740 6372 2746 6384
rect 2777 6375 2835 6381
rect 2777 6372 2789 6375
rect 2740 6344 2789 6372
rect 2740 6332 2746 6344
rect 2777 6341 2789 6344
rect 2823 6341 2835 6375
rect 2777 6335 2835 6341
rect 3697 6375 3755 6381
rect 3697 6341 3709 6375
rect 3743 6372 3755 6375
rect 3878 6372 3884 6384
rect 3743 6344 3884 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7006 6372 7012 6384
rect 6871 6344 7012 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 15188 6375 15246 6381
rect 15188 6341 15200 6375
rect 15234 6372 15246 6375
rect 16022 6372 16028 6384
rect 15234 6344 16028 6372
rect 15234 6341 15246 6344
rect 15188 6335 15246 6341
rect 16022 6332 16028 6344
rect 16080 6332 16086 6384
rect 19788 6375 19846 6381
rect 19788 6341 19800 6375
rect 19834 6372 19846 6375
rect 21266 6372 21272 6384
rect 19834 6344 21272 6372
rect 19834 6341 19846 6344
rect 19788 6335 19846 6341
rect 21266 6332 21272 6344
rect 21324 6332 21330 6384
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 28902 6381 28908 6384
rect 24682 6375 24740 6381
rect 24682 6372 24694 6375
rect 23624 6344 24694 6372
rect 23624 6332 23630 6344
rect 24682 6341 24694 6344
rect 24728 6341 24740 6375
rect 28896 6372 28908 6381
rect 28863 6344 28908 6372
rect 24682 6335 24740 6341
rect 28896 6335 28908 6344
rect 28902 6332 28908 6335
rect 28960 6332 28966 6384
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 28350 6264 28356 6316
rect 28408 6304 28414 6316
rect 28629 6307 28687 6313
rect 28629 6304 28641 6307
rect 28408 6276 28641 6304
rect 28408 6264 28414 6276
rect 28629 6273 28641 6276
rect 28675 6273 28687 6307
rect 28629 6267 28687 6273
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 5868 6208 6653 6236
rect 5868 6196 5874 6208
rect 6641 6205 6653 6208
rect 6687 6236 6699 6239
rect 12342 6236 12348 6248
rect 6687 6208 12348 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12400 6208 12725 6236
rect 12400 6196 12406 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 14918 6196 14924 6248
rect 14976 6196 14982 6248
rect 19518 6196 19524 6248
rect 19576 6196 19582 6248
rect 24949 6239 25007 6245
rect 24949 6205 24961 6239
rect 24995 6205 25007 6239
rect 24949 6199 25007 6205
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 7331 6140 13492 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 3970 6100 3976 6112
rect 3835 6072 3976 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 13464 6100 13492 6140
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 23569 6171 23627 6177
rect 23569 6168 23581 6171
rect 23532 6140 23581 6168
rect 23532 6128 23538 6140
rect 23569 6137 23581 6140
rect 23615 6137 23627 6171
rect 23569 6131 23627 6137
rect 18414 6100 18420 6112
rect 13464 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24964 6100 24992 6199
rect 24728 6072 24992 6100
rect 24728 6060 24734 6072
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 20162 5896 20168 5908
rect 13412 5868 20168 5896
rect 13412 5856 13418 5868
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 25958 5856 25964 5908
rect 26016 5856 26022 5908
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 16945 5831 17003 5837
rect 16945 5828 16957 5831
rect 16632 5800 16957 5828
rect 16632 5788 16638 5800
rect 16945 5797 16957 5800
rect 16991 5797 17003 5831
rect 16945 5791 17003 5797
rect 3970 5720 3976 5772
rect 4028 5720 4034 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4387 5732 5764 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5736 5692 5764 5732
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 12768 5732 14565 5760
rect 12768 5720 12774 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 6638 5692 6644 5704
rect 5736 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 12400 5664 14289 5692
rect 12400 5652 12406 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 14976 5664 15577 5692
rect 14976 5652 14982 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5692 24639 5695
rect 24670 5692 24676 5704
rect 24627 5664 24676 5692
rect 24627 5661 24639 5664
rect 24581 5655 24639 5661
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 24848 5695 24906 5701
rect 24848 5661 24860 5695
rect 24894 5692 24906 5695
rect 25590 5692 25596 5704
rect 24894 5664 25596 5692
rect 24894 5661 24906 5664
rect 24848 5655 24906 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 15832 5627 15890 5633
rect 15832 5593 15844 5627
rect 15878 5624 15890 5627
rect 15930 5624 15936 5636
rect 15878 5596 15936 5624
rect 15878 5593 15890 5596
rect 15832 5587 15890 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 14553 5559 14611 5565
rect 14553 5556 14565 5559
rect 14332 5528 14565 5556
rect 14332 5516 14338 5528
rect 14553 5525 14565 5528
rect 14599 5525 14611 5559
rect 14553 5519 14611 5525
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 10410 5352 10416 5364
rect 9631 5324 10416 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 10502 5312 10508 5364
rect 10560 5312 10566 5364
rect 13449 5355 13507 5361
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 14918 5352 14924 5364
rect 13495 5324 14924 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 19518 5312 19524 5364
rect 19576 5312 19582 5364
rect 24670 5312 24676 5364
rect 24728 5312 24734 5364
rect 29730 5312 29736 5364
rect 29788 5312 29794 5364
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 4062 5284 4068 5296
rect 3016 5256 4068 5284
rect 3016 5244 3022 5256
rect 4062 5244 4068 5256
rect 4120 5284 4126 5296
rect 4341 5287 4399 5293
rect 4120 5256 4200 5284
rect 4120 5244 4126 5256
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 4172 5225 4200 5256
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4706 5284 4712 5296
rect 4387 5256 4712 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9493 5287 9551 5293
rect 9493 5284 9505 5287
rect 9364 5256 9505 5284
rect 9364 5244 9370 5256
rect 9493 5253 9505 5256
rect 9539 5253 9551 5287
rect 9493 5247 9551 5253
rect 14737 5287 14795 5293
rect 14737 5253 14749 5287
rect 14783 5284 14795 5287
rect 15838 5284 15844 5296
rect 14783 5256 15844 5284
rect 14783 5253 14795 5256
rect 14737 5247 14795 5253
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 18230 5244 18236 5296
rect 18288 5244 18294 5296
rect 23382 5244 23388 5296
rect 23440 5244 23446 5296
rect 28620 5287 28678 5293
rect 28620 5253 28632 5287
rect 28666 5284 28678 5287
rect 28718 5284 28724 5296
rect 28666 5256 28724 5284
rect 28666 5253 28678 5256
rect 28620 5247 28678 5253
rect 28718 5244 28724 5256
rect 28776 5244 28782 5296
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3200 5188 3985 5216
rect 3200 5176 3206 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 5810 5176 5816 5228
rect 5868 5176 5874 5228
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11054 5216 11060 5228
rect 10643 5188 11060 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 25774 5176 25780 5228
rect 25832 5176 25838 5228
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5185 26019 5219
rect 29178 5216 29184 5228
rect 25961 5179 26019 5185
rect 28368 5188 29184 5216
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6638 5148 6644 5160
rect 5951 5120 6644 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 6696 5120 9321 5148
rect 6696 5108 6702 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 13262 5108 13268 5160
rect 13320 5148 13326 5160
rect 25038 5148 25044 5160
rect 13320 5120 25044 5148
rect 13320 5108 13326 5120
rect 25038 5108 25044 5120
rect 25096 5148 25102 5160
rect 25976 5148 26004 5179
rect 26694 5148 26700 5160
rect 25096 5120 26700 5148
rect 25096 5108 25102 5120
rect 26694 5108 26700 5120
rect 26752 5108 26758 5160
rect 28368 5157 28396 5188
rect 29178 5176 29184 5188
rect 29236 5216 29242 5228
rect 29914 5216 29920 5228
rect 29236 5188 29920 5216
rect 29236 5176 29242 5188
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 28353 5151 28411 5157
rect 28353 5117 28365 5151
rect 28399 5117 28411 5151
rect 28353 5111 28411 5117
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 13262 5012 13268 5024
rect 9999 4984 13268 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 15286 4972 15292 5024
rect 15344 4972 15350 5024
rect 25593 5015 25651 5021
rect 25593 4981 25605 5015
rect 25639 5012 25651 5015
rect 25682 5012 25688 5024
rect 25639 4984 25688 5012
rect 25639 4981 25651 4984
rect 25593 4975 25651 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 11698 4808 11704 4820
rect 7208 4780 11704 4808
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 7208 4681 7236 4780
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 22462 4808 22468 4820
rect 13320 4780 22468 4808
rect 13320 4768 13326 4780
rect 22462 4768 22468 4780
rect 22520 4768 22526 4820
rect 13081 4743 13139 4749
rect 13081 4709 13093 4743
rect 13127 4740 13139 4743
rect 14366 4740 14372 4752
rect 13127 4712 14372 4740
rect 13127 4709 13139 4712
rect 13081 4703 13139 4709
rect 14366 4700 14372 4712
rect 14424 4700 14430 4752
rect 14553 4743 14611 4749
rect 14553 4709 14565 4743
rect 14599 4740 14611 4743
rect 20990 4740 20996 4752
rect 14599 4712 20996 4740
rect 14599 4709 14611 4712
rect 14553 4703 14611 4709
rect 20990 4700 20996 4712
rect 21048 4700 21054 4752
rect 24670 4700 24676 4752
rect 24728 4700 24734 4752
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 5132 4644 7205 4672
rect 5132 4632 5138 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8996 4644 9137 4672
rect 8996 4632 9002 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 9447 4644 11836 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 7466 4613 7472 4616
rect 7460 4604 7472 4613
rect 7427 4576 7472 4604
rect 7460 4567 7472 4576
rect 7466 4564 7472 4567
rect 7524 4564 7530 4616
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 11698 4564 11704 4616
rect 11756 4564 11762 4616
rect 11808 4604 11836 4644
rect 14568 4644 16221 4672
rect 14568 4616 14596 4644
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 17586 4672 17592 4684
rect 16255 4644 17592 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 17586 4632 17592 4644
rect 17644 4672 17650 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 17644 4644 18705 4672
rect 17644 4632 17650 4644
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 18739 4644 20453 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20441 4641 20453 4644
rect 20487 4672 20499 4675
rect 21174 4672 21180 4684
rect 20487 4644 21180 4672
rect 20487 4641 20499 4644
rect 20441 4635 20499 4641
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 25038 4632 25044 4684
rect 25096 4632 25102 4684
rect 11974 4613 11980 4616
rect 11968 4604 11980 4613
rect 11808 4576 11980 4604
rect 11968 4567 11980 4576
rect 11974 4564 11980 4567
rect 12032 4564 12038 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17092 4576 17417 4604
rect 17092 4564 17098 4576
rect 17405 4573 17417 4576
rect 17451 4604 17463 4607
rect 18322 4604 18328 4616
rect 17451 4576 18328 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 18414 4564 18420 4616
rect 18472 4564 18478 4616
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21637 4607 21695 4613
rect 21637 4604 21649 4607
rect 20956 4576 21649 4604
rect 20956 4564 20962 4576
rect 21637 4573 21649 4576
rect 21683 4604 21695 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21683 4576 22293 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22281 4573 22293 4576
rect 22327 4604 22339 4607
rect 24394 4604 24400 4616
rect 22327 4576 24400 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 24394 4564 24400 4576
rect 24452 4564 24458 4616
rect 25958 4564 25964 4616
rect 26016 4604 26022 4616
rect 26053 4607 26111 4613
rect 26053 4604 26065 4607
rect 26016 4576 26065 4604
rect 26016 4564 26022 4576
rect 26053 4573 26065 4576
rect 26099 4604 26111 4607
rect 27154 4604 27160 4616
rect 26099 4576 27160 4604
rect 26099 4573 26111 4576
rect 26053 4567 26111 4573
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 15933 4539 15991 4545
rect 15933 4536 15945 4539
rect 13228 4508 15945 4536
rect 13228 4496 13234 4508
rect 15933 4505 15945 4508
rect 15979 4505 15991 4539
rect 15933 4499 15991 4505
rect 26320 4539 26378 4545
rect 26320 4505 26332 4539
rect 26366 4536 26378 4539
rect 26602 4536 26608 4548
rect 26366 4508 26608 4536
rect 26366 4505 26378 4508
rect 26320 4499 26378 4505
rect 26602 4496 26608 4508
rect 26660 4496 26666 4548
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9766 4468 9772 4480
rect 8619 4440 9772 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 11054 4468 11060 4480
rect 10919 4440 11060 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 14366 4428 14372 4480
rect 14424 4428 14430 4480
rect 15562 4428 15568 4480
rect 15620 4428 15626 4480
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 16298 4468 16304 4480
rect 16071 4440 16304 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17494 4428 17500 4480
rect 17552 4428 17558 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18230 4468 18236 4480
rect 18095 4440 18236 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 19058 4468 19064 4480
rect 18555 4440 19064 4468
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19702 4428 19708 4480
rect 19760 4468 19766 4480
rect 19797 4471 19855 4477
rect 19797 4468 19809 4471
rect 19760 4440 19809 4468
rect 19760 4428 19766 4440
rect 19797 4437 19809 4440
rect 19843 4437 19855 4471
rect 19797 4431 19855 4437
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20622 4468 20628 4480
rect 20303 4440 20628 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21542 4428 21548 4480
rect 21600 4428 21606 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22189 4471 22247 4477
rect 22189 4468 22201 4471
rect 22152 4440 22201 4468
rect 22152 4428 22158 4440
rect 22189 4437 22201 4440
rect 22235 4437 22247 4471
rect 22189 4431 22247 4437
rect 24578 4428 24584 4480
rect 24636 4428 24642 4480
rect 26786 4428 26792 4480
rect 26844 4468 26850 4480
rect 27433 4471 27491 4477
rect 27433 4468 27445 4471
rect 26844 4440 27445 4468
rect 26844 4428 26850 4440
rect 27433 4437 27445 4440
rect 27479 4437 27491 4471
rect 27433 4431 27491 4437
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8168 4236 9260 4264
rect 8168 4224 8174 4236
rect 7377 4199 7435 4205
rect 7377 4165 7389 4199
rect 7423 4196 7435 4199
rect 7466 4196 7472 4208
rect 7423 4168 7472 4196
rect 7423 4165 7435 4168
rect 7377 4159 7435 4165
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 7926 4156 7932 4208
rect 7984 4156 7990 4208
rect 9232 4196 9260 4236
rect 9306 4224 9312 4276
rect 9364 4224 9370 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10410 4264 10416 4276
rect 9732 4236 10416 4264
rect 9732 4224 9738 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 26145 4267 26203 4273
rect 26145 4233 26157 4267
rect 26191 4264 26203 4267
rect 26602 4264 26608 4276
rect 26191 4236 26608 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26602 4224 26608 4236
rect 26660 4224 26666 4276
rect 13357 4199 13415 4205
rect 13357 4196 13369 4199
rect 9232 4168 13369 4196
rect 13357 4165 13369 4168
rect 13403 4165 13415 4199
rect 15286 4196 15292 4208
rect 13357 4159 13415 4165
rect 15120 4168 15292 4196
rect 8938 4128 8944 4140
rect 8588 4100 8944 4128
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4060 7159 4063
rect 8588 4060 8616 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 7147 4032 8616 4060
rect 8849 4063 8907 4069
rect 7147 4029 7159 4032
rect 7101 4023 7159 4029
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9674 4060 9680 4072
rect 8895 4032 9680 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 9876 3924 9904 4023
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10796 4060 10824 4091
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11112 4100 11897 4128
rect 11112 4088 11118 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13998 4128 14004 4140
rect 13495 4100 14004 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15120 4128 15148 4168
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 17948 4199 18006 4205
rect 17948 4165 17960 4199
rect 17994 4196 18006 4199
rect 18230 4196 18236 4208
rect 17994 4168 18236 4196
rect 17994 4165 18006 4168
rect 17948 4159 18006 4165
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 24394 4156 24400 4208
rect 24452 4196 24458 4208
rect 25958 4196 25964 4208
rect 24452 4168 25964 4196
rect 24452 4156 24458 4168
rect 25958 4156 25964 4168
rect 26016 4156 26022 4208
rect 14967 4100 15148 4128
rect 15188 4131 15246 4137
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15188 4097 15200 4131
rect 15234 4128 15246 4131
rect 15562 4128 15568 4140
rect 15234 4100 15568 4128
rect 15234 4097 15246 4100
rect 15188 4091 15246 4097
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17552 4100 17693 4128
rect 17552 4088 17558 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21186 4131 21244 4137
rect 21186 4128 21198 4131
rect 20772 4100 21198 4128
rect 20772 4088 20778 4100
rect 21186 4097 21198 4100
rect 21232 4097 21244 4131
rect 21186 4091 21244 4097
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 21542 4128 21548 4140
rect 21499 4100 21548 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22278 4137 22284 4140
rect 22272 4091 22284 4137
rect 22278 4088 22284 4091
rect 22336 4088 22342 4140
rect 10008 4032 10824 4060
rect 13633 4063 13691 4069
rect 10008 4020 10014 4032
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14182 4060 14188 4072
rect 13679 4032 14188 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14182 4020 14188 4032
rect 14240 4060 14246 4072
rect 14550 4060 14556 4072
rect 14240 4032 14556 4060
rect 14240 4020 14246 4032
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4060 24363 4063
rect 24412 4060 24440 4156
rect 24578 4137 24584 4140
rect 24572 4128 24584 4137
rect 24539 4100 24584 4128
rect 24572 4091 24584 4100
rect 24578 4088 24584 4091
rect 24636 4088 24642 4140
rect 27154 4088 27160 4140
rect 27212 4088 27218 4140
rect 27430 4137 27436 4140
rect 27424 4091 27436 4137
rect 27430 4088 27436 4091
rect 27488 4088 27494 4140
rect 24351 4032 24440 4060
rect 26605 4063 26663 4069
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 26605 4029 26617 4063
rect 26651 4060 26663 4063
rect 26694 4060 26700 4072
rect 26651 4032 26700 4060
rect 26651 4029 26663 4032
rect 26605 4023 26663 4029
rect 26694 4020 26700 4032
rect 26752 4020 26758 4072
rect 12437 3995 12495 4001
rect 12437 3961 12449 3995
rect 12483 3992 12495 3995
rect 14366 3992 14372 4004
rect 12483 3964 14372 3992
rect 12483 3961 12495 3964
rect 12437 3955 12495 3961
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 26237 3995 26295 4001
rect 26237 3961 26249 3995
rect 26283 3992 26295 3995
rect 26283 3964 26317 3992
rect 26283 3961 26295 3964
rect 26237 3955 26295 3961
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 9876 3896 11989 3924
rect 11977 3893 11989 3896
rect 12023 3924 12035 3927
rect 12710 3924 12716 3936
rect 12023 3896 12716 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 16298 3884 16304 3936
rect 16356 3884 16362 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16724 3896 16957 3924
rect 16724 3884 16730 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 19058 3884 19064 3936
rect 19116 3884 19122 3936
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 21082 3924 21088 3936
rect 20119 3896 21088 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 23382 3884 23388 3936
rect 23440 3884 23446 3936
rect 25685 3927 25743 3933
rect 25685 3893 25697 3927
rect 25731 3924 25743 3927
rect 26252 3924 26280 3955
rect 26602 3924 26608 3936
rect 25731 3896 26608 3924
rect 25731 3893 25743 3896
rect 25685 3887 25743 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 28350 3884 28356 3936
rect 28408 3924 28414 3936
rect 28537 3927 28595 3933
rect 28537 3924 28549 3927
rect 28408 3896 28549 3924
rect 28408 3884 28414 3896
rect 28537 3893 28549 3896
rect 28583 3893 28595 3927
rect 28537 3887 28595 3893
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 7926 3680 7932 3732
rect 7984 3680 7990 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 20809 3723 20867 3729
rect 20809 3720 20821 3723
rect 20680 3692 20821 3720
rect 20680 3680 20686 3692
rect 20809 3689 20821 3692
rect 20855 3689 20867 3723
rect 20809 3683 20867 3689
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22370 3720 22376 3732
rect 22143 3692 22376 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 24581 3723 24639 3729
rect 24581 3689 24593 3723
rect 24627 3720 24639 3723
rect 24670 3720 24676 3732
rect 24627 3692 24676 3720
rect 24627 3689 24639 3692
rect 24581 3683 24639 3689
rect 24670 3680 24676 3692
rect 24728 3720 24734 3732
rect 25038 3720 25044 3732
rect 24728 3692 25044 3720
rect 24728 3680 24734 3692
rect 25038 3680 25044 3692
rect 25096 3720 25102 3732
rect 25096 3692 26188 3720
rect 25096 3680 25102 3692
rect 9950 3584 9956 3596
rect 7944 3556 9956 3584
rect 7944 3525 7972 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 16666 3544 16672 3596
rect 16724 3544 16730 3596
rect 22738 3544 22744 3596
rect 22796 3544 22802 3596
rect 25958 3544 25964 3596
rect 26016 3544 26022 3596
rect 26160 3584 26188 3692
rect 26786 3680 26792 3732
rect 26844 3680 26850 3732
rect 26234 3612 26240 3664
rect 26292 3652 26298 3664
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26292 3624 26893 3652
rect 26292 3612 26298 3624
rect 26881 3621 26893 3624
rect 26927 3652 26939 3655
rect 28350 3652 28356 3664
rect 26927 3624 28356 3652
rect 26927 3621 26939 3624
rect 26881 3615 26939 3621
rect 28350 3612 28356 3624
rect 28408 3612 28414 3664
rect 26973 3587 27031 3593
rect 26973 3584 26985 3587
rect 26160 3556 26985 3584
rect 26973 3553 26985 3556
rect 27019 3553 27031 3587
rect 26973 3547 27031 3553
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 12342 3476 12348 3528
rect 12400 3476 12406 3528
rect 12612 3519 12670 3525
rect 12612 3485 12624 3519
rect 12658 3516 12670 3519
rect 12986 3516 12992 3528
rect 12658 3488 12992 3516
rect 12658 3485 12670 3488
rect 12612 3479 12670 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 19702 3525 19708 3528
rect 19696 3516 19708 3525
rect 19663 3488 19708 3516
rect 19696 3479 19708 3488
rect 19702 3476 19708 3479
rect 19760 3476 19766 3528
rect 22462 3476 22468 3528
rect 22520 3476 22526 3528
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 23382 3516 23388 3528
rect 22603 3488 23388 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 25682 3476 25688 3528
rect 25740 3525 25746 3528
rect 25740 3516 25752 3525
rect 26421 3519 26479 3525
rect 25740 3488 25785 3516
rect 25740 3479 25752 3488
rect 26421 3485 26433 3519
rect 26467 3516 26479 3519
rect 26602 3516 26608 3528
rect 26467 3488 26608 3516
rect 26467 3485 26479 3488
rect 26421 3479 26479 3485
rect 25740 3476 25746 3479
rect 26602 3476 26608 3488
rect 26660 3476 26666 3528
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 16942 3457 16948 3460
rect 15390 3451 15448 3457
rect 15390 3448 15402 3451
rect 14792 3420 15402 3448
rect 14792 3408 14798 3420
rect 15390 3417 15402 3420
rect 15436 3417 15448 3451
rect 15390 3411 15448 3417
rect 16936 3411 16948 3457
rect 16942 3408 16948 3411
rect 17000 3408 17006 3460
rect 27341 3451 27399 3457
rect 27341 3448 27353 3451
rect 17052 3420 18368 3448
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 13998 3380 14004 3392
rect 13771 3352 14004 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 14274 3340 14280 3392
rect 14332 3340 14338 3392
rect 16850 3340 16856 3392
rect 16908 3380 16914 3392
rect 17052 3380 17080 3420
rect 16908 3352 17080 3380
rect 18049 3383 18107 3389
rect 16908 3340 16914 3352
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18230 3380 18236 3392
rect 18095 3352 18236 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 18340 3380 18368 3420
rect 22066 3420 27353 3448
rect 22066 3380 22094 3420
rect 27341 3417 27353 3420
rect 27387 3417 27399 3451
rect 27341 3411 27399 3417
rect 18340 3352 22094 3380
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12400 3148 12541 3176
rect 12400 3136 12406 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 14734 3136 14740 3188
rect 14792 3136 14798 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15654 3176 15660 3188
rect 15335 3148 15660 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18230 3176 18236 3188
rect 17451 3148 18236 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19484 3148 19625 3176
rect 19484 3136 19490 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 20714 3136 20720 3188
rect 20772 3136 20778 3188
rect 21082 3136 21088 3188
rect 21140 3136 21146 3188
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 27488 3148 27629 3176
rect 27488 3136 27494 3148
rect 27617 3145 27629 3148
rect 27663 3145 27675 3179
rect 27617 3139 27675 3145
rect 29914 3136 29920 3188
rect 29972 3136 29978 3188
rect 12636 3080 14504 3108
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 12636 3049 12664 3080
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 10008 3012 12633 3040
rect 10008 3000 10014 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 14476 3040 14504 3080
rect 26694 3068 26700 3120
rect 26752 3108 26758 3120
rect 27157 3111 27215 3117
rect 27157 3108 27169 3111
rect 26752 3080 27169 3108
rect 26752 3068 26758 3080
rect 27157 3077 27169 3080
rect 27203 3077 27215 3111
rect 27157 3071 27215 3077
rect 28629 3111 28687 3117
rect 28629 3077 28641 3111
rect 28675 3108 28687 3111
rect 28810 3108 28816 3120
rect 28675 3080 28816 3108
rect 28675 3077 28687 3080
rect 28629 3071 28687 3077
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 15194 3040 15200 3052
rect 14476 3012 15200 3040
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 16546 3012 17325 3040
rect 14182 2932 14188 2984
rect 14240 2932 14246 2984
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 15470 2972 15476 2984
rect 14332 2944 15476 2972
rect 14332 2932 14338 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 16546 2904 16574 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20806 3040 20812 3052
rect 19751 3012 20812 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3040 20959 3043
rect 20990 3040 20996 3052
rect 20947 3012 20996 3040
rect 20947 3009 20959 3012
rect 20901 3003 20959 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21174 3000 21180 3052
rect 21232 3040 21238 3052
rect 22738 3040 22744 3052
rect 21232 3012 22744 3040
rect 21232 3000 21238 3012
rect 22738 3000 22744 3012
rect 22796 3040 22802 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 22796 3012 25145 3040
rect 22796 3000 22802 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 17586 2932 17592 2984
rect 17644 2932 17650 2984
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 25096 2944 25513 2972
rect 25096 2932 25102 2944
rect 25501 2941 25513 2944
rect 25547 2941 25559 2975
rect 25501 2935 25559 2941
rect 11020 2876 16574 2904
rect 25593 2907 25651 2913
rect 11020 2864 11026 2876
rect 25593 2873 25605 2907
rect 25639 2904 25651 2907
rect 26053 2907 26111 2913
rect 25639 2876 26004 2904
rect 25639 2873 25651 2876
rect 25593 2867 25651 2873
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2836 25743 2839
rect 25774 2836 25780 2848
rect 25731 2808 25780 2836
rect 25731 2805 25743 2808
rect 25685 2799 25743 2805
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 25976 2836 26004 2876
rect 26053 2873 26065 2907
rect 26099 2904 26111 2907
rect 26786 2904 26792 2916
rect 26099 2876 26792 2904
rect 26099 2873 26111 2876
rect 26053 2867 26111 2873
rect 26786 2864 26792 2876
rect 26844 2904 26850 2916
rect 27433 2907 27491 2913
rect 27433 2904 27445 2907
rect 26844 2876 27445 2904
rect 26844 2864 26850 2876
rect 27172 2848 27200 2876
rect 27433 2873 27445 2876
rect 27479 2873 27491 2907
rect 27433 2867 27491 2873
rect 26234 2836 26240 2848
rect 25976 2808 26240 2836
rect 26234 2796 26240 2808
rect 26292 2836 26298 2848
rect 26602 2836 26608 2848
rect 26292 2808 26608 2836
rect 26292 2796 26298 2808
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27154 2796 27160 2848
rect 27212 2796 27218 2848
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 14366 2632 14372 2644
rect 3068 2604 14372 2632
rect 3068 2437 3096 2604
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 10134 2564 10140 2576
rect 5644 2536 10140 2564
rect 5644 2437 5672 2536
rect 10134 2524 10140 2536
rect 10192 2564 10198 2576
rect 10962 2564 10968 2576
rect 10192 2536 10968 2564
rect 10192 2524 10198 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 18230 2456 18236 2508
rect 18288 2456 18294 2508
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 5629 2431 5687 2437
rect 4479 2400 5580 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1268 2332 1777 2360
rect 1268 2320 1274 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2056 2292 2084 2391
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2556 2332 2789 2360
rect 2556 2320 2562 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 4154 2320 4160 2372
rect 4212 2320 4218 2372
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5132 2332 5365 2360
rect 5132 2320 5138 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5552 2360 5580 2400
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7650 2388 7656 2440
rect 7708 2428 7714 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7708 2400 7757 2428
rect 7708 2388 7714 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8996 2400 9137 2428
rect 8996 2388 9002 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10284 2400 10333 2428
rect 10284 2388 10290 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11572 2400 11713 2428
rect 11572 2388 11578 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12860 2400 12909 2428
rect 12860 2388 12866 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 18248 2428 18276 2456
rect 18095 2400 18276 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19116 2400 19441 2428
rect 19116 2388 19122 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20622 2388 20628 2440
rect 20680 2388 20686 2440
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21140 2400 22017 2428
rect 21140 2388 21146 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23382 2428 23388 2440
rect 23247 2400 23388 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 25038 2388 25044 2440
rect 25096 2388 25102 2440
rect 26234 2388 26240 2440
rect 26292 2388 26298 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 28350 2388 28356 2440
rect 28408 2388 28414 2440
rect 29546 2388 29552 2440
rect 29604 2428 29610 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29604 2400 29745 2428
rect 29604 2388 29610 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30892 2400 30941 2428
rect 30892 2388 30898 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 32122 2388 32128 2440
rect 32180 2428 32186 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32180 2400 32321 2428
rect 32180 2388 32186 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33505 2431 33563 2437
rect 33505 2428 33517 2431
rect 33468 2400 33517 2428
rect 33468 2388 33474 2400
rect 33505 2397 33517 2400
rect 33551 2397 33563 2431
rect 33505 2391 33563 2397
rect 13170 2360 13176 2372
rect 5552 2332 13176 2360
rect 5353 2323 5411 2329
rect 13170 2320 13176 2332
rect 13228 2320 13234 2372
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14148 2332 14565 2360
rect 14148 2320 14154 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15436 2332 15761 2360
rect 15436 2320 15442 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16724 2332 17141 2360
rect 16724 2320 16730 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18288 2332 18337 2360
rect 18288 2320 18294 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19392 2332 19717 2360
rect 19392 2320 19398 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 20901 2363 20959 2369
rect 20901 2360 20913 2363
rect 20772 2332 20913 2360
rect 20772 2320 20778 2332
rect 20901 2329 20913 2332
rect 20947 2329 20959 2363
rect 20901 2323 20959 2329
rect 22094 2320 22100 2372
rect 22152 2360 22158 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 22152 2332 22293 2360
rect 22152 2320 22158 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 23474 2320 23480 2372
rect 23532 2320 23538 2372
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24765 2363 24823 2369
rect 24765 2360 24777 2363
rect 24452 2332 24777 2360
rect 24452 2320 24458 2332
rect 24765 2329 24777 2332
rect 24811 2329 24823 2363
rect 24765 2323 24823 2329
rect 25682 2320 25688 2372
rect 25740 2360 25746 2372
rect 25961 2363 26019 2369
rect 25961 2360 25973 2363
rect 25740 2332 25973 2360
rect 25740 2320 25746 2332
rect 25961 2329 25973 2332
rect 26007 2329 26019 2363
rect 25961 2323 26019 2329
rect 26970 2320 26976 2372
rect 27028 2360 27034 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27028 2332 27445 2360
rect 27028 2320 27034 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28258 2320 28264 2372
rect 28316 2360 28322 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28316 2332 28641 2360
rect 28316 2320 28322 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 8110 2292 8116 2304
rect 2056 2264 8116 2292
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 34333 2295 34391 2301
rect 34333 2261 34345 2295
rect 34379 2292 34391 2295
rect 34606 2292 34612 2304
rect 34379 2264 34612 2292
rect 34379 2261 34391 2264
rect 34333 2255 34391 2261
rect 34606 2252 34612 2264
rect 34664 2252 34670 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
<< via1 >>
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 4896 33575 4948 33584
rect 4896 33541 4905 33575
rect 4905 33541 4939 33575
rect 4939 33541 4948 33575
rect 4896 33532 4948 33541
rect 7840 33575 7892 33584
rect 7840 33541 7849 33575
rect 7849 33541 7883 33575
rect 7883 33541 7892 33575
rect 7840 33532 7892 33541
rect 10600 33532 10652 33584
rect 13820 33532 13872 33584
rect 16580 33532 16632 33584
rect 19432 33532 19484 33584
rect 22376 33532 22428 33584
rect 25596 33575 25648 33584
rect 25596 33541 25605 33575
rect 25605 33541 25639 33575
rect 25639 33541 25648 33575
rect 25596 33532 25648 33541
rect 28540 33575 28592 33584
rect 28540 33541 28549 33575
rect 28549 33541 28583 33575
rect 28583 33541 28592 33575
rect 28540 33532 28592 33541
rect 31484 33575 31536 33584
rect 31484 33541 31493 33575
rect 31493 33541 31527 33575
rect 31527 33541 31536 33575
rect 31484 33532 31536 33541
rect 34244 33575 34296 33584
rect 34244 33541 34253 33575
rect 34253 33541 34287 33575
rect 34287 33541 34296 33575
rect 34244 33532 34296 33541
rect 12256 33328 12308 33380
rect 14280 33371 14332 33380
rect 14280 33337 14289 33371
rect 14289 33337 14323 33371
rect 14323 33337 14332 33371
rect 14280 33328 14332 33337
rect 16856 33371 16908 33380
rect 16856 33337 16865 33371
rect 16865 33337 16899 33371
rect 16899 33337 16908 33371
rect 16856 33328 16908 33337
rect 19524 33371 19576 33380
rect 19524 33337 19533 33371
rect 19533 33337 19567 33371
rect 19567 33337 19576 33371
rect 19524 33328 19576 33337
rect 22468 33371 22520 33380
rect 22468 33337 22477 33371
rect 22477 33337 22511 33371
rect 22511 33337 22520 33371
rect 22468 33328 22520 33337
rect 25412 33371 25464 33380
rect 25412 33337 25421 33371
rect 25421 33337 25455 33371
rect 25455 33337 25464 33371
rect 25412 33328 25464 33337
rect 28356 33371 28408 33380
rect 28356 33337 28365 33371
rect 28365 33337 28399 33371
rect 28399 33337 28408 33371
rect 28356 33328 28408 33337
rect 31300 33371 31352 33380
rect 31300 33337 31309 33371
rect 31309 33337 31343 33371
rect 31343 33337 31352 33371
rect 31300 33328 31352 33337
rect 33324 33328 33376 33380
rect 4988 33303 5040 33312
rect 4988 33269 4997 33303
rect 4997 33269 5031 33303
rect 5031 33269 5040 33303
rect 4988 33260 5040 33269
rect 11612 33260 11664 33312
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 10508 32852 10560 32904
rect 16856 32920 16908 32972
rect 28356 33056 28408 33108
rect 20628 32963 20680 32972
rect 20628 32929 20637 32963
rect 20637 32929 20671 32963
rect 20671 32929 20680 32963
rect 20628 32920 20680 32929
rect 24768 32920 24820 32972
rect 15476 32784 15528 32836
rect 16764 32784 16816 32836
rect 18328 32784 18380 32836
rect 22836 32852 22888 32904
rect 10140 32759 10192 32768
rect 10140 32725 10149 32759
rect 10149 32725 10183 32759
rect 10183 32725 10192 32759
rect 10140 32716 10192 32725
rect 13268 32716 13320 32768
rect 25412 32784 25464 32836
rect 21272 32716 21324 32768
rect 22008 32716 22060 32768
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 12256 32555 12308 32564
rect 12256 32521 12265 32555
rect 12265 32521 12299 32555
rect 12299 32521 12308 32555
rect 12256 32512 12308 32521
rect 11796 32444 11848 32496
rect 13268 32487 13320 32496
rect 13268 32453 13277 32487
rect 13277 32453 13311 32487
rect 13311 32453 13320 32487
rect 13268 32444 13320 32453
rect 14280 32512 14332 32564
rect 16764 32512 16816 32564
rect 22468 32512 22520 32564
rect 10416 32419 10468 32428
rect 10416 32385 10425 32419
rect 10425 32385 10459 32419
rect 10459 32385 10468 32419
rect 10416 32376 10468 32385
rect 10508 32419 10560 32428
rect 10508 32385 10517 32419
rect 10517 32385 10551 32419
rect 10551 32385 10560 32419
rect 10508 32376 10560 32385
rect 15936 32376 15988 32428
rect 16856 32376 16908 32428
rect 17868 32376 17920 32428
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 8576 32240 8628 32292
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22652 32376 22704 32428
rect 23388 32444 23440 32496
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 24584 32376 24636 32428
rect 24768 32376 24820 32428
rect 27712 32419 27764 32428
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 27712 32376 27764 32385
rect 28080 32419 28132 32428
rect 28080 32385 28089 32419
rect 28089 32385 28123 32419
rect 28123 32385 28132 32419
rect 28080 32376 28132 32385
rect 31300 32376 31352 32428
rect 33324 32419 33376 32428
rect 33324 32385 33333 32419
rect 33333 32385 33367 32419
rect 33367 32385 33376 32419
rect 33324 32376 33376 32385
rect 21272 32351 21324 32360
rect 21272 32317 21281 32351
rect 21281 32317 21315 32351
rect 21315 32317 21324 32351
rect 21272 32308 21324 32317
rect 22836 32308 22888 32360
rect 21088 32240 21140 32292
rect 10048 32172 10100 32224
rect 10600 32215 10652 32224
rect 10600 32181 10609 32215
rect 10609 32181 10643 32215
rect 10643 32181 10652 32215
rect 10600 32172 10652 32181
rect 11888 32172 11940 32224
rect 13176 32172 13228 32224
rect 13360 32172 13412 32224
rect 19524 32172 19576 32224
rect 25044 32172 25096 32224
rect 30196 32172 30248 32224
rect 33140 32215 33192 32224
rect 33140 32181 33149 32215
rect 33149 32181 33183 32215
rect 33183 32181 33192 32215
rect 33140 32172 33192 32181
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 15844 31968 15896 32020
rect 15936 32011 15988 32020
rect 15936 31977 15945 32011
rect 15945 31977 15979 32011
rect 15979 31977 15988 32011
rect 15936 31968 15988 31977
rect 18236 31968 18288 32020
rect 20628 31968 20680 32020
rect 23204 31968 23256 32020
rect 8760 31900 8812 31952
rect 11704 31900 11756 31952
rect 9864 31875 9916 31884
rect 9864 31841 9873 31875
rect 9873 31841 9907 31875
rect 9907 31841 9916 31875
rect 9864 31832 9916 31841
rect 13360 31832 13412 31884
rect 8576 31807 8628 31816
rect 8576 31773 8585 31807
rect 8585 31773 8619 31807
rect 8619 31773 8628 31807
rect 8576 31764 8628 31773
rect 10140 31764 10192 31816
rect 10508 31764 10560 31816
rect 15660 31900 15712 31952
rect 17132 31875 17184 31884
rect 17132 31841 17141 31875
rect 17141 31841 17175 31875
rect 17175 31841 17184 31875
rect 17132 31832 17184 31841
rect 20536 31900 20588 31952
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 14648 31764 14700 31816
rect 11612 31739 11664 31748
rect 11612 31705 11621 31739
rect 11621 31705 11655 31739
rect 11655 31705 11664 31739
rect 11612 31696 11664 31705
rect 11796 31696 11848 31748
rect 10048 31628 10100 31680
rect 15752 31671 15804 31680
rect 15752 31637 15777 31671
rect 15777 31637 15804 31671
rect 15936 31696 15988 31748
rect 17316 31807 17368 31816
rect 17316 31773 17325 31807
rect 17325 31773 17359 31807
rect 17359 31773 17368 31807
rect 17316 31764 17368 31773
rect 17868 31764 17920 31816
rect 21088 31832 21140 31884
rect 22652 31900 22704 31952
rect 15752 31628 15804 31637
rect 16672 31628 16724 31680
rect 18328 31628 18380 31680
rect 20812 31764 20864 31816
rect 21180 31764 21232 31816
rect 21364 31764 21416 31816
rect 22928 31832 22980 31884
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 25136 31875 25188 31884
rect 25136 31841 25145 31875
rect 25145 31841 25179 31875
rect 25179 31841 25188 31875
rect 25136 31832 25188 31841
rect 21088 31739 21140 31748
rect 21088 31705 21097 31739
rect 21097 31705 21131 31739
rect 21131 31705 21140 31739
rect 21088 31696 21140 31705
rect 22836 31807 22888 31816
rect 22836 31773 22845 31807
rect 22845 31773 22879 31807
rect 22879 31773 22888 31807
rect 22836 31764 22888 31773
rect 23756 31807 23808 31816
rect 23756 31773 23765 31807
rect 23765 31773 23799 31807
rect 23799 31773 23808 31807
rect 23756 31764 23808 31773
rect 23388 31696 23440 31748
rect 26608 31807 26660 31816
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 26700 31696 26752 31748
rect 27712 31696 27764 31748
rect 23480 31671 23532 31680
rect 23480 31637 23489 31671
rect 23489 31637 23523 31671
rect 23523 31637 23532 31671
rect 23480 31628 23532 31637
rect 24768 31628 24820 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 9864 31424 9916 31476
rect 14280 31424 14332 31476
rect 15844 31424 15896 31476
rect 17316 31424 17368 31476
rect 20812 31467 20864 31476
rect 20812 31433 20846 31467
rect 20846 31433 20864 31467
rect 20812 31424 20864 31433
rect 25136 31424 25188 31476
rect 26608 31424 26660 31476
rect 27344 31424 27396 31476
rect 10048 31356 10100 31408
rect 10600 31356 10652 31408
rect 8852 31288 8904 31340
rect 9956 31288 10008 31340
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 12716 31288 12768 31340
rect 15660 31356 15712 31408
rect 16028 31356 16080 31408
rect 14096 31331 14148 31340
rect 14096 31297 14105 31331
rect 14105 31297 14139 31331
rect 14139 31297 14148 31331
rect 14096 31288 14148 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 9404 31220 9456 31272
rect 9496 31220 9548 31272
rect 12440 31220 12492 31272
rect 13268 31263 13320 31272
rect 13268 31229 13277 31263
rect 13277 31229 13311 31263
rect 13311 31229 13320 31263
rect 13268 31220 13320 31229
rect 14648 31220 14700 31272
rect 15568 31288 15620 31340
rect 16672 31356 16724 31408
rect 17132 31331 17184 31340
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 17684 31288 17736 31340
rect 20352 31288 20404 31340
rect 24492 31356 24544 31408
rect 24676 31356 24728 31408
rect 20996 31288 21048 31340
rect 22652 31331 22704 31340
rect 22652 31297 22661 31331
rect 22661 31297 22695 31331
rect 22695 31297 22704 31331
rect 22652 31288 22704 31297
rect 22928 31331 22980 31340
rect 22928 31297 22937 31331
rect 22937 31297 22971 31331
rect 22971 31297 22980 31331
rect 22928 31288 22980 31297
rect 23020 31331 23072 31340
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 15752 31220 15804 31272
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 21364 31220 21416 31272
rect 21456 31220 21508 31272
rect 23480 31331 23532 31340
rect 23480 31297 23489 31331
rect 23489 31297 23523 31331
rect 23523 31297 23532 31331
rect 23480 31288 23532 31297
rect 24584 31288 24636 31340
rect 24860 31288 24912 31340
rect 25320 31288 25372 31340
rect 25688 31331 25740 31340
rect 25688 31297 25697 31331
rect 25697 31297 25731 31331
rect 25731 31297 25740 31331
rect 25688 31288 25740 31297
rect 26700 31288 26752 31340
rect 27344 31331 27396 31340
rect 27344 31297 27353 31331
rect 27353 31297 27387 31331
rect 27387 31297 27396 31331
rect 27344 31288 27396 31297
rect 25596 31263 25648 31272
rect 25596 31229 25605 31263
rect 25605 31229 25639 31263
rect 25639 31229 25648 31263
rect 25596 31220 25648 31229
rect 29092 31263 29144 31272
rect 29092 31229 29101 31263
rect 29101 31229 29135 31263
rect 29135 31229 29144 31263
rect 29092 31220 29144 31229
rect 10692 31152 10744 31204
rect 16856 31195 16908 31204
rect 16856 31161 16865 31195
rect 16865 31161 16899 31195
rect 16899 31161 16908 31195
rect 16856 31152 16908 31161
rect 14280 31127 14332 31136
rect 14280 31093 14289 31127
rect 14289 31093 14323 31127
rect 14323 31093 14332 31127
rect 14280 31084 14332 31093
rect 25780 31084 25832 31136
rect 29000 31127 29052 31136
rect 29000 31093 29009 31127
rect 29009 31093 29043 31127
rect 29043 31093 29052 31127
rect 29000 31084 29052 31093
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 9404 30923 9456 30932
rect 9404 30889 9413 30923
rect 9413 30889 9447 30923
rect 9447 30889 9456 30923
rect 9404 30880 9456 30889
rect 10048 30923 10100 30932
rect 10048 30889 10057 30923
rect 10057 30889 10091 30923
rect 10091 30889 10100 30923
rect 10048 30880 10100 30889
rect 10232 30880 10284 30932
rect 13268 30880 13320 30932
rect 20996 30923 21048 30932
rect 20996 30889 21005 30923
rect 21005 30889 21039 30923
rect 21039 30889 21048 30923
rect 20996 30880 21048 30889
rect 23020 30880 23072 30932
rect 10508 30744 10560 30796
rect 14832 30812 14884 30864
rect 9496 30719 9548 30728
rect 9496 30685 9505 30719
rect 9505 30685 9539 30719
rect 9539 30685 9548 30719
rect 9496 30676 9548 30685
rect 9956 30719 10008 30728
rect 9956 30685 9965 30719
rect 9965 30685 9999 30719
rect 9999 30685 10008 30719
rect 9956 30676 10008 30685
rect 10140 30719 10192 30728
rect 10140 30685 10149 30719
rect 10149 30685 10183 30719
rect 10183 30685 10192 30719
rect 10140 30676 10192 30685
rect 10416 30676 10468 30728
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 10600 30676 10652 30685
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 14096 30676 14148 30728
rect 14556 30676 14608 30728
rect 14924 30676 14976 30728
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 16028 30719 16080 30728
rect 16028 30685 16037 30719
rect 16037 30685 16071 30719
rect 16071 30685 16080 30719
rect 16028 30676 16080 30685
rect 23388 30812 23440 30864
rect 23756 30744 23808 30796
rect 24676 30744 24728 30796
rect 25228 30744 25280 30796
rect 21456 30676 21508 30728
rect 22928 30719 22980 30728
rect 22928 30685 22937 30719
rect 22937 30685 22971 30719
rect 22971 30685 22980 30719
rect 22928 30676 22980 30685
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 25044 30719 25096 30728
rect 25044 30685 25053 30719
rect 25053 30685 25087 30719
rect 25087 30685 25096 30719
rect 25044 30676 25096 30685
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 25780 30719 25832 30728
rect 25780 30685 25789 30719
rect 25789 30685 25823 30719
rect 25823 30685 25832 30719
rect 25780 30676 25832 30685
rect 29092 30744 29144 30796
rect 27712 30719 27764 30728
rect 27712 30685 27721 30719
rect 27721 30685 27755 30719
rect 27755 30685 27764 30719
rect 27712 30676 27764 30685
rect 17592 30608 17644 30660
rect 20996 30608 21048 30660
rect 26148 30651 26200 30660
rect 26148 30617 26157 30651
rect 26157 30617 26191 30651
rect 26191 30617 26200 30651
rect 26148 30608 26200 30617
rect 27620 30608 27672 30660
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 28724 30608 28776 30660
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 29000 30336 29052 30388
rect 29092 30336 29144 30388
rect 16028 30268 16080 30320
rect 25044 30268 25096 30320
rect 25688 30268 25740 30320
rect 14280 30243 14332 30252
rect 14280 30209 14289 30243
rect 14289 30209 14323 30243
rect 14323 30209 14332 30243
rect 14280 30200 14332 30209
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 20168 30200 20220 30252
rect 20812 30200 20864 30252
rect 20904 30200 20956 30252
rect 24676 30243 24728 30252
rect 24676 30209 24685 30243
rect 24685 30209 24719 30243
rect 24719 30209 24728 30243
rect 24676 30200 24728 30209
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 25228 30200 25280 30252
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 27712 30268 27764 30320
rect 28080 30311 28132 30320
rect 28080 30277 28089 30311
rect 28089 30277 28123 30311
rect 28123 30277 28132 30311
rect 28080 30268 28132 30277
rect 25596 30132 25648 30184
rect 27528 30200 27580 30252
rect 28448 30200 28500 30252
rect 26148 30132 26200 30184
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 29000 30243 29052 30252
rect 29000 30209 29009 30243
rect 29009 30209 29043 30243
rect 29043 30209 29052 30243
rect 29000 30200 29052 30209
rect 29184 30243 29236 30252
rect 29184 30209 29193 30243
rect 29193 30209 29227 30243
rect 29227 30209 29236 30243
rect 29184 30200 29236 30209
rect 29644 30243 29696 30252
rect 29644 30209 29653 30243
rect 29653 30209 29687 30243
rect 29687 30209 29696 30243
rect 29644 30200 29696 30209
rect 25780 30064 25832 30116
rect 28080 30064 28132 30116
rect 12900 29996 12952 30048
rect 20628 29996 20680 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 25044 29835 25096 29844
rect 25044 29801 25053 29835
rect 25053 29801 25087 29835
rect 25087 29801 25096 29835
rect 25044 29792 25096 29801
rect 25136 29792 25188 29844
rect 9036 29724 9088 29776
rect 10692 29656 10744 29708
rect 10416 29631 10468 29640
rect 10416 29597 10425 29631
rect 10425 29597 10459 29631
rect 10459 29597 10468 29631
rect 10416 29588 10468 29597
rect 10140 29520 10192 29572
rect 12900 29588 12952 29640
rect 10692 29563 10744 29572
rect 10692 29529 10701 29563
rect 10701 29529 10735 29563
rect 10735 29529 10744 29563
rect 10692 29520 10744 29529
rect 15016 29588 15068 29640
rect 19616 29631 19668 29640
rect 19616 29597 19625 29631
rect 19625 29597 19659 29631
rect 19659 29597 19668 29631
rect 20536 29656 20588 29708
rect 20812 29656 20864 29708
rect 23204 29724 23256 29776
rect 27712 29767 27764 29776
rect 27712 29733 27721 29767
rect 27721 29733 27755 29767
rect 27755 29733 27764 29767
rect 27712 29724 27764 29733
rect 27160 29656 27212 29708
rect 19616 29588 19668 29597
rect 20352 29588 20404 29640
rect 20720 29588 20772 29640
rect 14188 29520 14240 29572
rect 15108 29563 15160 29572
rect 15108 29529 15117 29563
rect 15117 29529 15151 29563
rect 15151 29529 15160 29563
rect 15108 29520 15160 29529
rect 20904 29520 20956 29572
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 27528 29631 27580 29640
rect 27528 29597 27537 29631
rect 27537 29597 27571 29631
rect 27571 29597 27580 29631
rect 27528 29588 27580 29597
rect 27620 29631 27672 29640
rect 27620 29597 27629 29631
rect 27629 29597 27663 29631
rect 27663 29597 27672 29631
rect 27620 29588 27672 29597
rect 21640 29520 21692 29572
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 28908 29724 28960 29776
rect 29000 29656 29052 29708
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 29184 29588 29236 29640
rect 9312 29452 9364 29504
rect 9956 29452 10008 29504
rect 10416 29452 10468 29504
rect 12716 29452 12768 29504
rect 12808 29495 12860 29504
rect 12808 29461 12817 29495
rect 12817 29461 12851 29495
rect 12851 29461 12860 29495
rect 12808 29452 12860 29461
rect 19524 29495 19576 29504
rect 19524 29461 19533 29495
rect 19533 29461 19567 29495
rect 19567 29461 19576 29495
rect 19524 29452 19576 29461
rect 21456 29452 21508 29504
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 12900 29248 12952 29300
rect 14556 29291 14608 29300
rect 14556 29257 14565 29291
rect 14565 29257 14599 29291
rect 14599 29257 14608 29291
rect 14556 29248 14608 29257
rect 14924 29248 14976 29300
rect 9036 29155 9088 29164
rect 9036 29121 9045 29155
rect 9045 29121 9079 29155
rect 9079 29121 9088 29155
rect 9036 29112 9088 29121
rect 9312 29155 9364 29164
rect 9312 29121 9321 29155
rect 9321 29121 9355 29155
rect 9355 29121 9364 29155
rect 9312 29112 9364 29121
rect 9496 29155 9548 29164
rect 9496 29121 9505 29155
rect 9505 29121 9539 29155
rect 9539 29121 9548 29155
rect 9496 29112 9548 29121
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 15108 29180 15160 29232
rect 20168 29291 20220 29300
rect 20168 29257 20177 29291
rect 20177 29257 20211 29291
rect 20211 29257 20220 29291
rect 20168 29248 20220 29257
rect 21364 29248 21416 29300
rect 27160 29248 27212 29300
rect 27528 29248 27580 29300
rect 27620 29248 27672 29300
rect 28356 29248 28408 29300
rect 29184 29248 29236 29300
rect 12716 29112 12768 29164
rect 12808 29112 12860 29164
rect 13360 29112 13412 29164
rect 15568 29155 15620 29164
rect 15568 29121 15577 29155
rect 15577 29121 15611 29155
rect 15611 29121 15620 29155
rect 15568 29112 15620 29121
rect 16396 29112 16448 29164
rect 19340 29112 19392 29164
rect 19524 29155 19576 29164
rect 19524 29121 19533 29155
rect 19533 29121 19567 29155
rect 19567 29121 19576 29155
rect 19524 29112 19576 29121
rect 20536 29180 20588 29232
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 20628 29155 20680 29164
rect 20628 29121 20637 29155
rect 20637 29121 20671 29155
rect 20671 29121 20680 29155
rect 20628 29112 20680 29121
rect 20720 29155 20772 29164
rect 20720 29121 20729 29155
rect 20729 29121 20763 29155
rect 20763 29121 20772 29155
rect 20720 29112 20772 29121
rect 21640 29180 21692 29232
rect 12440 29087 12492 29096
rect 12440 29053 12449 29087
rect 12449 29053 12483 29087
rect 12483 29053 12492 29087
rect 12440 29044 12492 29053
rect 15016 29044 15068 29096
rect 22376 29112 22428 29164
rect 25228 29223 25280 29232
rect 25228 29189 25237 29223
rect 25237 29189 25271 29223
rect 25271 29189 25280 29223
rect 25228 29180 25280 29189
rect 22744 29155 22796 29164
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 23480 29112 23532 29164
rect 24492 29112 24544 29164
rect 26056 29112 26108 29164
rect 27160 29155 27212 29164
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 28080 29155 28132 29164
rect 28080 29121 28089 29155
rect 28089 29121 28123 29155
rect 28123 29121 28132 29155
rect 28080 29112 28132 29121
rect 26792 29044 26844 29096
rect 21272 29019 21324 29028
rect 21272 28985 21281 29019
rect 21281 28985 21315 29019
rect 21315 28985 21324 29019
rect 21272 28976 21324 28985
rect 8944 28908 8996 28960
rect 20720 28908 20772 28960
rect 23204 28976 23256 29028
rect 27436 28976 27488 29028
rect 29644 29044 29696 29096
rect 28908 28951 28960 28960
rect 28908 28917 28917 28951
rect 28917 28917 28951 28951
rect 28951 28917 28960 28951
rect 28908 28908 28960 28917
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 21180 28747 21232 28756
rect 21180 28713 21189 28747
rect 21189 28713 21223 28747
rect 21223 28713 21232 28747
rect 21180 28704 21232 28713
rect 28908 28704 28960 28756
rect 12440 28636 12492 28688
rect 12808 28636 12860 28688
rect 9496 28568 9548 28620
rect 11888 28568 11940 28620
rect 12532 28568 12584 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 15016 28568 15068 28620
rect 20812 28568 20864 28620
rect 9036 28432 9088 28484
rect 10692 28500 10744 28552
rect 12440 28500 12492 28552
rect 12624 28432 12676 28484
rect 13268 28543 13320 28552
rect 13268 28509 13277 28543
rect 13277 28509 13311 28543
rect 13311 28509 13320 28543
rect 13268 28500 13320 28509
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 15108 28500 15160 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 15752 28500 15804 28552
rect 16396 28500 16448 28552
rect 19616 28500 19668 28552
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 19984 28543 20036 28552
rect 19984 28509 19993 28543
rect 19993 28509 20027 28543
rect 20027 28509 20036 28543
rect 19984 28500 20036 28509
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 9312 28364 9364 28416
rect 12348 28364 12400 28416
rect 15936 28432 15988 28484
rect 18420 28432 18472 28484
rect 20720 28543 20772 28552
rect 20720 28509 20729 28543
rect 20729 28509 20763 28543
rect 20763 28509 20772 28543
rect 20720 28500 20772 28509
rect 20904 28543 20956 28552
rect 20904 28509 20913 28543
rect 20913 28509 20947 28543
rect 20947 28509 20956 28543
rect 20904 28500 20956 28509
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 23388 28500 23440 28552
rect 27344 28636 27396 28688
rect 26700 28568 26752 28620
rect 28356 28568 28408 28620
rect 27896 28500 27948 28552
rect 28724 28543 28776 28552
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 28724 28500 28776 28509
rect 23664 28432 23716 28484
rect 24676 28432 24728 28484
rect 22744 28364 22796 28416
rect 27252 28407 27304 28416
rect 27252 28373 27261 28407
rect 27261 28373 27295 28407
rect 27295 28373 27304 28407
rect 27252 28364 27304 28373
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 8944 28160 8996 28212
rect 13360 28160 13412 28212
rect 15384 28203 15436 28212
rect 15384 28169 15393 28203
rect 15393 28169 15427 28203
rect 15427 28169 15436 28203
rect 15384 28160 15436 28169
rect 8852 28092 8904 28144
rect 9128 28024 9180 28076
rect 12624 28092 12676 28144
rect 8760 27999 8812 28008
rect 8760 27965 8769 27999
rect 8769 27965 8803 27999
rect 8803 27965 8812 27999
rect 8760 27956 8812 27965
rect 8852 27999 8904 28008
rect 8852 27965 8861 27999
rect 8861 27965 8895 27999
rect 8895 27965 8904 27999
rect 8852 27956 8904 27965
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 10692 28024 10744 28076
rect 12348 28024 12400 28076
rect 12532 28067 12584 28076
rect 12532 28033 12541 28067
rect 12541 28033 12575 28067
rect 12575 28033 12584 28067
rect 12532 28024 12584 28033
rect 15016 28092 15068 28144
rect 15568 28092 15620 28144
rect 16028 28092 16080 28144
rect 13268 28024 13320 28076
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 14188 28067 14240 28076
rect 14188 28033 14197 28067
rect 14197 28033 14231 28067
rect 14231 28033 14240 28067
rect 14188 28024 14240 28033
rect 15752 28024 15804 28076
rect 19616 28160 19668 28212
rect 19892 28160 19944 28212
rect 19340 28092 19392 28144
rect 20904 28092 20956 28144
rect 22376 28160 22428 28212
rect 23204 28203 23256 28212
rect 23204 28169 23213 28203
rect 23213 28169 23247 28203
rect 23247 28169 23256 28203
rect 23204 28160 23256 28169
rect 26608 28092 26660 28144
rect 27344 28092 27396 28144
rect 31116 28092 31168 28144
rect 23664 28067 23716 28076
rect 8944 27956 8996 27965
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 14556 27956 14608 28008
rect 19984 27956 20036 28008
rect 9128 27820 9180 27872
rect 9312 27820 9364 27872
rect 9588 27820 9640 27872
rect 9772 27863 9824 27872
rect 9772 27829 9781 27863
rect 9781 27829 9815 27863
rect 9815 27829 9824 27863
rect 9772 27820 9824 27829
rect 23664 28033 23673 28067
rect 23673 28033 23707 28067
rect 23707 28033 23716 28067
rect 23664 28024 23716 28033
rect 25044 28067 25096 28076
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 25412 28024 25464 28076
rect 27068 28024 27120 28076
rect 27712 28024 27764 28076
rect 30012 28067 30064 28076
rect 30012 28033 30021 28067
rect 30021 28033 30055 28067
rect 30055 28033 30064 28067
rect 30012 28024 30064 28033
rect 32680 28024 32732 28076
rect 25136 27956 25188 28008
rect 26056 27999 26108 28008
rect 26056 27965 26065 27999
rect 26065 27965 26099 27999
rect 26099 27965 26108 27999
rect 26056 27956 26108 27965
rect 26516 27956 26568 28008
rect 23388 27931 23440 27940
rect 23388 27897 23397 27931
rect 23397 27897 23431 27931
rect 23431 27897 23440 27931
rect 23388 27888 23440 27897
rect 25872 27888 25924 27940
rect 24676 27820 24728 27872
rect 29828 27863 29880 27872
rect 29828 27829 29837 27863
rect 29837 27829 29871 27863
rect 29871 27829 29880 27863
rect 29828 27820 29880 27829
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 16028 27548 16080 27600
rect 24860 27548 24912 27600
rect 9036 27480 9088 27532
rect 12532 27480 12584 27532
rect 9128 27412 9180 27464
rect 9588 27412 9640 27464
rect 14004 27480 14056 27532
rect 14188 27412 14240 27464
rect 17224 27480 17276 27532
rect 8208 27344 8260 27396
rect 12348 27344 12400 27396
rect 12716 27344 12768 27396
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 20904 27480 20956 27532
rect 20996 27480 21048 27532
rect 21916 27480 21968 27532
rect 25044 27480 25096 27532
rect 25320 27480 25372 27532
rect 18236 27455 18288 27464
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 22008 27455 22060 27464
rect 22008 27421 22017 27455
rect 22017 27421 22051 27455
rect 22051 27421 22060 27455
rect 22008 27412 22060 27421
rect 26056 27548 26108 27600
rect 20260 27344 20312 27396
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 26516 27480 26568 27532
rect 25596 27344 25648 27396
rect 26148 27412 26200 27464
rect 27896 27591 27948 27600
rect 27896 27557 27905 27591
rect 27905 27557 27939 27591
rect 27939 27557 27948 27591
rect 27896 27548 27948 27557
rect 19800 27276 19852 27328
rect 21916 27276 21968 27328
rect 22376 27276 22428 27328
rect 25872 27276 25924 27328
rect 27528 27412 27580 27464
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 27068 27276 27120 27328
rect 29920 27412 29972 27464
rect 32220 27344 32272 27396
rect 28724 27276 28776 27328
rect 32588 27276 32640 27328
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 12072 27072 12124 27124
rect 12900 27072 12952 27124
rect 18236 27072 18288 27124
rect 19800 27072 19852 27124
rect 9128 27004 9180 27056
rect 10600 27004 10652 27056
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 9772 26936 9824 26988
rect 12716 27004 12768 27056
rect 13452 27004 13504 27056
rect 12072 26979 12124 26988
rect 12072 26945 12081 26979
rect 12081 26945 12115 26979
rect 12115 26945 12124 26979
rect 12072 26936 12124 26945
rect 12440 26936 12492 26988
rect 14188 27004 14240 27056
rect 31116 27115 31168 27124
rect 31116 27081 31125 27115
rect 31125 27081 31159 27115
rect 31159 27081 31168 27115
rect 31116 27072 31168 27081
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 16396 26936 16448 26988
rect 18328 26936 18380 26988
rect 20904 26936 20956 26988
rect 9128 26911 9180 26920
rect 9128 26877 9137 26911
rect 9137 26877 9171 26911
rect 9171 26877 9180 26911
rect 9128 26868 9180 26877
rect 21364 26936 21416 26988
rect 22008 26936 22060 26988
rect 22928 27004 22980 27056
rect 25412 27004 25464 27056
rect 24768 26936 24820 26988
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 26148 27004 26200 27056
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 29828 26936 29880 26988
rect 26148 26868 26200 26920
rect 28356 26868 28408 26920
rect 29920 26868 29972 26920
rect 8760 26732 8812 26784
rect 21640 26800 21692 26852
rect 27160 26800 27212 26852
rect 27528 26800 27580 26852
rect 9220 26732 9272 26784
rect 11152 26732 11204 26784
rect 12624 26732 12676 26784
rect 18420 26732 18472 26784
rect 20904 26732 20956 26784
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 12440 26528 12492 26580
rect 12900 26528 12952 26580
rect 13360 26528 13412 26580
rect 15660 26528 15712 26580
rect 17132 26528 17184 26580
rect 25136 26528 25188 26580
rect 27068 26571 27120 26580
rect 27068 26537 27077 26571
rect 27077 26537 27111 26571
rect 27111 26537 27120 26571
rect 27068 26528 27120 26537
rect 32220 26571 32272 26580
rect 32220 26537 32229 26571
rect 32229 26537 32263 26571
rect 32263 26537 32272 26571
rect 32220 26528 32272 26537
rect 9312 26460 9364 26512
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 26700 26460 26752 26512
rect 14740 26392 14792 26444
rect 18236 26392 18288 26444
rect 19340 26392 19392 26444
rect 12624 26367 12676 26376
rect 12624 26333 12633 26367
rect 12633 26333 12667 26367
rect 12667 26333 12676 26367
rect 12624 26324 12676 26333
rect 24584 26392 24636 26444
rect 28632 26460 28684 26512
rect 9036 26256 9088 26308
rect 12532 26256 12584 26308
rect 13452 26299 13504 26308
rect 13452 26265 13463 26299
rect 13463 26265 13504 26299
rect 13452 26256 13504 26265
rect 13544 26256 13596 26308
rect 16856 26256 16908 26308
rect 18236 26256 18288 26308
rect 20076 26324 20128 26376
rect 21364 26324 21416 26376
rect 25320 26324 25372 26376
rect 25504 26367 25556 26376
rect 25504 26333 25513 26367
rect 25513 26333 25547 26367
rect 25547 26333 25556 26367
rect 25504 26324 25556 26333
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 20260 26256 20312 26308
rect 22560 26299 22612 26308
rect 22560 26265 22569 26299
rect 22569 26265 22603 26299
rect 22603 26265 22612 26299
rect 22560 26256 22612 26265
rect 22744 26256 22796 26308
rect 9312 26188 9364 26240
rect 21180 26188 21232 26240
rect 26516 26367 26568 26376
rect 26516 26333 26525 26367
rect 26525 26333 26559 26367
rect 26559 26333 26568 26367
rect 26516 26324 26568 26333
rect 26792 26367 26844 26376
rect 26792 26333 26801 26367
rect 26801 26333 26835 26367
rect 26835 26333 26844 26367
rect 26792 26324 26844 26333
rect 26884 26367 26936 26376
rect 26884 26333 26893 26367
rect 26893 26333 26927 26367
rect 26927 26333 26936 26367
rect 26884 26324 26936 26333
rect 32404 26367 32456 26376
rect 32404 26333 32413 26367
rect 32413 26333 32447 26367
rect 32447 26333 32456 26367
rect 32404 26324 32456 26333
rect 32588 26367 32640 26376
rect 32588 26333 32597 26367
rect 32597 26333 32631 26367
rect 32631 26333 32640 26367
rect 32588 26324 32640 26333
rect 32680 26367 32732 26376
rect 32680 26333 32689 26367
rect 32689 26333 32723 26367
rect 32723 26333 32732 26367
rect 32680 26324 32732 26333
rect 27620 26256 27672 26308
rect 29092 26256 29144 26308
rect 26608 26188 26660 26240
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 9220 25984 9272 26036
rect 9312 25848 9364 25900
rect 12348 26027 12400 26036
rect 12348 25993 12357 26027
rect 12357 25993 12391 26027
rect 12391 25993 12400 26027
rect 12348 25984 12400 25993
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 12440 25984 12492 25993
rect 12072 25959 12124 25968
rect 12072 25925 12081 25959
rect 12081 25925 12115 25959
rect 12115 25925 12124 25959
rect 12072 25916 12124 25925
rect 12532 25916 12584 25968
rect 16856 26027 16908 26036
rect 16856 25993 16865 26027
rect 16865 25993 16899 26027
rect 16899 25993 16908 26027
rect 16856 25984 16908 25993
rect 17132 25984 17184 26036
rect 25688 25984 25740 26036
rect 27252 25984 27304 26036
rect 29920 26027 29972 26036
rect 29920 25993 29929 26027
rect 29929 25993 29963 26027
rect 29963 25993 29972 26027
rect 29920 25984 29972 25993
rect 13360 25959 13412 25968
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 21916 25916 21968 25968
rect 25504 25916 25556 25968
rect 26792 25916 26844 25968
rect 9220 25780 9272 25832
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 12348 25848 12400 25900
rect 13452 25891 13504 25900
rect 13452 25857 13466 25891
rect 13466 25857 13500 25891
rect 13500 25857 13504 25891
rect 13452 25848 13504 25857
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17224 25848 17276 25900
rect 17684 25848 17736 25900
rect 19616 25891 19668 25900
rect 19616 25857 19625 25891
rect 19625 25857 19659 25891
rect 19659 25857 19668 25891
rect 19616 25848 19668 25857
rect 14648 25780 14700 25832
rect 14464 25712 14516 25764
rect 21180 25848 21232 25900
rect 22376 25848 22428 25900
rect 23572 25848 23624 25900
rect 23480 25823 23532 25832
rect 23480 25789 23489 25823
rect 23489 25789 23523 25823
rect 23523 25789 23532 25823
rect 23480 25780 23532 25789
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 24860 25848 24912 25900
rect 26516 25891 26568 25900
rect 26516 25857 26525 25891
rect 26525 25857 26559 25891
rect 26559 25857 26568 25891
rect 26516 25848 26568 25857
rect 26884 25848 26936 25900
rect 28632 25891 28684 25900
rect 28632 25857 28641 25891
rect 28641 25857 28675 25891
rect 28675 25857 28684 25891
rect 28632 25848 28684 25857
rect 31944 25848 31996 25900
rect 32680 25891 32732 25900
rect 32680 25857 32689 25891
rect 32689 25857 32723 25891
rect 32723 25857 32732 25891
rect 32680 25848 32732 25857
rect 32772 25891 32824 25900
rect 32772 25857 32781 25891
rect 32781 25857 32815 25891
rect 32815 25857 32824 25891
rect 32772 25848 32824 25857
rect 25228 25780 25280 25832
rect 25136 25712 25188 25764
rect 27068 25780 27120 25832
rect 27620 25823 27672 25832
rect 27620 25789 27629 25823
rect 27629 25789 27663 25823
rect 27663 25789 27672 25823
rect 27620 25780 27672 25789
rect 28264 25780 28316 25832
rect 12716 25644 12768 25696
rect 13084 25687 13136 25696
rect 13084 25653 13093 25687
rect 13093 25653 13127 25687
rect 13127 25653 13136 25687
rect 13084 25644 13136 25653
rect 18328 25687 18380 25696
rect 18328 25653 18337 25687
rect 18337 25653 18371 25687
rect 18371 25653 18380 25687
rect 18328 25644 18380 25653
rect 25872 25644 25924 25696
rect 26056 25644 26108 25696
rect 32312 25687 32364 25696
rect 32312 25653 32321 25687
rect 32321 25653 32355 25687
rect 32355 25653 32364 25687
rect 32312 25644 32364 25653
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 15660 25440 15712 25492
rect 19800 25483 19852 25492
rect 19800 25449 19809 25483
rect 19809 25449 19843 25483
rect 19843 25449 19852 25483
rect 19800 25440 19852 25449
rect 25596 25440 25648 25492
rect 26700 25440 26752 25492
rect 28264 25483 28316 25492
rect 28264 25449 28273 25483
rect 28273 25449 28307 25483
rect 28307 25449 28316 25483
rect 28264 25440 28316 25449
rect 3332 25236 3384 25288
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 4804 25236 4856 25288
rect 6828 25236 6880 25288
rect 7472 25236 7524 25288
rect 10692 25236 10744 25288
rect 13084 25304 13136 25356
rect 16304 25415 16356 25424
rect 16304 25381 16313 25415
rect 16313 25381 16347 25415
rect 16347 25381 16356 25415
rect 16304 25372 16356 25381
rect 26608 25415 26660 25424
rect 26608 25381 26617 25415
rect 26617 25381 26651 25415
rect 26651 25381 26660 25415
rect 26608 25372 26660 25381
rect 3976 25211 4028 25220
rect 3976 25177 3985 25211
rect 3985 25177 4019 25211
rect 4019 25177 4028 25211
rect 3976 25168 4028 25177
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 15384 25236 15436 25288
rect 2872 25100 2924 25152
rect 5540 25100 5592 25152
rect 13452 25100 13504 25152
rect 15200 25143 15252 25152
rect 15200 25109 15209 25143
rect 15209 25109 15243 25143
rect 15243 25109 15252 25143
rect 15200 25100 15252 25109
rect 15936 25236 15988 25288
rect 21180 25347 21232 25356
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 20904 25279 20956 25288
rect 20904 25245 20922 25279
rect 20922 25245 20956 25279
rect 20904 25236 20956 25245
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 27344 25279 27396 25288
rect 27344 25245 27352 25279
rect 27352 25245 27386 25279
rect 27386 25245 27396 25279
rect 27344 25236 27396 25245
rect 21088 25168 21140 25220
rect 24860 25211 24912 25220
rect 24860 25177 24869 25211
rect 24869 25177 24903 25211
rect 24903 25177 24912 25211
rect 24860 25168 24912 25177
rect 25228 25168 25280 25220
rect 26516 25168 26568 25220
rect 28908 25236 28960 25288
rect 30104 25279 30156 25288
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 15752 25100 15804 25152
rect 18420 25100 18472 25152
rect 22560 25100 22612 25152
rect 27068 25143 27120 25152
rect 27068 25109 27077 25143
rect 27077 25109 27111 25143
rect 27111 25109 27120 25143
rect 27068 25100 27120 25109
rect 30380 25211 30432 25220
rect 30380 25177 30414 25211
rect 30414 25177 30432 25211
rect 30380 25168 30432 25177
rect 30932 25100 30984 25152
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 17040 24896 17092 24948
rect 5080 24828 5132 24880
rect 2780 24692 2832 24744
rect 3976 24760 4028 24812
rect 6828 24760 6880 24812
rect 7472 24760 7524 24812
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 4712 24735 4764 24744
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 8392 24692 8444 24744
rect 15200 24760 15252 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 15476 24692 15528 24744
rect 6736 24624 6788 24676
rect 16304 24760 16356 24812
rect 17684 24760 17736 24812
rect 17316 24692 17368 24744
rect 18236 24760 18288 24812
rect 20812 24760 20864 24812
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 20904 24692 20956 24744
rect 21364 24760 21416 24812
rect 25136 24939 25188 24948
rect 25136 24905 25145 24939
rect 25145 24905 25179 24939
rect 25179 24905 25188 24939
rect 25136 24896 25188 24905
rect 23572 24760 23624 24812
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 25320 24803 25372 24812
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 25320 24760 25372 24769
rect 27068 24828 27120 24880
rect 28724 24760 28776 24812
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 32312 24760 32364 24812
rect 21272 24624 21324 24676
rect 4068 24556 4120 24608
rect 4344 24556 4396 24608
rect 14924 24556 14976 24608
rect 21548 24556 21600 24608
rect 27160 24692 27212 24744
rect 30104 24735 30156 24744
rect 30104 24701 30113 24735
rect 30113 24701 30147 24735
rect 30147 24701 30156 24735
rect 30104 24692 30156 24701
rect 26608 24624 26660 24676
rect 23480 24556 23532 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 28908 24556 28960 24608
rect 32680 24624 32732 24676
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 2780 24395 2832 24404
rect 2780 24361 2789 24395
rect 2789 24361 2823 24395
rect 2823 24361 2832 24395
rect 2780 24352 2832 24361
rect 6828 24395 6880 24404
rect 6828 24361 6837 24395
rect 6837 24361 6871 24395
rect 6871 24361 6880 24395
rect 6828 24352 6880 24361
rect 2780 24216 2832 24268
rect 2320 24123 2372 24132
rect 2320 24089 2329 24123
rect 2329 24089 2363 24123
rect 2363 24089 2372 24123
rect 2320 24080 2372 24089
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 5080 24216 5132 24268
rect 7288 24216 7340 24268
rect 13452 24216 13504 24268
rect 3424 24123 3476 24132
rect 3424 24089 3433 24123
rect 3433 24089 3467 24123
rect 3467 24089 3476 24123
rect 3424 24080 3476 24089
rect 4252 24012 4304 24064
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 7012 24148 7064 24200
rect 8208 24148 8260 24200
rect 9312 24148 9364 24200
rect 11980 24148 12032 24200
rect 12440 24148 12492 24200
rect 13268 24148 13320 24200
rect 7840 24080 7892 24132
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 15016 24216 15068 24268
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 16396 24148 16448 24200
rect 20904 24352 20956 24404
rect 21824 24352 21876 24404
rect 24584 24352 24636 24404
rect 30380 24352 30432 24404
rect 30012 24284 30064 24336
rect 21088 24216 21140 24268
rect 23848 24216 23900 24268
rect 32404 24216 32456 24268
rect 17960 24148 18012 24200
rect 20628 24191 20680 24200
rect 20628 24157 20637 24191
rect 20637 24157 20671 24191
rect 20671 24157 20680 24191
rect 20628 24148 20680 24157
rect 5816 24012 5868 24064
rect 10508 24012 10560 24064
rect 12624 24012 12676 24064
rect 12900 24012 12952 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 18696 24080 18748 24132
rect 19708 24080 19760 24132
rect 21272 24148 21324 24200
rect 23572 24148 23624 24200
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 25872 24148 25924 24200
rect 30840 24148 30892 24200
rect 30932 24191 30984 24200
rect 30932 24157 30941 24191
rect 30941 24157 30975 24191
rect 30975 24157 30984 24191
rect 30932 24148 30984 24157
rect 15660 24012 15712 24064
rect 17132 24055 17184 24064
rect 17132 24021 17141 24055
rect 17141 24021 17175 24055
rect 17175 24021 17184 24055
rect 17132 24012 17184 24021
rect 17592 24012 17644 24064
rect 20812 24012 20864 24064
rect 23664 24055 23716 24064
rect 23664 24021 23673 24055
rect 23673 24021 23707 24055
rect 23707 24021 23716 24055
rect 23664 24012 23716 24021
rect 25320 24055 25372 24064
rect 25320 24021 25329 24055
rect 25329 24021 25363 24055
rect 25363 24021 25372 24055
rect 25320 24012 25372 24021
rect 25504 24080 25556 24132
rect 32772 24148 32824 24200
rect 26792 24012 26844 24064
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 2320 23808 2372 23860
rect 4712 23740 4764 23792
rect 4804 23740 4856 23792
rect 4528 23672 4580 23724
rect 5816 23740 5868 23792
rect 3332 23536 3384 23588
rect 4344 23536 4396 23588
rect 4896 23468 4948 23520
rect 7196 23672 7248 23724
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 15292 23808 15344 23860
rect 18236 23808 18288 23860
rect 18420 23808 18472 23860
rect 21364 23808 21416 23860
rect 8392 23740 8444 23792
rect 15016 23740 15068 23792
rect 20904 23740 20956 23792
rect 21916 23740 21968 23792
rect 25228 23808 25280 23860
rect 30104 23851 30156 23860
rect 30104 23817 30113 23851
rect 30113 23817 30147 23851
rect 30147 23817 30156 23851
rect 30104 23808 30156 23817
rect 28632 23783 28684 23792
rect 28632 23749 28641 23783
rect 28641 23749 28675 23783
rect 28675 23749 28684 23783
rect 28632 23740 28684 23749
rect 10048 23715 10100 23724
rect 10048 23681 10057 23715
rect 10057 23681 10091 23715
rect 10091 23681 10100 23715
rect 10048 23672 10100 23681
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 15476 23672 15528 23724
rect 17132 23672 17184 23724
rect 19524 23672 19576 23724
rect 6736 23604 6788 23656
rect 7104 23647 7156 23656
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 8300 23604 8352 23656
rect 9588 23604 9640 23656
rect 10508 23604 10560 23656
rect 7840 23536 7892 23588
rect 13176 23647 13228 23656
rect 13176 23613 13185 23647
rect 13185 23613 13219 23647
rect 13219 23613 13228 23647
rect 13176 23604 13228 23613
rect 14648 23604 14700 23656
rect 15200 23647 15252 23656
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 15384 23604 15436 23656
rect 16488 23604 16540 23656
rect 14188 23536 14240 23588
rect 19708 23536 19760 23588
rect 20720 23715 20772 23724
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 21548 23672 21600 23724
rect 23480 23672 23532 23724
rect 23664 23672 23716 23724
rect 24860 23672 24912 23724
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 28816 23536 28868 23588
rect 7472 23468 7524 23520
rect 15476 23511 15528 23520
rect 15476 23477 15485 23511
rect 15485 23477 15519 23511
rect 15519 23477 15528 23511
rect 15476 23468 15528 23477
rect 24952 23468 25004 23520
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 2872 23264 2924 23316
rect 3424 23264 3476 23316
rect 4436 23264 4488 23316
rect 4804 23264 4856 23316
rect 7104 23264 7156 23316
rect 10324 23307 10376 23316
rect 4896 23196 4948 23248
rect 10324 23273 10333 23307
rect 10333 23273 10367 23307
rect 10367 23273 10376 23307
rect 10324 23264 10376 23273
rect 11980 23264 12032 23316
rect 18696 23307 18748 23316
rect 18696 23273 18705 23307
rect 18705 23273 18739 23307
rect 18739 23273 18748 23307
rect 18696 23264 18748 23273
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 31852 23264 31904 23316
rect 33140 23264 33192 23316
rect 3976 23128 4028 23180
rect 8668 23196 8720 23248
rect 8300 23171 8352 23180
rect 8300 23137 8309 23171
rect 8309 23137 8343 23171
rect 8343 23137 8352 23171
rect 8300 23128 8352 23137
rect 8484 23128 8536 23180
rect 19616 23196 19668 23248
rect 19984 23196 20036 23248
rect 28724 23196 28776 23248
rect 3148 23103 3200 23112
rect 3148 23069 3157 23103
rect 3157 23069 3191 23103
rect 3191 23069 3200 23103
rect 3148 23060 3200 23069
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 7196 23103 7248 23112
rect 7196 23069 7205 23103
rect 7205 23069 7239 23103
rect 7239 23069 7248 23103
rect 7196 23060 7248 23069
rect 7564 23103 7616 23112
rect 7564 23069 7573 23103
rect 7573 23069 7607 23103
rect 7607 23069 7616 23103
rect 7564 23060 7616 23069
rect 14924 23128 14976 23180
rect 15200 23171 15252 23180
rect 15200 23137 15209 23171
rect 15209 23137 15243 23171
rect 15243 23137 15252 23171
rect 15200 23128 15252 23137
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 15476 23128 15528 23180
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 25320 23171 25372 23180
rect 25320 23137 25329 23171
rect 25329 23137 25363 23171
rect 25363 23137 25372 23171
rect 25320 23128 25372 23137
rect 31392 23128 31444 23180
rect 32680 23171 32732 23180
rect 32680 23137 32689 23171
rect 32689 23137 32723 23171
rect 32723 23137 32732 23171
rect 32680 23128 32732 23137
rect 33140 23171 33192 23180
rect 33140 23137 33149 23171
rect 33149 23137 33183 23171
rect 33183 23137 33192 23171
rect 33140 23128 33192 23137
rect 4344 23035 4396 23044
rect 4344 23001 4353 23035
rect 4353 23001 4387 23035
rect 4387 23001 4396 23035
rect 4344 22992 4396 23001
rect 3976 22967 4028 22976
rect 3976 22933 3985 22967
rect 3985 22933 4019 22967
rect 4019 22933 4028 22967
rect 3976 22924 4028 22933
rect 4712 22924 4764 22976
rect 8668 22992 8720 23044
rect 9312 23060 9364 23112
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 9772 22992 9824 23044
rect 11520 22992 11572 23044
rect 14648 23060 14700 23112
rect 15016 23060 15068 23112
rect 17592 23103 17644 23112
rect 17592 23069 17626 23103
rect 17626 23069 17644 23103
rect 17592 23060 17644 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20812 23060 20864 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 27528 23103 27580 23112
rect 27528 23069 27537 23103
rect 27537 23069 27571 23103
rect 27571 23069 27580 23103
rect 27528 23060 27580 23069
rect 28080 23103 28132 23112
rect 28080 23069 28089 23103
rect 28089 23069 28123 23103
rect 28123 23069 28132 23103
rect 28080 23060 28132 23069
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 31760 23103 31812 23112
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32036 23103 32088 23112
rect 32036 23069 32045 23103
rect 32045 23069 32079 23103
rect 32079 23069 32088 23103
rect 32036 23060 32088 23069
rect 32404 23060 32456 23112
rect 33324 23060 33376 23112
rect 7840 22924 7892 22976
rect 8208 22924 8260 22976
rect 10232 22924 10284 22976
rect 10416 22924 10468 22976
rect 10876 22924 10928 22976
rect 25320 22992 25372 23044
rect 27620 22992 27672 23044
rect 14648 22924 14700 22976
rect 25136 22967 25188 22976
rect 25136 22933 25145 22967
rect 25145 22933 25179 22967
rect 25179 22933 25188 22967
rect 25136 22924 25188 22933
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 29736 22924 29788 22976
rect 33508 22924 33560 22976
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 7564 22720 7616 22772
rect 7840 22720 7892 22772
rect 7104 22652 7156 22704
rect 10048 22720 10100 22772
rect 8392 22652 8444 22704
rect 9312 22652 9364 22704
rect 4252 22584 4304 22636
rect 7012 22584 7064 22636
rect 7472 22584 7524 22636
rect 9772 22652 9824 22704
rect 4528 22491 4580 22500
rect 4528 22457 4537 22491
rect 4537 22457 4571 22491
rect 4571 22457 4580 22491
rect 4528 22448 4580 22457
rect 8484 22448 8536 22500
rect 10416 22584 10468 22636
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 12440 22584 12492 22636
rect 12624 22584 12676 22636
rect 11796 22516 11848 22568
rect 11980 22448 12032 22500
rect 12900 22448 12952 22500
rect 13452 22584 13504 22636
rect 31852 22720 31904 22772
rect 32036 22720 32088 22772
rect 15016 22652 15068 22704
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 15292 22627 15344 22636
rect 15292 22593 15301 22627
rect 15301 22593 15335 22627
rect 15335 22593 15344 22627
rect 15292 22584 15344 22593
rect 14188 22516 14240 22568
rect 15660 22584 15712 22636
rect 16304 22584 16356 22636
rect 17132 22584 17184 22636
rect 18144 22652 18196 22704
rect 18696 22652 18748 22704
rect 20168 22652 20220 22704
rect 20628 22652 20680 22704
rect 19984 22627 20036 22636
rect 15936 22516 15988 22568
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 18236 22559 18288 22568
rect 18236 22525 18245 22559
rect 18245 22525 18279 22559
rect 18279 22525 18288 22559
rect 18236 22516 18288 22525
rect 18052 22448 18104 22500
rect 20536 22584 20588 22636
rect 25228 22695 25280 22704
rect 25228 22661 25237 22695
rect 25237 22661 25271 22695
rect 25271 22661 25280 22695
rect 25228 22652 25280 22661
rect 27620 22652 27672 22704
rect 27160 22584 27212 22636
rect 28172 22627 28224 22636
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 28172 22584 28224 22593
rect 28264 22584 28316 22636
rect 23848 22516 23900 22568
rect 26148 22516 26200 22568
rect 29736 22559 29788 22568
rect 29736 22525 29745 22559
rect 29745 22525 29779 22559
rect 29779 22525 29788 22559
rect 29736 22516 29788 22525
rect 25780 22448 25832 22500
rect 27988 22448 28040 22500
rect 31116 22559 31168 22568
rect 31116 22525 31125 22559
rect 31125 22525 31159 22559
rect 31159 22525 31168 22559
rect 31116 22516 31168 22525
rect 31208 22559 31260 22568
rect 31208 22525 31217 22559
rect 31217 22525 31251 22559
rect 31251 22525 31260 22559
rect 31208 22516 31260 22525
rect 33140 22652 33192 22704
rect 33508 22695 33560 22704
rect 33508 22661 33517 22695
rect 33517 22661 33551 22695
rect 33551 22661 33560 22695
rect 33508 22652 33560 22661
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33692 22627 33744 22636
rect 33692 22593 33701 22627
rect 33701 22593 33735 22627
rect 33735 22593 33744 22627
rect 33692 22584 33744 22593
rect 32404 22516 32456 22568
rect 33324 22516 33376 22568
rect 4344 22380 4396 22432
rect 9220 22380 9272 22432
rect 10232 22380 10284 22432
rect 10416 22380 10468 22432
rect 12992 22380 13044 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19800 22423 19852 22432
rect 19800 22389 19809 22423
rect 19809 22389 19843 22423
rect 19843 22389 19852 22423
rect 19800 22380 19852 22389
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 26976 22380 27028 22432
rect 30840 22423 30892 22432
rect 30840 22389 30849 22423
rect 30849 22389 30883 22423
rect 30883 22389 30892 22423
rect 30840 22380 30892 22389
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 4988 22176 5040 22228
rect 11520 22176 11572 22228
rect 11704 22219 11756 22228
rect 11704 22185 11725 22219
rect 11725 22185 11756 22219
rect 11704 22176 11756 22185
rect 15292 22176 15344 22228
rect 12440 22108 12492 22160
rect 17960 22108 18012 22160
rect 19248 22108 19300 22160
rect 21640 22108 21692 22160
rect 22652 22176 22704 22228
rect 33692 22176 33744 22228
rect 3148 22040 3200 22092
rect 11060 22040 11112 22092
rect 11612 22040 11664 22092
rect 12072 22040 12124 22092
rect 7104 21972 7156 22024
rect 7472 21972 7524 22024
rect 9312 21972 9364 22024
rect 11704 21904 11756 21956
rect 12900 22015 12952 22024
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 25228 22040 25280 22092
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 29920 22040 29972 22092
rect 30380 22108 30432 22160
rect 30840 22108 30892 22160
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 19432 21972 19484 22024
rect 20904 21972 20956 22024
rect 22928 21972 22980 22024
rect 24584 21972 24636 22024
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 10692 21836 10744 21888
rect 16488 21836 16540 21888
rect 19616 21904 19668 21956
rect 20260 21904 20312 21956
rect 21088 21904 21140 21956
rect 25964 21972 26016 22024
rect 25136 21904 25188 21956
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 25044 21836 25096 21888
rect 27068 21972 27120 22024
rect 27344 21972 27396 22024
rect 27528 21904 27580 21956
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 31024 22015 31076 22024
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31024 21972 31076 21981
rect 31208 21972 31260 22024
rect 33140 22083 33192 22092
rect 33140 22049 33149 22083
rect 33149 22049 33183 22083
rect 33183 22049 33192 22083
rect 33140 22040 33192 22049
rect 31576 22015 31628 22024
rect 31576 21981 31585 22015
rect 31585 21981 31619 22015
rect 31619 21981 31628 22015
rect 31576 21972 31628 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 30288 21904 30340 21956
rect 26976 21836 27028 21888
rect 27068 21836 27120 21888
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 31024 21836 31076 21888
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 9864 21632 9916 21684
rect 11704 21607 11756 21616
rect 11704 21573 11713 21607
rect 11713 21573 11747 21607
rect 11747 21573 11756 21607
rect 11704 21564 11756 21573
rect 3976 21496 4028 21548
rect 4528 21496 4580 21548
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 27068 21632 27120 21684
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 29092 21632 29144 21684
rect 30288 21675 30340 21684
rect 30288 21641 30297 21675
rect 30297 21641 30331 21675
rect 30331 21641 30340 21675
rect 30288 21632 30340 21641
rect 31760 21632 31812 21684
rect 15844 21496 15896 21548
rect 17684 21496 17736 21548
rect 19524 21539 19576 21548
rect 19524 21505 19533 21539
rect 19533 21505 19567 21539
rect 19567 21505 19576 21539
rect 19524 21496 19576 21505
rect 19800 21539 19852 21548
rect 19800 21505 19809 21539
rect 19809 21505 19843 21539
rect 19843 21505 19852 21539
rect 19800 21496 19852 21505
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 18236 21428 18288 21480
rect 4068 21360 4120 21412
rect 19156 21360 19208 21412
rect 22284 21539 22336 21548
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 23572 21428 23624 21480
rect 23940 21428 23992 21480
rect 27988 21496 28040 21548
rect 28448 21564 28500 21616
rect 27620 21428 27672 21480
rect 29736 21496 29788 21548
rect 30380 21564 30432 21616
rect 31024 21564 31076 21616
rect 31116 21496 31168 21548
rect 32588 21496 32640 21548
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3056 21292 3108 21301
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 16672 21292 16724 21344
rect 19432 21335 19484 21344
rect 19432 21301 19441 21335
rect 19441 21301 19475 21335
rect 19475 21301 19484 21335
rect 19432 21292 19484 21301
rect 23848 21292 23900 21344
rect 27896 21292 27948 21344
rect 28448 21292 28500 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 12900 21088 12952 21140
rect 17316 21088 17368 21140
rect 21272 21131 21324 21140
rect 21272 21097 21281 21131
rect 21281 21097 21315 21131
rect 21315 21097 21324 21131
rect 21272 21088 21324 21097
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 23848 21088 23900 21140
rect 31944 21088 31996 21140
rect 32404 21131 32456 21140
rect 32404 21097 32413 21131
rect 32413 21097 32447 21131
rect 32447 21097 32456 21131
rect 32404 21088 32456 21097
rect 25872 21020 25924 21072
rect 31116 21020 31168 21072
rect 4528 20952 4580 21004
rect 7472 20952 7524 21004
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 3516 20884 3568 20936
rect 7288 20884 7340 20936
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 11888 20952 11940 21004
rect 19432 20952 19484 21004
rect 19984 20952 20036 21004
rect 21180 20952 21232 21004
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 13452 20884 13504 20936
rect 14464 20884 14516 20936
rect 18328 20884 18380 20936
rect 19156 20884 19208 20936
rect 28448 20952 28500 21004
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 3148 20748 3200 20800
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 21364 20816 21416 20868
rect 21640 20816 21692 20868
rect 23848 20884 23900 20936
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 24032 20927 24084 20936
rect 24032 20893 24041 20927
rect 24041 20893 24075 20927
rect 24075 20893 24084 20927
rect 24032 20884 24084 20893
rect 23388 20816 23440 20868
rect 24952 20884 25004 20936
rect 25136 20884 25188 20936
rect 25504 20884 25556 20936
rect 21088 20748 21140 20800
rect 30932 20816 30984 20868
rect 32128 20884 32180 20936
rect 32312 20884 32364 20936
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 32772 20816 32824 20868
rect 33048 20816 33100 20868
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 7840 20587 7892 20596
rect 7840 20553 7849 20587
rect 7849 20553 7883 20587
rect 7883 20553 7892 20587
rect 7840 20544 7892 20553
rect 3056 20476 3108 20528
rect 3424 20476 3476 20528
rect 3608 20519 3660 20528
rect 3608 20485 3617 20519
rect 3617 20485 3651 20519
rect 3651 20485 3660 20519
rect 3608 20476 3660 20485
rect 7748 20476 7800 20528
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3976 20408 4028 20460
rect 5080 20408 5132 20460
rect 7288 20408 7340 20460
rect 8024 20408 8076 20460
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 8392 20408 8444 20460
rect 10232 20408 10284 20460
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 14188 20544 14240 20596
rect 19892 20544 19944 20596
rect 20904 20544 20956 20596
rect 24860 20544 24912 20596
rect 31576 20587 31628 20596
rect 31576 20553 31585 20587
rect 31585 20553 31619 20587
rect 31619 20553 31628 20587
rect 31576 20544 31628 20553
rect 32588 20587 32640 20596
rect 32588 20553 32597 20587
rect 32597 20553 32631 20587
rect 32631 20553 32640 20587
rect 32588 20544 32640 20553
rect 14372 20476 14424 20528
rect 2412 20272 2464 20324
rect 9036 20340 9088 20392
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 13360 20340 13412 20392
rect 15568 20476 15620 20528
rect 12808 20272 12860 20324
rect 14188 20340 14240 20392
rect 14924 20340 14976 20392
rect 14096 20272 14148 20324
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 21364 20476 21416 20528
rect 22376 20476 22428 20528
rect 29092 20476 29144 20528
rect 32128 20476 32180 20528
rect 20076 20408 20128 20460
rect 20628 20408 20680 20460
rect 21272 20408 21324 20460
rect 27896 20451 27948 20460
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 18788 20272 18840 20324
rect 20996 20340 21048 20392
rect 32496 20408 32548 20460
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33048 20451 33100 20460
rect 33048 20417 33057 20451
rect 33057 20417 33091 20451
rect 33091 20417 33100 20451
rect 33048 20408 33100 20417
rect 31944 20340 31996 20392
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 6920 20204 6972 20256
rect 7840 20204 7892 20256
rect 16856 20204 16908 20256
rect 18236 20204 18288 20256
rect 20812 20272 20864 20324
rect 19708 20204 19760 20256
rect 27620 20315 27672 20324
rect 27620 20281 27629 20315
rect 27629 20281 27663 20315
rect 27663 20281 27672 20315
rect 27620 20272 27672 20281
rect 32312 20272 32364 20324
rect 32956 20315 33008 20324
rect 32956 20281 32965 20315
rect 32965 20281 32999 20315
rect 32999 20281 33008 20315
rect 32956 20272 33008 20281
rect 28264 20204 28316 20256
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 3976 20043 4028 20052
rect 3976 20009 3985 20043
rect 3985 20009 4019 20043
rect 4019 20009 4028 20043
rect 3976 20000 4028 20009
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 3240 19907 3292 19916
rect 3240 19873 3249 19907
rect 3249 19873 3283 19907
rect 3283 19873 3292 19907
rect 3240 19864 3292 19873
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3516 19796 3568 19848
rect 3332 19728 3384 19780
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 6920 19932 6972 19984
rect 7104 19975 7156 19984
rect 7104 19941 7113 19975
rect 7113 19941 7147 19975
rect 7147 19941 7156 19975
rect 7104 19932 7156 19941
rect 7656 20000 7708 20052
rect 15660 20000 15712 20052
rect 19248 20000 19300 20052
rect 7748 19975 7800 19984
rect 7748 19941 7757 19975
rect 7757 19941 7791 19975
rect 7791 19941 7800 19975
rect 7748 19932 7800 19941
rect 9220 19932 9272 19984
rect 4252 19771 4304 19780
rect 4252 19737 4261 19771
rect 4261 19737 4295 19771
rect 4295 19737 4304 19771
rect 4252 19728 4304 19737
rect 4896 19728 4948 19780
rect 5080 19771 5132 19780
rect 5080 19737 5089 19771
rect 5089 19737 5123 19771
rect 5123 19737 5132 19771
rect 5080 19728 5132 19737
rect 7380 19796 7432 19848
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 8392 19796 8444 19848
rect 11888 19907 11940 19916
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 14096 19864 14148 19916
rect 7288 19728 7340 19780
rect 9036 19728 9088 19780
rect 9772 19728 9824 19780
rect 10232 19728 10284 19780
rect 10692 19728 10744 19780
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13452 19796 13504 19848
rect 19616 19864 19668 19916
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 16856 19839 16908 19848
rect 16856 19805 16865 19839
rect 16865 19805 16899 19839
rect 16899 19805 16908 19839
rect 16856 19796 16908 19805
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19524 19839 19576 19848
rect 19524 19805 19534 19839
rect 19534 19805 19568 19839
rect 19568 19805 19576 19839
rect 19524 19796 19576 19805
rect 19800 20000 19852 20052
rect 19892 19932 19944 19984
rect 24768 20000 24820 20052
rect 20628 19932 20680 19984
rect 32312 19975 32364 19984
rect 32312 19941 32321 19975
rect 32321 19941 32355 19975
rect 32355 19941 32364 19975
rect 32312 19932 32364 19941
rect 19892 19839 19944 19848
rect 19892 19805 19906 19839
rect 19906 19805 19940 19839
rect 19940 19805 19944 19839
rect 21272 19864 21324 19916
rect 23204 19864 23256 19916
rect 32128 19864 32180 19916
rect 19892 19796 19944 19805
rect 31944 19839 31996 19848
rect 31944 19805 31953 19839
rect 31953 19805 31987 19839
rect 31987 19805 31996 19839
rect 31944 19796 31996 19805
rect 32220 19839 32272 19848
rect 32220 19805 32229 19839
rect 32229 19805 32263 19839
rect 32263 19805 32272 19839
rect 32220 19796 32272 19805
rect 32404 19839 32456 19848
rect 32404 19805 32413 19839
rect 32413 19805 32447 19839
rect 32447 19805 32456 19839
rect 32404 19796 32456 19805
rect 32496 19796 32548 19848
rect 15660 19771 15712 19780
rect 15660 19737 15669 19771
rect 15669 19737 15703 19771
rect 15703 19737 15712 19771
rect 15660 19728 15712 19737
rect 16028 19728 16080 19780
rect 4712 19660 4764 19712
rect 4988 19660 5040 19712
rect 11520 19703 11572 19712
rect 11520 19669 11529 19703
rect 11529 19669 11563 19703
rect 11563 19669 11572 19703
rect 11520 19660 11572 19669
rect 19432 19660 19484 19712
rect 19616 19660 19668 19712
rect 20812 19771 20864 19780
rect 20812 19737 20821 19771
rect 20821 19737 20855 19771
rect 20855 19737 20864 19771
rect 20812 19728 20864 19737
rect 24676 19660 24728 19712
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 1860 19456 1912 19508
rect 5080 19456 5132 19508
rect 19524 19456 19576 19508
rect 20996 19456 21048 19508
rect 29184 19456 29236 19508
rect 32496 19456 32548 19508
rect 33048 19456 33100 19508
rect 2964 19388 3016 19440
rect 3516 19320 3568 19372
rect 12440 19431 12492 19440
rect 12440 19397 12449 19431
rect 12449 19397 12483 19431
rect 12483 19397 12492 19431
rect 12440 19388 12492 19397
rect 15844 19388 15896 19440
rect 16028 19388 16080 19440
rect 4620 19363 4672 19372
rect 4620 19329 4629 19363
rect 4629 19329 4663 19363
rect 4663 19329 4672 19363
rect 4620 19320 4672 19329
rect 6644 19320 6696 19372
rect 6736 19320 6788 19372
rect 7656 19320 7708 19372
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 9772 19320 9824 19372
rect 10324 19320 10376 19372
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 17684 19320 17736 19372
rect 19432 19388 19484 19440
rect 20076 19388 20128 19440
rect 4252 19184 4304 19236
rect 7012 19252 7064 19304
rect 11060 19252 11112 19304
rect 11520 19252 11572 19304
rect 14740 19252 14792 19304
rect 21088 19320 21140 19372
rect 21180 19320 21232 19372
rect 24952 19388 25004 19440
rect 28172 19388 28224 19440
rect 23204 19320 23256 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27896 19320 27948 19372
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 31300 19320 31352 19372
rect 32220 19388 32272 19440
rect 31944 19320 31996 19372
rect 32404 19320 32456 19372
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 28540 19252 28592 19304
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 31392 19227 31444 19236
rect 31392 19193 31401 19227
rect 31401 19193 31435 19227
rect 31435 19193 31444 19227
rect 31392 19184 31444 19193
rect 8576 19116 8628 19168
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 10600 19116 10652 19125
rect 14924 19116 14976 19168
rect 19340 19116 19392 19168
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 14924 18912 14976 18964
rect 16212 18912 16264 18964
rect 18236 18912 18288 18964
rect 19340 18912 19392 18964
rect 2964 18844 3016 18896
rect 7104 18776 7156 18828
rect 8392 18844 8444 18896
rect 19800 18912 19852 18964
rect 20904 18912 20956 18964
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 33324 18912 33376 18964
rect 9128 18776 9180 18828
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 10140 18708 10192 18760
rect 3240 18640 3292 18692
rect 7196 18640 7248 18692
rect 9772 18640 9824 18692
rect 10600 18708 10652 18760
rect 12440 18708 12492 18760
rect 14740 18708 14792 18760
rect 15384 18708 15436 18760
rect 12072 18640 12124 18692
rect 16948 18708 17000 18760
rect 21824 18776 21876 18828
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 15752 18640 15804 18692
rect 19524 18640 19576 18692
rect 20720 18708 20772 18760
rect 23756 18751 23808 18760
rect 23756 18717 23765 18751
rect 23765 18717 23799 18751
rect 23799 18717 23808 18751
rect 23756 18708 23808 18717
rect 19708 18683 19760 18692
rect 19708 18649 19742 18683
rect 19742 18649 19760 18683
rect 25136 18708 25188 18760
rect 27712 18844 27764 18896
rect 27252 18776 27304 18828
rect 29092 18776 29144 18828
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 19708 18640 19760 18649
rect 15200 18572 15252 18624
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 19892 18572 19944 18624
rect 23572 18615 23624 18624
rect 23572 18581 23581 18615
rect 23581 18581 23615 18615
rect 23615 18581 23624 18615
rect 23572 18572 23624 18581
rect 24492 18572 24544 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 25688 18640 25740 18692
rect 27160 18708 27212 18760
rect 27528 18708 27580 18760
rect 27896 18751 27948 18760
rect 27896 18717 27905 18751
rect 27905 18717 27939 18751
rect 27939 18717 27948 18751
rect 27896 18708 27948 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 28632 18708 28684 18760
rect 27344 18683 27396 18692
rect 27344 18649 27353 18683
rect 27353 18649 27387 18683
rect 27387 18649 27396 18683
rect 27344 18640 27396 18649
rect 29276 18708 29328 18760
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 32496 18776 32548 18828
rect 32588 18776 32640 18828
rect 29368 18640 29420 18692
rect 32864 18708 32916 18760
rect 32404 18640 32456 18692
rect 26148 18572 26200 18624
rect 26240 18572 26292 18624
rect 28356 18615 28408 18624
rect 28356 18581 28365 18615
rect 28365 18581 28399 18615
rect 28399 18581 28408 18615
rect 28356 18572 28408 18581
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 9036 18368 9088 18420
rect 15752 18411 15804 18420
rect 15752 18377 15761 18411
rect 15761 18377 15795 18411
rect 15795 18377 15804 18411
rect 15752 18368 15804 18377
rect 16212 18368 16264 18420
rect 19432 18368 19484 18420
rect 19800 18368 19852 18420
rect 25688 18411 25740 18420
rect 25688 18377 25697 18411
rect 25697 18377 25731 18411
rect 25731 18377 25740 18411
rect 25688 18368 25740 18377
rect 32864 18368 32916 18420
rect 6460 18300 6512 18352
rect 12072 18300 12124 18352
rect 6644 18232 6696 18284
rect 8576 18232 8628 18284
rect 9772 18232 9824 18284
rect 11060 18232 11112 18284
rect 11796 18232 11848 18284
rect 12348 18232 12400 18284
rect 14740 18343 14792 18352
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 15844 18300 15896 18352
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 15660 18232 15712 18284
rect 18512 18300 18564 18352
rect 24952 18300 25004 18352
rect 28448 18300 28500 18352
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 24584 18232 24636 18284
rect 25320 18275 25372 18284
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 28356 18232 28408 18284
rect 28724 18275 28776 18284
rect 28724 18241 28733 18275
rect 28733 18241 28767 18275
rect 28767 18241 28776 18275
rect 28724 18232 28776 18241
rect 29092 18275 29144 18284
rect 29092 18241 29101 18275
rect 29101 18241 29135 18275
rect 29135 18241 29144 18275
rect 29092 18232 29144 18241
rect 29184 18232 29236 18284
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 17132 18164 17184 18216
rect 23112 18164 23164 18216
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 27528 18207 27580 18216
rect 27528 18173 27537 18207
rect 27537 18173 27571 18207
rect 27571 18173 27580 18207
rect 27528 18164 27580 18173
rect 29000 18164 29052 18216
rect 32312 18207 32364 18216
rect 32312 18173 32321 18207
rect 32321 18173 32355 18207
rect 32355 18173 32364 18207
rect 32312 18164 32364 18173
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 35072 18164 35124 18216
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 28540 18096 28592 18148
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 18236 18028 18288 18080
rect 25228 18028 25280 18080
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 6736 17824 6788 17876
rect 15384 17824 15436 17876
rect 3516 17756 3568 17808
rect 11612 17688 11664 17740
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 7104 17620 7156 17672
rect 15200 17663 15252 17672
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 17408 17620 17460 17672
rect 2688 17552 2740 17604
rect 12164 17552 12216 17604
rect 12808 17595 12860 17604
rect 12808 17561 12817 17595
rect 12817 17561 12851 17595
rect 12851 17561 12860 17595
rect 12808 17552 12860 17561
rect 16212 17552 16264 17604
rect 19248 17620 19300 17672
rect 21824 17824 21876 17876
rect 27988 17867 28040 17876
rect 27988 17833 27997 17867
rect 27997 17833 28031 17867
rect 28031 17833 28040 17867
rect 27988 17824 28040 17833
rect 29000 17824 29052 17876
rect 23756 17756 23808 17808
rect 24676 17688 24728 17740
rect 25780 17688 25832 17740
rect 27896 17688 27948 17740
rect 25688 17620 25740 17672
rect 27712 17663 27764 17672
rect 27712 17629 27721 17663
rect 27721 17629 27755 17663
rect 27755 17629 27764 17663
rect 27712 17620 27764 17629
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 28540 17620 28592 17672
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 26608 17552 26660 17604
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 10968 17484 11020 17536
rect 12992 17484 13044 17536
rect 16580 17484 16632 17536
rect 17500 17484 17552 17536
rect 20904 17484 20956 17536
rect 24860 17484 24912 17536
rect 25964 17484 26016 17536
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 30932 17663 30984 17672
rect 30932 17629 30941 17663
rect 30941 17629 30975 17663
rect 30975 17629 30984 17663
rect 32312 17756 32364 17808
rect 30932 17620 30984 17629
rect 32588 17663 32640 17672
rect 32588 17629 32597 17663
rect 32597 17629 32631 17663
rect 32631 17629 32640 17663
rect 32588 17620 32640 17629
rect 33416 17663 33468 17672
rect 33416 17629 33425 17663
rect 33425 17629 33459 17663
rect 33459 17629 33468 17663
rect 33416 17620 33468 17629
rect 31116 17595 31168 17604
rect 31116 17561 31125 17595
rect 31125 17561 31159 17595
rect 31159 17561 31168 17595
rect 31116 17552 31168 17561
rect 31944 17484 31996 17536
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 6920 17280 6972 17332
rect 2964 17255 3016 17264
rect 2964 17221 2973 17255
rect 2973 17221 3007 17255
rect 3007 17221 3016 17255
rect 2964 17212 3016 17221
rect 4252 17144 4304 17196
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 6828 17144 6880 17196
rect 7472 17144 7524 17196
rect 7748 17144 7800 17196
rect 9220 17212 9272 17264
rect 10324 17212 10376 17264
rect 12256 17212 12308 17264
rect 13176 17212 13228 17264
rect 18236 17255 18288 17264
rect 18236 17221 18245 17255
rect 18245 17221 18279 17255
rect 18279 17221 18288 17255
rect 18236 17212 18288 17221
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 15384 17144 15436 17196
rect 16672 17144 16724 17196
rect 17224 17144 17276 17196
rect 19800 17255 19852 17264
rect 19800 17221 19809 17255
rect 19809 17221 19843 17255
rect 19843 17221 19852 17255
rect 19800 17212 19852 17221
rect 21180 17212 21232 17264
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 7012 17076 7064 17128
rect 10600 17076 10652 17128
rect 11612 17076 11664 17128
rect 15936 17119 15988 17128
rect 15936 17085 15945 17119
rect 15945 17085 15979 17119
rect 15979 17085 15988 17119
rect 15936 17076 15988 17085
rect 17408 17076 17460 17128
rect 21088 17144 21140 17196
rect 22744 17280 22796 17332
rect 23572 17212 23624 17264
rect 23756 17144 23808 17196
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25044 17144 25096 17153
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 27804 17280 27856 17332
rect 28816 17280 28868 17332
rect 30012 17280 30064 17332
rect 30932 17323 30984 17332
rect 30932 17289 30941 17323
rect 30941 17289 30975 17323
rect 30975 17289 30984 17323
rect 30932 17280 30984 17289
rect 25964 17212 26016 17264
rect 32220 17280 32272 17332
rect 32864 17280 32916 17332
rect 33416 17280 33468 17332
rect 22560 17076 22612 17128
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 6460 17008 6512 17060
rect 10416 17008 10468 17060
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 11152 16940 11204 16992
rect 19340 16940 19392 16992
rect 19524 16940 19576 16992
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 22468 16940 22520 16992
rect 24492 16983 24544 16992
rect 24492 16949 24501 16983
rect 24501 16949 24535 16983
rect 24535 16949 24544 16983
rect 24492 16940 24544 16949
rect 24768 16940 24820 16992
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 28540 17187 28592 17196
rect 28540 17153 28549 17187
rect 28549 17153 28583 17187
rect 28583 17153 28592 17187
rect 28540 17144 28592 17153
rect 28908 17144 28960 17196
rect 26608 17076 26660 17128
rect 30288 17076 30340 17128
rect 31300 17144 31352 17196
rect 31392 17144 31444 17196
rect 32588 17144 32640 17196
rect 32588 16940 32640 16992
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 2688 16736 2740 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 6644 16736 6696 16788
rect 8208 16736 8260 16788
rect 9864 16736 9916 16788
rect 10968 16736 11020 16788
rect 12256 16779 12308 16788
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 21088 16736 21140 16788
rect 25964 16779 26016 16788
rect 25964 16745 25973 16779
rect 25973 16745 26007 16779
rect 26007 16745 26016 16779
rect 25964 16736 26016 16745
rect 31116 16736 31168 16788
rect 32220 16779 32272 16788
rect 32220 16745 32229 16779
rect 32229 16745 32263 16779
rect 32263 16745 32272 16779
rect 32220 16736 32272 16745
rect 2596 16600 2648 16652
rect 6460 16668 6512 16720
rect 8300 16668 8352 16720
rect 12072 16668 12124 16720
rect 15200 16668 15252 16720
rect 17500 16668 17552 16720
rect 7104 16643 7156 16652
rect 7104 16609 7113 16643
rect 7113 16609 7147 16643
rect 7147 16609 7156 16643
rect 7104 16600 7156 16609
rect 3056 16464 3108 16516
rect 6644 16532 6696 16584
rect 9864 16600 9916 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10416 16600 10468 16652
rect 10048 16575 10100 16584
rect 10048 16541 10055 16575
rect 10055 16541 10089 16575
rect 10089 16541 10100 16575
rect 12440 16600 12492 16652
rect 14740 16600 14792 16652
rect 26148 16600 26200 16652
rect 10048 16532 10100 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 15384 16532 15436 16584
rect 16580 16532 16632 16584
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 5080 16464 5132 16516
rect 6552 16464 6604 16516
rect 11152 16464 11204 16516
rect 17040 16464 17092 16516
rect 6368 16396 6420 16448
rect 7104 16396 7156 16448
rect 7656 16396 7708 16448
rect 9680 16396 9732 16448
rect 10140 16396 10192 16448
rect 10416 16396 10468 16448
rect 15384 16396 15436 16448
rect 15936 16396 15988 16448
rect 16120 16396 16172 16448
rect 17408 16464 17460 16516
rect 19524 16532 19576 16584
rect 20444 16532 20496 16584
rect 17684 16396 17736 16448
rect 18696 16507 18748 16516
rect 18696 16473 18705 16507
rect 18705 16473 18739 16507
rect 18739 16473 18748 16507
rect 18696 16464 18748 16473
rect 19248 16464 19300 16516
rect 23296 16532 23348 16584
rect 21640 16464 21692 16516
rect 24584 16575 24636 16584
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 24860 16575 24912 16584
rect 24860 16541 24894 16575
rect 24894 16541 24912 16575
rect 24860 16532 24912 16541
rect 28908 16600 28960 16652
rect 29092 16600 29144 16652
rect 29736 16643 29788 16652
rect 29736 16609 29745 16643
rect 29745 16609 29779 16643
rect 29779 16609 29788 16643
rect 29736 16600 29788 16609
rect 31300 16668 31352 16720
rect 30012 16600 30064 16652
rect 31392 16600 31444 16652
rect 21180 16396 21232 16448
rect 26148 16396 26200 16448
rect 28356 16464 28408 16516
rect 28724 16464 28776 16516
rect 31300 16532 31352 16584
rect 32312 16600 32364 16652
rect 32772 16600 32824 16652
rect 32404 16575 32456 16584
rect 32404 16541 32413 16575
rect 32413 16541 32447 16575
rect 32447 16541 32456 16575
rect 32404 16532 32456 16541
rect 27804 16396 27856 16448
rect 28448 16396 28500 16448
rect 30012 16439 30064 16448
rect 30012 16405 30021 16439
rect 30021 16405 30055 16439
rect 30055 16405 30064 16439
rect 30012 16396 30064 16405
rect 30104 16439 30156 16448
rect 30104 16405 30113 16439
rect 30113 16405 30147 16439
rect 30147 16405 30156 16439
rect 30104 16396 30156 16405
rect 30288 16439 30340 16448
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 6736 16235 6788 16244
rect 6736 16201 6745 16235
rect 6745 16201 6779 16235
rect 6779 16201 6788 16235
rect 6736 16192 6788 16201
rect 12716 16192 12768 16244
rect 5724 16167 5776 16176
rect 5724 16133 5733 16167
rect 5733 16133 5767 16167
rect 5767 16133 5776 16167
rect 5724 16124 5776 16133
rect 6828 16124 6880 16176
rect 6460 16056 6512 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6644 16056 6696 16108
rect 9312 16056 9364 16108
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 19248 16192 19300 16244
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 20536 16192 20588 16244
rect 15200 16167 15252 16176
rect 15200 16133 15234 16167
rect 15234 16133 15252 16167
rect 15200 16124 15252 16133
rect 18236 16167 18288 16176
rect 18236 16133 18245 16167
rect 18245 16133 18279 16167
rect 18279 16133 18288 16167
rect 18236 16124 18288 16133
rect 18696 16124 18748 16176
rect 21180 16124 21232 16176
rect 22652 16235 22704 16244
rect 22652 16201 22661 16235
rect 22661 16201 22695 16235
rect 22695 16201 22704 16235
rect 22652 16192 22704 16201
rect 24492 16192 24544 16244
rect 14372 16056 14424 16108
rect 16212 16056 16264 16108
rect 16580 16056 16632 16108
rect 7104 15988 7156 16040
rect 14740 15988 14792 16040
rect 16396 15988 16448 16040
rect 20260 16056 20312 16108
rect 20168 15988 20220 16040
rect 5540 15920 5592 15972
rect 15936 15920 15988 15972
rect 20904 16099 20956 16108
rect 20904 16065 20949 16099
rect 20949 16065 20956 16099
rect 20904 16056 20956 16065
rect 21824 16056 21876 16108
rect 26056 16124 26108 16176
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22836 16056 22888 16108
rect 25136 16099 25188 16108
rect 25136 16065 25145 16099
rect 25145 16065 25179 16099
rect 25179 16065 25188 16099
rect 25136 16056 25188 16065
rect 26148 16056 26200 16108
rect 26608 16099 26660 16108
rect 26608 16065 26617 16099
rect 26617 16065 26651 16099
rect 26651 16065 26660 16099
rect 26608 16056 26660 16065
rect 27988 15988 28040 16040
rect 28724 16192 28776 16244
rect 32772 16192 32824 16244
rect 28448 16056 28500 16108
rect 30104 16124 30156 16176
rect 28908 16099 28960 16108
rect 28908 16065 28917 16099
rect 28917 16065 28951 16099
rect 28951 16065 28960 16099
rect 28908 16056 28960 16065
rect 29092 16056 29144 16108
rect 30288 16056 30340 16108
rect 32404 16056 32456 16108
rect 33876 16056 33928 16108
rect 32312 16031 32364 16040
rect 32312 15997 32321 16031
rect 32321 15997 32355 16031
rect 32355 15997 32364 16031
rect 32312 15988 32364 15997
rect 26056 15920 26108 15972
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 17040 15852 17092 15904
rect 19432 15852 19484 15904
rect 21640 15852 21692 15904
rect 24584 15852 24636 15904
rect 26148 15895 26200 15904
rect 26148 15861 26157 15895
rect 26157 15861 26191 15895
rect 26191 15861 26200 15895
rect 26148 15852 26200 15861
rect 28172 15852 28224 15904
rect 29460 15895 29512 15904
rect 29460 15861 29469 15895
rect 29469 15861 29503 15895
rect 29503 15861 29512 15895
rect 29460 15852 29512 15861
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 4988 15648 5040 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 11612 15648 11664 15700
rect 23848 15648 23900 15700
rect 25136 15648 25188 15700
rect 26056 15648 26108 15700
rect 27988 15691 28040 15700
rect 27988 15657 27997 15691
rect 27997 15657 28031 15691
rect 28031 15657 28040 15691
rect 27988 15648 28040 15657
rect 31760 15648 31812 15700
rect 32312 15648 32364 15700
rect 33876 15691 33928 15700
rect 33876 15657 33885 15691
rect 33885 15657 33919 15691
rect 33919 15657 33928 15691
rect 33876 15648 33928 15657
rect 13268 15580 13320 15632
rect 15108 15580 15160 15632
rect 22376 15580 22428 15632
rect 32680 15580 32732 15632
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 5080 15444 5132 15496
rect 5816 15444 5868 15496
rect 6644 15512 6696 15564
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 10600 15512 10652 15564
rect 6552 15444 6604 15496
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 2964 15419 3016 15428
rect 2964 15385 2973 15419
rect 2973 15385 3007 15419
rect 3007 15385 3016 15419
rect 2964 15376 3016 15385
rect 5540 15376 5592 15428
rect 7472 15444 7524 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 13452 15512 13504 15564
rect 14372 15444 14424 15496
rect 14556 15444 14608 15496
rect 15660 15444 15712 15496
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16396 15512 16448 15564
rect 19156 15512 19208 15564
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 4436 15308 4488 15360
rect 6092 15308 6144 15360
rect 17592 15376 17644 15428
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 22192 15444 22244 15496
rect 25780 15512 25832 15564
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 29460 15512 29512 15564
rect 19340 15376 19392 15428
rect 21916 15376 21968 15428
rect 24400 15376 24452 15428
rect 27712 15444 27764 15496
rect 28080 15444 28132 15496
rect 28448 15487 28500 15496
rect 28448 15453 28457 15487
rect 28457 15453 28491 15487
rect 28491 15453 28500 15487
rect 28448 15444 28500 15453
rect 25780 15376 25832 15428
rect 29552 15376 29604 15428
rect 32864 15444 32916 15496
rect 32956 15419 33008 15428
rect 32956 15385 32965 15419
rect 32965 15385 32999 15419
rect 32999 15385 33008 15419
rect 32956 15376 33008 15385
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 12532 15308 12584 15360
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 24768 15308 24820 15360
rect 32772 15308 32824 15360
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 5724 15104 5776 15156
rect 8484 15104 8536 15156
rect 9956 15104 10008 15156
rect 2964 15036 3016 15088
rect 5816 15079 5868 15088
rect 5816 15045 5825 15079
rect 5825 15045 5859 15079
rect 5859 15045 5868 15079
rect 5816 15036 5868 15045
rect 16488 15104 16540 15156
rect 17132 15104 17184 15156
rect 12716 15036 12768 15088
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2688 14900 2740 14952
rect 3240 14832 3292 14884
rect 4528 14968 4580 15020
rect 9956 14968 10008 15020
rect 10324 14968 10376 15020
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 15660 14968 15712 15020
rect 16856 14968 16908 15020
rect 17684 15036 17736 15088
rect 12072 14900 12124 14952
rect 16580 14900 16632 14952
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 22468 15104 22520 15156
rect 32956 15104 33008 15156
rect 23940 15036 23992 15088
rect 24768 15036 24820 15088
rect 30840 15036 30892 15088
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 22192 15011 22244 15020
rect 22192 14977 22201 15011
rect 22201 14977 22235 15011
rect 22235 14977 22244 15011
rect 22192 14968 22244 14977
rect 25136 15011 25188 15020
rect 25136 14977 25154 15011
rect 25154 14977 25188 15011
rect 25136 14968 25188 14977
rect 29000 14968 29052 15020
rect 29920 14968 29972 15020
rect 13268 14832 13320 14884
rect 26424 14900 26476 14952
rect 24400 14832 24452 14884
rect 29644 14875 29696 14884
rect 29644 14841 29653 14875
rect 29653 14841 29687 14875
rect 29687 14841 29696 14875
rect 29644 14832 29696 14841
rect 4252 14764 4304 14816
rect 6552 14764 6604 14816
rect 11980 14764 12032 14816
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 20996 14764 21048 14816
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 6828 14560 6880 14612
rect 6092 14492 6144 14544
rect 9128 14560 9180 14612
rect 19892 14560 19944 14612
rect 8484 14535 8536 14544
rect 8484 14501 8493 14535
rect 8493 14501 8527 14535
rect 8527 14501 8536 14535
rect 8484 14492 8536 14501
rect 8852 14492 8904 14544
rect 9312 14492 9364 14544
rect 1768 14424 1820 14476
rect 20260 14492 20312 14544
rect 22468 14560 22520 14612
rect 25964 14603 26016 14612
rect 25964 14569 25973 14603
rect 25973 14569 26007 14603
rect 26007 14569 26016 14603
rect 25964 14560 26016 14569
rect 22192 14492 22244 14544
rect 23756 14492 23808 14544
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 3056 14356 3108 14408
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 5724 14288 5776 14340
rect 8116 14356 8168 14408
rect 6460 14288 6512 14340
rect 7104 14288 7156 14340
rect 7472 14288 7524 14340
rect 7932 14331 7984 14340
rect 7932 14297 7941 14331
rect 7941 14297 7975 14331
rect 7975 14297 7984 14331
rect 7932 14288 7984 14297
rect 3792 14220 3844 14272
rect 5816 14220 5868 14272
rect 6920 14220 6972 14272
rect 7840 14220 7892 14272
rect 8576 14288 8628 14340
rect 9220 14356 9272 14408
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 9496 14331 9548 14340
rect 9496 14297 9505 14331
rect 9505 14297 9539 14331
rect 9539 14297 9548 14331
rect 9496 14288 9548 14297
rect 10692 14288 10744 14340
rect 12440 14288 12492 14340
rect 13728 14356 13780 14408
rect 20536 14424 20588 14476
rect 24584 14467 24636 14476
rect 24584 14433 24593 14467
rect 24593 14433 24627 14467
rect 24627 14433 24636 14467
rect 24584 14424 24636 14433
rect 31760 14424 31812 14476
rect 32312 14424 32364 14476
rect 17592 14356 17644 14408
rect 18420 14356 18472 14408
rect 19708 14356 19760 14408
rect 20996 14399 21048 14408
rect 20996 14365 21030 14399
rect 21030 14365 21048 14399
rect 20996 14356 21048 14365
rect 26148 14356 26200 14408
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 26976 14356 27028 14408
rect 27528 14356 27580 14408
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 30104 14356 30156 14408
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32128 14356 32180 14365
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 19340 14288 19392 14340
rect 19524 14288 19576 14340
rect 22744 14288 22796 14340
rect 29736 14331 29788 14340
rect 29736 14297 29745 14331
rect 29745 14297 29779 14331
rect 29779 14297 29788 14331
rect 29736 14288 29788 14297
rect 10232 14220 10284 14272
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 19892 14220 19944 14272
rect 23848 14220 23900 14272
rect 27804 14263 27856 14272
rect 27804 14229 27813 14263
rect 27813 14229 27847 14263
rect 27847 14229 27856 14263
rect 27804 14220 27856 14229
rect 31300 14220 31352 14272
rect 33232 14263 33284 14272
rect 33232 14229 33241 14263
rect 33241 14229 33275 14263
rect 33275 14229 33284 14263
rect 33232 14220 33284 14229
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 1676 14016 1728 14068
rect 7932 14016 7984 14068
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 6460 13948 6512 14000
rect 3056 13880 3108 13932
rect 4068 13880 4120 13932
rect 5540 13880 5592 13932
rect 5816 13880 5868 13932
rect 7104 13948 7156 14000
rect 12440 14016 12492 14068
rect 12808 14016 12860 14068
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 5080 13812 5132 13864
rect 8300 13880 8352 13932
rect 9220 13880 9272 13932
rect 11980 13948 12032 14000
rect 13084 13948 13136 14000
rect 13728 13880 13780 13932
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 19892 14016 19944 14068
rect 20812 14016 20864 14068
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 15936 13880 15988 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 8392 13812 8444 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 8576 13744 8628 13796
rect 10324 13744 10376 13796
rect 17684 13880 17736 13932
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 19064 13991 19116 14000
rect 19064 13957 19073 13991
rect 19073 13957 19107 13991
rect 19107 13957 19116 13991
rect 19064 13948 19116 13957
rect 20444 13948 20496 14000
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 21180 14016 21232 14068
rect 22284 14016 22336 14068
rect 24032 14016 24084 14068
rect 25136 14016 25188 14068
rect 26608 14016 26660 14068
rect 27528 14016 27580 14068
rect 27712 13991 27764 14000
rect 27712 13957 27721 13991
rect 27721 13957 27755 13991
rect 27755 13957 27764 13991
rect 27712 13948 27764 13957
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 22468 13880 22520 13932
rect 23296 13923 23348 13932
rect 23296 13889 23305 13923
rect 23305 13889 23339 13923
rect 23339 13889 23348 13923
rect 23296 13880 23348 13889
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 24768 13880 24820 13932
rect 26792 13880 26844 13932
rect 27620 13923 27672 13932
rect 27620 13889 27629 13923
rect 27629 13889 27663 13923
rect 27663 13889 27672 13923
rect 27620 13880 27672 13889
rect 28080 14016 28132 14068
rect 29920 14016 29972 14068
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 30840 14016 30892 14068
rect 31300 14016 31352 14068
rect 32588 14016 32640 14068
rect 27988 13948 28040 14000
rect 28172 13880 28224 13932
rect 28908 13880 28960 13932
rect 2964 13676 3016 13728
rect 4252 13676 4304 13728
rect 6828 13676 6880 13728
rect 13452 13676 13504 13728
rect 23848 13812 23900 13864
rect 25780 13812 25832 13864
rect 26884 13812 26936 13864
rect 28632 13812 28684 13864
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 29736 13923 29788 13932
rect 29736 13889 29745 13923
rect 29745 13889 29779 13923
rect 29779 13889 29788 13923
rect 29736 13880 29788 13889
rect 27620 13744 27672 13796
rect 28172 13744 28224 13796
rect 28356 13744 28408 13796
rect 30380 13744 30432 13796
rect 19892 13676 19944 13728
rect 20904 13676 20956 13728
rect 28908 13719 28960 13728
rect 28908 13685 28917 13719
rect 28917 13685 28951 13719
rect 28951 13685 28960 13719
rect 28908 13676 28960 13685
rect 31392 13880 31444 13932
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 32772 13676 32824 13728
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 4160 13472 4212 13524
rect 2596 13404 2648 13456
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 3884 13268 3936 13320
rect 5264 13336 5316 13388
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 5632 13472 5684 13524
rect 10876 13472 10928 13524
rect 15660 13515 15712 13524
rect 15660 13481 15669 13515
rect 15669 13481 15703 13515
rect 15703 13481 15712 13515
rect 15660 13472 15712 13481
rect 26976 13472 27028 13524
rect 32312 13472 32364 13524
rect 14556 13404 14608 13456
rect 17592 13404 17644 13456
rect 5080 13268 5132 13320
rect 8484 13336 8536 13388
rect 9036 13336 9088 13388
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 3976 13200 4028 13252
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 3240 13132 3292 13184
rect 8576 13243 8628 13252
rect 8576 13209 8585 13243
rect 8585 13209 8619 13243
rect 8619 13209 8628 13243
rect 8576 13200 8628 13209
rect 9864 13200 9916 13252
rect 8944 13132 8996 13184
rect 15384 13336 15436 13388
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 16856 13336 16908 13388
rect 12072 13243 12124 13252
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 14096 13200 14148 13252
rect 13084 13132 13136 13184
rect 15752 13268 15804 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 19616 13336 19668 13388
rect 22836 13336 22888 13388
rect 28080 13336 28132 13388
rect 18328 13268 18380 13320
rect 19800 13268 19852 13320
rect 26056 13311 26108 13320
rect 26056 13277 26065 13311
rect 26065 13277 26099 13311
rect 26099 13277 26108 13311
rect 26056 13268 26108 13277
rect 32956 13311 33008 13320
rect 32956 13277 32965 13311
rect 32965 13277 32999 13311
rect 32999 13277 33008 13311
rect 32956 13268 33008 13277
rect 15568 13200 15620 13252
rect 20352 13200 20404 13252
rect 15936 13132 15988 13184
rect 18236 13132 18288 13184
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 2596 12928 2648 12980
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 3976 12928 4028 12980
rect 9128 12928 9180 12980
rect 17500 12928 17552 12980
rect 3056 12860 3108 12912
rect 8576 12860 8628 12912
rect 4068 12792 4120 12844
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 11796 12860 11848 12912
rect 12992 12903 13044 12912
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 14740 12903 14792 12912
rect 14740 12869 14749 12903
rect 14749 12869 14783 12903
rect 14783 12869 14792 12903
rect 14740 12860 14792 12869
rect 18420 12860 18472 12912
rect 15200 12792 15252 12844
rect 15568 12792 15620 12844
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 5816 12724 5868 12776
rect 8852 12724 8904 12776
rect 16396 12792 16448 12844
rect 17592 12835 17644 12844
rect 10876 12656 10928 12708
rect 12992 12656 13044 12708
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 19432 12860 19484 12912
rect 19892 12928 19944 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 16120 12724 16172 12733
rect 17224 12724 17276 12776
rect 19800 12792 19852 12844
rect 20352 12792 20404 12844
rect 19616 12724 19668 12776
rect 7564 12588 7616 12640
rect 14372 12588 14424 12640
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 24768 12860 24820 12912
rect 22468 12724 22520 12776
rect 26700 12792 26752 12844
rect 27804 12928 27856 12980
rect 28448 12928 28500 12980
rect 32128 12928 32180 12980
rect 33232 12928 33284 12980
rect 27988 12860 28040 12912
rect 23756 12724 23808 12776
rect 28356 12792 28408 12844
rect 28724 12835 28776 12844
rect 28724 12801 28733 12835
rect 28733 12801 28767 12835
rect 28767 12801 28776 12835
rect 28724 12792 28776 12801
rect 29644 12792 29696 12844
rect 31944 12792 31996 12844
rect 32864 12792 32916 12844
rect 30196 12724 30248 12776
rect 27712 12656 27764 12708
rect 19984 12588 20036 12640
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 25780 12588 25832 12640
rect 28908 12656 28960 12708
rect 28356 12631 28408 12640
rect 28356 12597 28365 12631
rect 28365 12597 28399 12631
rect 28399 12597 28408 12631
rect 28356 12588 28408 12597
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 19800 12384 19852 12436
rect 21916 12384 21968 12436
rect 22560 12384 22612 12436
rect 15936 12316 15988 12368
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 14372 12180 14424 12232
rect 14740 12180 14792 12232
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 15752 12180 15804 12232
rect 19340 12316 19392 12368
rect 19708 12316 19760 12368
rect 21824 12316 21876 12368
rect 24676 12384 24728 12436
rect 28540 12384 28592 12436
rect 25688 12316 25740 12368
rect 27896 12316 27948 12368
rect 16856 12180 16908 12232
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 18052 12248 18104 12300
rect 21088 12248 21140 12300
rect 16580 12112 16632 12164
rect 17224 12112 17276 12164
rect 18696 12112 18748 12164
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 20904 12180 20956 12232
rect 21548 12180 21600 12232
rect 22744 12180 22796 12232
rect 20536 12112 20588 12164
rect 24584 12180 24636 12232
rect 24676 12180 24728 12232
rect 28172 12223 28224 12232
rect 28172 12189 28176 12223
rect 28176 12189 28210 12223
rect 28210 12189 28224 12223
rect 20628 12044 20680 12096
rect 24032 12112 24084 12164
rect 28172 12180 28224 12189
rect 28724 12248 28776 12300
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 24768 12044 24820 12096
rect 28448 12112 28500 12164
rect 30380 12112 30432 12164
rect 31392 12112 31444 12164
rect 31208 12044 31260 12096
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 22376 11883 22428 11892
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 13452 11704 13504 11756
rect 15200 11772 15252 11824
rect 15752 11815 15804 11824
rect 15752 11781 15761 11815
rect 15761 11781 15795 11815
rect 15795 11781 15804 11815
rect 15752 11772 15804 11781
rect 14556 11747 14608 11756
rect 14556 11713 14565 11747
rect 14565 11713 14599 11747
rect 14599 11713 14608 11747
rect 14556 11704 14608 11713
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 18328 11704 18380 11756
rect 20904 11704 20956 11756
rect 22744 11815 22796 11824
rect 22744 11781 22753 11815
rect 22753 11781 22787 11815
rect 22787 11781 22796 11815
rect 22744 11772 22796 11781
rect 23480 11772 23532 11824
rect 24584 11772 24636 11824
rect 24768 11840 24820 11892
rect 25320 11840 25372 11892
rect 28448 11840 28500 11892
rect 28724 11883 28776 11892
rect 28724 11849 28733 11883
rect 28733 11849 28767 11883
rect 28767 11849 28776 11883
rect 28724 11840 28776 11849
rect 31208 11883 31260 11892
rect 31208 11849 31217 11883
rect 31217 11849 31251 11883
rect 31251 11849 31260 11883
rect 31208 11840 31260 11849
rect 32680 11883 32732 11892
rect 32680 11849 32689 11883
rect 32689 11849 32723 11883
rect 32723 11849 32732 11883
rect 32680 11840 32732 11849
rect 33692 11840 33744 11892
rect 25136 11772 25188 11824
rect 25688 11815 25740 11824
rect 25688 11781 25697 11815
rect 25697 11781 25731 11815
rect 25731 11781 25740 11815
rect 25688 11772 25740 11781
rect 28356 11772 28408 11824
rect 19800 11636 19852 11688
rect 19984 11636 20036 11688
rect 23664 11704 23716 11756
rect 27896 11704 27948 11756
rect 30196 11704 30248 11756
rect 31392 11747 31444 11756
rect 31392 11713 31401 11747
rect 31401 11713 31435 11747
rect 31435 11713 31444 11747
rect 31392 11704 31444 11713
rect 21364 11568 21416 11620
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 27344 11679 27396 11688
rect 27344 11645 27353 11679
rect 27353 11645 27387 11679
rect 27387 11645 27396 11679
rect 27344 11636 27396 11645
rect 28540 11636 28592 11688
rect 33416 11704 33468 11756
rect 32496 11568 32548 11620
rect 17868 11500 17920 11552
rect 22468 11500 22520 11552
rect 25320 11500 25372 11552
rect 25780 11500 25832 11552
rect 26056 11543 26108 11552
rect 26056 11509 26065 11543
rect 26065 11509 26099 11543
rect 26099 11509 26108 11543
rect 26056 11500 26108 11509
rect 32404 11500 32456 11552
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 4528 11296 4580 11348
rect 20628 11296 20680 11348
rect 20904 11296 20956 11348
rect 21088 11296 21140 11348
rect 26792 11296 26844 11348
rect 31208 11296 31260 11348
rect 17868 11271 17920 11280
rect 17868 11237 17877 11271
rect 17877 11237 17911 11271
rect 17911 11237 17920 11271
rect 17868 11228 17920 11237
rect 19892 11228 19944 11280
rect 12348 11160 12400 11212
rect 17040 11160 17092 11212
rect 5080 11092 5132 11144
rect 7196 11092 7248 11144
rect 11060 11092 11112 11144
rect 11980 11092 12032 11144
rect 12532 11092 12584 11144
rect 12900 11092 12952 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13268 11092 13320 11144
rect 3976 11067 4028 11076
rect 3976 11033 3985 11067
rect 3985 11033 4019 11067
rect 4019 11033 4028 11067
rect 3976 11024 4028 11033
rect 4252 11024 4304 11076
rect 5816 11067 5868 11076
rect 5816 11033 5850 11067
rect 5850 11033 5868 11067
rect 5816 11024 5868 11033
rect 11152 11024 11204 11076
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 7288 10956 7340 11008
rect 7840 10956 7892 11008
rect 9220 10956 9272 11008
rect 12440 11024 12492 11076
rect 12624 11067 12676 11076
rect 12624 11033 12633 11067
rect 12633 11033 12667 11067
rect 12667 11033 12676 11067
rect 12624 11024 12676 11033
rect 13176 11024 13228 11076
rect 12808 10956 12860 11008
rect 12992 10956 13044 11008
rect 13268 10956 13320 11008
rect 16672 11024 16724 11076
rect 17224 11092 17276 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 18328 11092 18380 11144
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 23664 11228 23716 11280
rect 20352 11135 20404 11144
rect 20352 11101 20366 11135
rect 20366 11101 20400 11135
rect 20400 11101 20404 11135
rect 20352 11092 20404 11101
rect 20720 11092 20772 11144
rect 21916 11160 21968 11212
rect 24676 11228 24728 11280
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 21548 11092 21600 11144
rect 23756 11135 23808 11144
rect 23756 11101 23765 11135
rect 23765 11101 23799 11135
rect 23799 11101 23808 11135
rect 23756 11092 23808 11101
rect 25964 11160 26016 11212
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 29552 11092 29604 11144
rect 29828 11092 29880 11144
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 24860 11024 24912 11076
rect 32312 11024 32364 11076
rect 32496 11067 32548 11076
rect 32496 11033 32514 11067
rect 32514 11033 32548 11067
rect 32496 11024 32548 11033
rect 26608 10956 26660 11008
rect 29000 10956 29052 11008
rect 30104 10999 30156 11008
rect 30104 10965 30113 10999
rect 30113 10965 30147 10999
rect 30147 10965 30156 10999
rect 30104 10956 30156 10965
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 6644 10752 6696 10804
rect 3332 10684 3384 10736
rect 2780 10616 2832 10668
rect 3792 10616 3844 10668
rect 6736 10684 6788 10736
rect 6920 10684 6972 10736
rect 7288 10684 7340 10736
rect 7564 10727 7616 10736
rect 7564 10693 7573 10727
rect 7573 10693 7607 10727
rect 7607 10693 7616 10727
rect 7564 10684 7616 10693
rect 4252 10616 4304 10668
rect 8208 10752 8260 10804
rect 8944 10752 8996 10804
rect 8852 10727 8904 10736
rect 8852 10693 8861 10727
rect 8861 10693 8895 10727
rect 8895 10693 8904 10727
rect 8852 10684 8904 10693
rect 9496 10684 9548 10736
rect 10324 10752 10376 10804
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 12716 10752 12768 10804
rect 25964 10795 26016 10804
rect 25964 10761 25973 10795
rect 25973 10761 26007 10795
rect 26007 10761 26016 10795
rect 25964 10752 26016 10761
rect 29092 10752 29144 10804
rect 30104 10752 30156 10804
rect 33692 10795 33744 10804
rect 33692 10761 33701 10795
rect 33701 10761 33735 10795
rect 33735 10761 33744 10795
rect 33692 10752 33744 10761
rect 12900 10727 12952 10736
rect 12900 10693 12909 10727
rect 12909 10693 12943 10727
rect 12943 10693 12952 10727
rect 12900 10684 12952 10693
rect 13452 10684 13504 10736
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 19984 10727 20036 10736
rect 19984 10693 19993 10727
rect 19993 10693 20027 10727
rect 20027 10693 20036 10727
rect 19984 10684 20036 10693
rect 24860 10727 24912 10736
rect 24860 10693 24894 10727
rect 24894 10693 24912 10727
rect 24860 10684 24912 10693
rect 29000 10684 29052 10736
rect 29368 10727 29420 10736
rect 29368 10693 29377 10727
rect 29377 10693 29411 10727
rect 29411 10693 29420 10727
rect 29368 10684 29420 10693
rect 9220 10616 9272 10625
rect 12440 10616 12492 10668
rect 28172 10616 28224 10668
rect 28724 10616 28776 10668
rect 32404 10616 32456 10668
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 3424 10548 3476 10600
rect 6644 10548 6696 10600
rect 9864 10548 9916 10600
rect 12348 10548 12400 10600
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 27344 10591 27396 10600
rect 27344 10557 27353 10591
rect 27353 10557 27387 10591
rect 27387 10557 27396 10591
rect 27344 10548 27396 10557
rect 32312 10591 32364 10600
rect 32312 10557 32321 10591
rect 32321 10557 32355 10591
rect 32355 10557 32364 10591
rect 32312 10548 32364 10557
rect 3240 10480 3292 10532
rect 4252 10480 4304 10532
rect 3608 10412 3660 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 10140 10455 10192 10464
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 14464 10412 14516 10464
rect 29184 10412 29236 10464
rect 30840 10412 30892 10464
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 2780 10208 2832 10260
rect 4528 10208 4580 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 9128 10208 9180 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 23848 10208 23900 10260
rect 24584 10208 24636 10260
rect 25412 10208 25464 10260
rect 27344 10251 27396 10260
rect 27344 10217 27353 10251
rect 27353 10217 27387 10251
rect 27387 10217 27396 10251
rect 27344 10208 27396 10217
rect 28264 10251 28316 10260
rect 28264 10217 28273 10251
rect 28273 10217 28307 10251
rect 28307 10217 28316 10251
rect 28264 10208 28316 10217
rect 28448 10208 28500 10260
rect 29920 10208 29972 10260
rect 2964 10140 3016 10192
rect 4252 10072 4304 10124
rect 7196 10115 7248 10124
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 11060 10072 11112 10124
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4344 10004 4396 10056
rect 3148 9936 3200 9988
rect 4068 9936 4120 9988
rect 3792 9868 3844 9920
rect 5908 10004 5960 10056
rect 12072 10004 12124 10056
rect 25136 10047 25188 10056
rect 25136 10013 25140 10047
rect 25140 10013 25174 10047
rect 25174 10013 25188 10047
rect 5816 9936 5868 9988
rect 7472 9979 7524 9988
rect 7472 9945 7506 9979
rect 7506 9945 7524 9979
rect 7472 9936 7524 9945
rect 9036 9936 9088 9988
rect 25136 10004 25188 10013
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 28540 10072 28592 10124
rect 25228 9979 25280 9988
rect 25228 9945 25237 9979
rect 25237 9945 25271 9979
rect 25271 9945 25280 9979
rect 25228 9936 25280 9945
rect 25964 9936 26016 9988
rect 26608 10004 26660 10056
rect 27712 10004 27764 10056
rect 28448 10004 28500 10056
rect 29092 10072 29144 10124
rect 28908 10047 28960 10056
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10004 28960 10013
rect 32312 10208 32364 10260
rect 30380 10072 30432 10124
rect 30932 10072 30984 10124
rect 28724 9936 28776 9988
rect 30288 10047 30340 10056
rect 30288 10013 30297 10047
rect 30297 10013 30331 10047
rect 30331 10013 30340 10047
rect 30288 10004 30340 10013
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33416 10004 33468 10013
rect 29092 9868 29144 9920
rect 31208 9979 31260 9988
rect 31208 9945 31217 9979
rect 31217 9945 31251 9979
rect 31251 9945 31260 9979
rect 31208 9936 31260 9945
rect 33692 9868 33744 9920
rect 33876 9911 33928 9920
rect 33876 9877 33885 9911
rect 33885 9877 33919 9911
rect 33919 9877 33928 9911
rect 33876 9868 33928 9877
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 2964 9664 3016 9716
rect 4344 9664 4396 9716
rect 8852 9664 8904 9716
rect 28908 9664 28960 9716
rect 3148 9528 3200 9580
rect 3516 9528 3568 9580
rect 2780 9460 2832 9512
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 2688 9392 2740 9444
rect 3240 9392 3292 9444
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 4252 9528 4304 9580
rect 4068 9392 4120 9444
rect 5908 9596 5960 9648
rect 4528 9571 4580 9580
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4528 9528 4580 9537
rect 7472 9571 7524 9580
rect 7472 9537 7506 9571
rect 7506 9537 7524 9571
rect 7472 9528 7524 9537
rect 12072 9596 12124 9648
rect 16212 9596 16264 9648
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17224 9639 17276 9648
rect 17224 9605 17233 9639
rect 17233 9605 17267 9639
rect 17267 9605 17276 9639
rect 17224 9596 17276 9605
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17776 9528 17828 9580
rect 10784 9460 10836 9512
rect 17868 9460 17920 9512
rect 19800 9571 19852 9580
rect 19800 9537 19809 9571
rect 19809 9537 19843 9571
rect 19843 9537 19852 9571
rect 19800 9528 19852 9537
rect 21272 9596 21324 9648
rect 25136 9596 25188 9648
rect 30840 9596 30892 9648
rect 20812 9528 20864 9580
rect 21088 9571 21140 9580
rect 21088 9537 21102 9571
rect 21102 9537 21136 9571
rect 21136 9537 21140 9571
rect 21088 9528 21140 9537
rect 5080 9392 5132 9444
rect 12808 9392 12860 9444
rect 16028 9392 16080 9444
rect 18604 9392 18656 9444
rect 19892 9392 19944 9444
rect 20996 9460 21048 9512
rect 21180 9392 21232 9444
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 17592 9324 17644 9376
rect 19340 9324 19392 9376
rect 21364 9324 21416 9376
rect 22468 9571 22520 9580
rect 22468 9537 22477 9571
rect 22477 9537 22511 9571
rect 22511 9537 22520 9571
rect 22468 9528 22520 9537
rect 25964 9528 26016 9580
rect 28724 9528 28776 9580
rect 30196 9528 30248 9580
rect 31300 9571 31352 9580
rect 31300 9537 31312 9571
rect 31312 9537 31346 9571
rect 31346 9537 31352 9571
rect 31300 9528 31352 9537
rect 31392 9571 31444 9580
rect 31392 9537 31401 9571
rect 31401 9537 31435 9571
rect 31435 9537 31444 9571
rect 31392 9528 31444 9537
rect 31484 9528 31536 9580
rect 23756 9392 23808 9444
rect 31392 9392 31444 9444
rect 31944 9392 31996 9444
rect 25044 9324 25096 9376
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 12532 9120 12584 9172
rect 17224 9120 17276 9172
rect 17684 9120 17736 9172
rect 17316 9052 17368 9104
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 3608 8916 3660 8968
rect 4344 8916 4396 8968
rect 16856 8916 16908 8968
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 19616 9120 19668 9172
rect 19340 9052 19392 9104
rect 21272 9163 21324 9172
rect 21272 9129 21281 9163
rect 21281 9129 21315 9163
rect 21315 9129 21324 9163
rect 21272 9120 21324 9129
rect 21548 9120 21600 9172
rect 22468 9120 22520 9172
rect 33692 9163 33744 9172
rect 33692 9129 33701 9163
rect 33701 9129 33735 9163
rect 33735 9129 33744 9163
rect 33692 9120 33744 9129
rect 22744 9052 22796 9104
rect 2872 8848 2924 8900
rect 11152 8848 11204 8900
rect 15384 8848 15436 8900
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 18420 8848 18472 8900
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 16672 8780 16724 8832
rect 17868 8780 17920 8832
rect 18788 8848 18840 8900
rect 19984 8916 20036 8968
rect 21364 8916 21416 8968
rect 20628 8780 20680 8832
rect 20996 8848 21048 8900
rect 26700 8984 26752 9036
rect 24032 8916 24084 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 27620 8916 27672 8968
rect 29828 8984 29880 9036
rect 29000 8916 29052 8968
rect 30196 8916 30248 8968
rect 32312 8959 32364 8968
rect 32312 8925 32321 8959
rect 32321 8925 32355 8959
rect 32355 8925 32364 8959
rect 32312 8916 32364 8925
rect 33876 8916 33928 8968
rect 26056 8848 26108 8900
rect 21088 8780 21140 8832
rect 23664 8780 23716 8832
rect 24952 8780 25004 8832
rect 28724 8823 28776 8832
rect 28724 8789 28733 8823
rect 28733 8789 28767 8823
rect 28767 8789 28776 8823
rect 28724 8780 28776 8789
rect 29092 8823 29144 8832
rect 29092 8789 29101 8823
rect 29101 8789 29135 8823
rect 29135 8789 29144 8823
rect 29092 8780 29144 8789
rect 29736 8780 29788 8832
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 3516 8576 3568 8628
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 16580 8576 16632 8628
rect 17684 8576 17736 8628
rect 18420 8576 18472 8628
rect 9312 8508 9364 8560
rect 3240 8440 3292 8492
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 18328 8508 18380 8560
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 16212 8440 16264 8492
rect 16672 8440 16724 8492
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 20536 8508 20588 8560
rect 20628 8551 20680 8560
rect 20628 8517 20637 8551
rect 20637 8517 20671 8551
rect 20671 8517 20680 8551
rect 20628 8508 20680 8517
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 21180 8576 21232 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 23756 8576 23808 8628
rect 22468 8508 22520 8560
rect 22560 8508 22612 8560
rect 16488 8372 16540 8424
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 21088 8440 21140 8492
rect 15292 8304 15344 8356
rect 15844 8347 15896 8356
rect 15844 8313 15853 8347
rect 15853 8313 15887 8347
rect 15887 8313 15896 8347
rect 15844 8304 15896 8313
rect 16028 8304 16080 8356
rect 19800 8304 19852 8356
rect 24676 8508 24728 8560
rect 25228 8576 25280 8628
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 31392 8576 31444 8628
rect 24952 8440 25004 8492
rect 30012 8508 30064 8560
rect 30288 8508 30340 8560
rect 31760 8508 31812 8560
rect 26056 8440 26108 8492
rect 28172 8440 28224 8492
rect 28908 8440 28960 8492
rect 30380 8483 30432 8492
rect 30380 8449 30389 8483
rect 30389 8449 30423 8483
rect 30423 8449 30432 8483
rect 30380 8440 30432 8449
rect 31300 8440 31352 8492
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 32312 8415 32364 8424
rect 32312 8381 32321 8415
rect 32321 8381 32355 8415
rect 32355 8381 32364 8415
rect 32312 8372 32364 8381
rect 24032 8304 24084 8356
rect 25136 8304 25188 8356
rect 8300 8236 8352 8288
rect 9864 8236 9916 8288
rect 15200 8279 15252 8288
rect 15200 8245 15209 8279
rect 15209 8245 15243 8279
rect 15243 8245 15252 8279
rect 15200 8236 15252 8245
rect 19064 8236 19116 8288
rect 20628 8236 20680 8288
rect 27896 8236 27948 8288
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 22560 8032 22612 8084
rect 26884 8032 26936 8084
rect 29184 8032 29236 8084
rect 32312 8032 32364 8084
rect 23388 7964 23440 8016
rect 3056 7828 3108 7880
rect 8300 7896 8352 7948
rect 3608 7760 3660 7812
rect 4068 7760 4120 7812
rect 8208 7828 8260 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10600 7828 10652 7880
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 21548 7896 21600 7948
rect 19984 7828 20036 7880
rect 24032 7828 24084 7880
rect 31208 7871 31260 7880
rect 31208 7837 31217 7871
rect 31217 7837 31251 7871
rect 31251 7837 31260 7871
rect 31208 7828 31260 7837
rect 7380 7803 7432 7812
rect 7380 7769 7389 7803
rect 7389 7769 7423 7803
rect 7423 7769 7432 7803
rect 7380 7760 7432 7769
rect 10232 7760 10284 7812
rect 16304 7760 16356 7812
rect 19708 7760 19760 7812
rect 20536 7760 20588 7812
rect 22928 7760 22980 7812
rect 28816 7760 28868 7812
rect 29368 7760 29420 7812
rect 29920 7803 29972 7812
rect 29920 7769 29929 7803
rect 29929 7769 29963 7803
rect 29963 7769 29972 7803
rect 29920 7760 29972 7769
rect 18880 7692 18932 7744
rect 28356 7692 28408 7744
rect 30564 7692 30616 7744
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 15384 7488 15436 7540
rect 5816 7420 5868 7472
rect 6828 7463 6880 7472
rect 6828 7429 6837 7463
rect 6837 7429 6871 7463
rect 6871 7429 6880 7463
rect 6828 7420 6880 7429
rect 7380 7420 7432 7472
rect 10232 7420 10284 7472
rect 11152 7420 11204 7472
rect 16212 7488 16264 7540
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 21088 7488 21140 7540
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 27896 7488 27948 7540
rect 28172 7531 28224 7540
rect 28172 7497 28181 7531
rect 28181 7497 28215 7531
rect 28215 7497 28224 7531
rect 28172 7488 28224 7497
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 3884 7352 3936 7404
rect 8392 7284 8444 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 17408 7420 17460 7472
rect 18236 7463 18288 7472
rect 18236 7429 18245 7463
rect 18245 7429 18279 7463
rect 18279 7429 18288 7463
rect 18236 7420 18288 7429
rect 18880 7420 18932 7472
rect 19984 7463 20036 7472
rect 19984 7429 19993 7463
rect 19993 7429 20027 7463
rect 20027 7429 20036 7463
rect 19984 7420 20036 7429
rect 20904 7463 20956 7472
rect 20904 7429 20913 7463
rect 20913 7429 20947 7463
rect 20947 7429 20956 7463
rect 20904 7420 20956 7429
rect 23388 7463 23440 7472
rect 23388 7429 23397 7463
rect 23397 7429 23431 7463
rect 23431 7429 23440 7463
rect 23388 7420 23440 7429
rect 24860 7420 24912 7472
rect 15200 7352 15252 7404
rect 16948 7352 17000 7404
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 30564 7463 30616 7472
rect 30564 7429 30573 7463
rect 30573 7429 30607 7463
rect 30607 7429 30616 7463
rect 30564 7420 30616 7429
rect 27620 7284 27672 7336
rect 29000 7352 29052 7404
rect 28816 7327 28868 7336
rect 28816 7293 28825 7327
rect 28825 7293 28859 7327
rect 28859 7293 28868 7327
rect 28816 7284 28868 7293
rect 12900 7216 12952 7268
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 8392 7148 8444 7200
rect 10784 7148 10836 7200
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 20628 7148 20680 7200
rect 25596 7191 25648 7200
rect 25596 7157 25605 7191
rect 25605 7157 25639 7191
rect 25639 7157 25648 7191
rect 25596 7148 25648 7157
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 2504 6944 2556 6996
rect 2596 6944 2648 6996
rect 18328 6944 18380 6996
rect 20904 6944 20956 6996
rect 8208 6876 8260 6928
rect 10600 6876 10652 6928
rect 2688 6672 2740 6724
rect 3148 6672 3200 6724
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8392 6808 8444 6860
rect 10416 6808 10468 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 12716 6876 12768 6928
rect 4344 6740 4396 6792
rect 5080 6740 5132 6792
rect 6828 6740 6880 6792
rect 10508 6740 10560 6792
rect 13084 6740 13136 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 19524 6740 19576 6792
rect 19708 6783 19760 6792
rect 19708 6749 19742 6783
rect 19742 6749 19760 6783
rect 19708 6740 19760 6749
rect 23480 6808 23532 6860
rect 26056 6944 26108 6996
rect 27160 6944 27212 6996
rect 29368 6944 29420 6996
rect 21548 6740 21600 6792
rect 21916 6740 21968 6792
rect 27988 6808 28040 6860
rect 10784 6672 10836 6724
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 13360 6672 13412 6724
rect 20720 6672 20772 6724
rect 24676 6740 24728 6792
rect 25136 6740 25188 6792
rect 29184 6783 29236 6792
rect 29184 6749 29193 6783
rect 29193 6749 29227 6783
rect 29227 6749 29236 6783
rect 29184 6740 29236 6749
rect 12992 6604 13044 6656
rect 15844 6604 15896 6656
rect 16304 6604 16356 6656
rect 18788 6604 18840 6656
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 21272 6604 21324 6613
rect 23572 6647 23624 6656
rect 23572 6613 23581 6647
rect 23581 6613 23615 6647
rect 23615 6613 23624 6647
rect 23572 6604 23624 6613
rect 25872 6604 25924 6656
rect 30196 6783 30248 6792
rect 30196 6749 30205 6783
rect 30205 6749 30239 6783
rect 30239 6749 30248 6783
rect 30196 6740 30248 6749
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 7288 6400 7340 6452
rect 12900 6443 12952 6452
rect 12900 6409 12909 6443
rect 12909 6409 12943 6443
rect 12943 6409 12952 6443
rect 12900 6400 12952 6409
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 16488 6400 16540 6452
rect 20720 6400 20772 6452
rect 30012 6443 30064 6452
rect 30012 6409 30021 6443
rect 30021 6409 30055 6443
rect 30055 6409 30064 6443
rect 30012 6400 30064 6409
rect 2688 6332 2740 6384
rect 3884 6332 3936 6384
rect 7012 6332 7064 6384
rect 16028 6332 16080 6384
rect 21272 6332 21324 6384
rect 23572 6332 23624 6384
rect 28908 6375 28960 6384
rect 28908 6341 28942 6375
rect 28942 6341 28960 6375
rect 28908 6332 28960 6341
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 28356 6264 28408 6316
rect 5816 6196 5868 6248
rect 12348 6196 12400 6248
rect 14924 6239 14976 6248
rect 14924 6205 14933 6239
rect 14933 6205 14967 6239
rect 14967 6205 14976 6239
rect 14924 6196 14976 6205
rect 19524 6239 19576 6248
rect 19524 6205 19533 6239
rect 19533 6205 19567 6239
rect 19567 6205 19576 6239
rect 19524 6196 19576 6205
rect 3976 6060 4028 6112
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 23480 6128 23532 6180
rect 18420 6060 18472 6112
rect 24676 6060 24728 6112
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 13360 5856 13412 5908
rect 20168 5856 20220 5908
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 16580 5788 16632 5840
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 12716 5720 12768 5772
rect 6644 5652 6696 5704
rect 12348 5652 12400 5704
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 14924 5652 14976 5704
rect 24676 5652 24728 5704
rect 25596 5652 25648 5704
rect 4712 5584 4764 5636
rect 15936 5584 15988 5636
rect 14280 5516 14332 5568
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 10416 5312 10468 5364
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 14924 5312 14976 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 29736 5355 29788 5364
rect 29736 5321 29745 5355
rect 29745 5321 29779 5355
rect 29779 5321 29788 5355
rect 29736 5312 29788 5321
rect 2964 5244 3016 5296
rect 4068 5244 4120 5296
rect 3148 5176 3200 5228
rect 4712 5244 4764 5296
rect 9312 5244 9364 5296
rect 15844 5244 15896 5296
rect 18236 5287 18288 5296
rect 18236 5253 18245 5287
rect 18245 5253 18279 5287
rect 18279 5253 18288 5287
rect 18236 5244 18288 5253
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 28724 5244 28776 5296
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 11060 5176 11112 5228
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 6644 5108 6696 5160
rect 13268 5108 13320 5160
rect 25044 5108 25096 5160
rect 26700 5108 26752 5160
rect 29184 5176 29236 5228
rect 29920 5176 29972 5228
rect 13268 4972 13320 5024
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 25688 4972 25740 5024
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 5080 4632 5132 4684
rect 11704 4768 11756 4820
rect 13268 4768 13320 4820
rect 22468 4768 22520 4820
rect 14372 4700 14424 4752
rect 20996 4700 21048 4752
rect 24676 4743 24728 4752
rect 24676 4709 24685 4743
rect 24685 4709 24719 4743
rect 24719 4709 24728 4743
rect 24676 4700 24728 4709
rect 8944 4632 8996 4684
rect 7472 4607 7524 4616
rect 7472 4573 7506 4607
rect 7506 4573 7524 4607
rect 7472 4564 7524 4573
rect 10508 4564 10560 4616
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 17592 4632 17644 4684
rect 21180 4632 21232 4684
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 11980 4607 12032 4616
rect 11980 4573 12014 4607
rect 12014 4573 12032 4607
rect 11980 4564 12032 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 17040 4564 17092 4616
rect 18328 4564 18380 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20904 4564 20956 4616
rect 24400 4564 24452 4616
rect 25964 4564 26016 4616
rect 27160 4564 27212 4616
rect 13176 4496 13228 4548
rect 26608 4496 26660 4548
rect 9772 4428 9824 4480
rect 11060 4428 11112 4480
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16304 4428 16356 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 18236 4428 18288 4480
rect 19064 4428 19116 4480
rect 19708 4428 19760 4480
rect 20628 4428 20680 4480
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 22100 4428 22152 4480
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 26792 4428 26844 4480
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 8116 4224 8168 4276
rect 7472 4156 7524 4208
rect 7932 4156 7984 4208
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 10416 4224 10468 4276
rect 26608 4224 26660 4276
rect 8944 4088 8996 4140
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 9680 4020 9732 4072
rect 9956 4020 10008 4072
rect 11060 4088 11112 4140
rect 12348 4088 12400 4140
rect 14004 4088 14056 4140
rect 15292 4156 15344 4208
rect 18236 4156 18288 4208
rect 24400 4156 24452 4208
rect 25964 4156 26016 4208
rect 15568 4088 15620 4140
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17500 4088 17552 4140
rect 20720 4088 20772 4140
rect 21548 4088 21600 4140
rect 22100 4088 22152 4140
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 22284 4088 22336 4097
rect 14188 4020 14240 4072
rect 14556 4020 14608 4072
rect 24584 4131 24636 4140
rect 24584 4097 24618 4131
rect 24618 4097 24636 4131
rect 24584 4088 24636 4097
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 27436 4131 27488 4140
rect 27436 4097 27470 4131
rect 27470 4097 27488 4131
rect 27436 4088 27488 4097
rect 26700 4020 26752 4072
rect 14372 3952 14424 4004
rect 12716 3884 12768 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16672 3884 16724 3936
rect 19064 3927 19116 3936
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 21088 3884 21140 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 26608 3884 26660 3936
rect 28356 3884 28408 3936
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 20628 3680 20680 3732
rect 22376 3680 22428 3732
rect 24676 3680 24728 3732
rect 25044 3680 25096 3732
rect 9956 3544 10008 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 25964 3587 26016 3596
rect 25964 3553 25973 3587
rect 25973 3553 26007 3587
rect 26007 3553 26016 3587
rect 25964 3544 26016 3553
rect 26792 3723 26844 3732
rect 26792 3689 26801 3723
rect 26801 3689 26835 3723
rect 26835 3689 26844 3723
rect 26792 3680 26844 3689
rect 26240 3612 26292 3664
rect 28356 3612 28408 3664
rect 8208 3476 8260 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 12992 3476 13044 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19708 3519 19760 3528
rect 19708 3485 19742 3519
rect 19742 3485 19760 3519
rect 19708 3476 19760 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 23388 3476 23440 3528
rect 25688 3519 25740 3528
rect 25688 3485 25706 3519
rect 25706 3485 25740 3519
rect 25688 3476 25740 3485
rect 26608 3476 26660 3528
rect 14740 3408 14792 3460
rect 16948 3451 17000 3460
rect 16948 3417 16982 3451
rect 16982 3417 17000 3451
rect 16948 3408 17000 3417
rect 14004 3340 14056 3392
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 16856 3340 16908 3392
rect 18236 3340 18288 3392
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 12348 3136 12400 3188
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 15660 3136 15712 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 18236 3136 18288 3188
rect 19432 3136 19484 3188
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 27436 3136 27488 3188
rect 29920 3179 29972 3188
rect 29920 3145 29929 3179
rect 29929 3145 29963 3179
rect 29963 3145 29972 3179
rect 29920 3136 29972 3145
rect 9956 3000 10008 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 26700 3068 26752 3120
rect 28816 3068 28868 3120
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15476 2932 15528 2984
rect 10968 2864 11020 2916
rect 20812 3000 20864 3052
rect 20996 3000 21048 3052
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 22744 3000 22796 3052
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 25044 2932 25096 2984
rect 25780 2796 25832 2848
rect 26792 2864 26844 2916
rect 26240 2796 26292 2848
rect 26608 2796 26660 2848
rect 27160 2796 27212 2848
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 14372 2592 14424 2644
rect 10140 2524 10192 2576
rect 10968 2524 11020 2576
rect 18236 2456 18288 2508
rect 1216 2320 1268 2372
rect 2504 2320 2556 2372
rect 4160 2363 4212 2372
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 4160 2320 4212 2329
rect 5080 2320 5132 2372
rect 6368 2388 6420 2440
rect 7656 2388 7708 2440
rect 8944 2388 8996 2440
rect 10232 2388 10284 2440
rect 11520 2388 11572 2440
rect 12808 2388 12860 2440
rect 14004 2388 14056 2440
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16304 2388 16356 2440
rect 19064 2388 19116 2440
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 21088 2388 21140 2440
rect 23388 2388 23440 2440
rect 25044 2431 25096 2440
rect 25044 2397 25053 2431
rect 25053 2397 25087 2431
rect 25087 2397 25096 2431
rect 25044 2388 25096 2397
rect 26240 2431 26292 2440
rect 26240 2397 26249 2431
rect 26249 2397 26283 2431
rect 26283 2397 26292 2431
rect 26240 2388 26292 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 29552 2388 29604 2440
rect 30840 2388 30892 2440
rect 32128 2388 32180 2440
rect 33416 2388 33468 2440
rect 13176 2320 13228 2372
rect 14096 2320 14148 2372
rect 15384 2320 15436 2372
rect 16672 2320 16724 2372
rect 18236 2320 18288 2372
rect 19340 2320 19392 2372
rect 20720 2320 20772 2372
rect 22100 2320 22152 2372
rect 23480 2363 23532 2372
rect 23480 2329 23489 2363
rect 23489 2329 23523 2363
rect 23523 2329 23532 2363
rect 23480 2320 23532 2329
rect 24400 2320 24452 2372
rect 25688 2320 25740 2372
rect 26976 2320 27028 2372
rect 28264 2320 28316 2372
rect 8116 2252 8168 2304
rect 34612 2252 34664 2304
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
<< metal2 >>
rect 1766 35200 1822 36000
rect 4710 35306 4766 36000
rect 7654 35306 7710 36000
rect 4710 35278 4936 35306
rect 4710 35200 4766 35278
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14074 1716 14894
rect 1780 14482 1808 35200
rect 4908 33590 4936 35278
rect 7654 35278 7880 35306
rect 7654 35200 7710 35278
rect 7852 33590 7880 35278
rect 10598 35200 10654 36000
rect 13542 35306 13598 36000
rect 16486 35306 16542 36000
rect 13542 35278 13860 35306
rect 13542 35200 13598 35278
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 10612 33590 10640 35200
rect 13832 33590 13860 35278
rect 16486 35278 16620 35306
rect 16486 35200 16542 35278
rect 16592 33590 16620 35278
rect 19430 35200 19486 36000
rect 22374 35200 22430 36000
rect 25318 35306 25374 36000
rect 28262 35306 28318 36000
rect 31206 35306 31262 36000
rect 34150 35306 34206 36000
rect 25318 35278 25636 35306
rect 25318 35200 25374 35278
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 19444 33590 19472 35200
rect 22388 33590 22416 35200
rect 25608 33590 25636 35278
rect 28262 35278 28580 35306
rect 28262 35200 28318 35278
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 28552 33590 28580 35278
rect 31206 35278 31524 35306
rect 31206 35200 31262 35278
rect 31496 33590 31524 35278
rect 34150 35278 34284 35306
rect 34150 35200 34206 35278
rect 34256 33590 34284 35278
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 4896 33584 4948 33590
rect 4896 33526 4948 33532
rect 7840 33584 7892 33590
rect 7840 33526 7892 33532
rect 10600 33584 10652 33590
rect 10600 33526 10652 33532
rect 13820 33584 13872 33590
rect 13820 33526 13872 33532
rect 16580 33584 16632 33590
rect 16580 33526 16632 33532
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 31484 33584 31536 33590
rect 31484 33526 31536 33532
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 22468 33380 22520 33386
rect 22468 33322 22520 33328
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 28356 33380 28408 33386
rect 28356 33322 28408 33328
rect 31300 33380 31352 33386
rect 31300 33322 31352 33328
rect 33324 33380 33376 33386
rect 33324 33322 33376 33328
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 11612 33312 11664 33318
rect 11612 33254 11664 33260
rect 3332 25288 3384 25294
rect 3332 25230 3384 25236
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2792 24410 2820 24686
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2884 24290 2912 25094
rect 2792 24274 2912 24290
rect 2780 24268 2912 24274
rect 2832 24262 2912 24268
rect 2780 24210 2832 24216
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2332 23866 2360 24074
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2884 23322 2912 24262
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2976 21486 3004 24210
rect 3344 23594 3372 25230
rect 3976 25220 4028 25226
rect 3976 25162 4028 25168
rect 3988 24818 4016 25162
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3436 23322 3464 24074
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3988 23186 4016 24754
rect 4080 24614 4108 25230
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3160 22098 3188 23054
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3988 21554 4016 22918
rect 4264 22642 4292 24006
rect 4356 23594 4384 24550
rect 4724 23798 4752 24686
rect 4816 23798 4844 25230
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4804 23792 4856 23798
rect 4804 23734 4856 23740
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4356 23050 4384 23530
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4344 23044 4396 23050
rect 4344 22986 4396 22992
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4356 22438 4384 22986
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4448 22094 4476 23258
rect 4540 22506 4568 23666
rect 4724 22982 4752 23734
rect 4816 23322 4844 23734
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4908 23254 4936 23462
rect 4896 23248 4948 23254
rect 4896 23190 4948 23196
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4528 22500 4580 22506
rect 4528 22442 4580 22448
rect 4540 22386 4568 22442
rect 4540 22358 4752 22386
rect 4448 22066 4660 22094
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3068 20534 3096 21286
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 3160 20466 3188 20742
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2424 19922 2452 20266
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1872 19514 1900 19790
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 2976 19446 3004 20198
rect 3252 19922 3280 20878
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 17134 2728 17546
rect 2976 17270 3004 18838
rect 3344 18766 3372 19722
rect 3436 18766 3464 20470
rect 3528 19854 3556 20878
rect 3620 20534 3648 21286
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 20058 4016 20402
rect 4080 20398 4108 21354
rect 4540 21010 4568 21490
rect 4528 21004 4580 21010
rect 4528 20946 4580 20952
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4540 19854 4568 20946
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3252 17678 3280 18634
rect 3528 17814 3556 19314
rect 4264 19242 4292 19722
rect 4632 19378 4660 22066
rect 4724 19718 4752 22358
rect 4908 19786 4936 23190
rect 5000 22234 5028 33254
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 8588 31822 8616 32234
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8576 31816 8628 31822
rect 8576 31758 8628 31764
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 8772 28014 8800 31894
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 9876 31482 9904 31826
rect 10060 31686 10088 32166
rect 10152 31822 10180 32710
rect 10520 32434 10548 32846
rect 10416 32428 10468 32434
rect 10416 32370 10468 32376
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10048 31680 10100 31686
rect 10048 31622 10100 31628
rect 10060 31498 10088 31622
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9968 31470 10088 31498
rect 9968 31346 9996 31470
rect 10048 31408 10100 31414
rect 10048 31350 10100 31356
rect 8852 31340 8904 31346
rect 8852 31282 8904 31288
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 8864 28150 8892 31282
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9416 30938 9444 31214
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9508 30734 9536 31214
rect 10060 30938 10088 31350
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10244 30938 10272 31282
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10428 30734 10456 32370
rect 10520 31822 10548 32370
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10520 30802 10548 31758
rect 10612 31414 10640 32166
rect 11624 31754 11652 33254
rect 12268 32570 12296 33322
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 13280 32502 13308 32710
rect 14292 32570 14320 33322
rect 16868 32978 16896 33322
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 15476 32836 15528 32842
rect 15476 32778 15528 32784
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 18328 32836 18380 32842
rect 18328 32778 18380 32784
rect 14280 32564 14332 32570
rect 14280 32506 14332 32512
rect 11796 32496 11848 32502
rect 11796 32438 11848 32444
rect 13268 32496 13320 32502
rect 13268 32438 13320 32444
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 11612 31748 11664 31754
rect 11612 31690 11664 31696
rect 10600 31408 10652 31414
rect 10600 31350 10652 31356
rect 10692 31204 10744 31210
rect 10692 31146 10744 31152
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 9036 29776 9088 29782
rect 9036 29718 9088 29724
rect 9048 29170 9076 29718
rect 9968 29510 9996 30670
rect 10152 29578 10180 30670
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10428 29510 10456 29582
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 9324 29170 9352 29446
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 8944 28960 8996 28966
rect 8944 28902 8996 28908
rect 8956 28218 8984 28902
rect 9048 28490 9076 29106
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 9324 28422 9352 29106
rect 9508 28626 9536 29106
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 8944 28212 8996 28218
rect 8944 28154 8996 28160
rect 8852 28144 8904 28150
rect 8852 28086 8904 28092
rect 8864 28014 8892 28086
rect 8956 28014 8984 28154
rect 9140 28082 9168 28358
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 8220 26994 8248 27338
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8772 26790 8800 27950
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9036 27532 9088 27538
rect 9036 27474 9088 27480
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 9048 26314 9076 27474
rect 9140 27470 9168 27814
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9140 26926 9168 26998
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9036 26308 9088 26314
rect 9036 26250 9088 26256
rect 9232 26042 9260 26726
rect 9324 26518 9352 27814
rect 9600 27470 9628 27814
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 9784 26994 9812 27814
rect 10612 27062 10640 30670
rect 10704 29714 10732 31146
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10704 29578 10732 29650
rect 10692 29572 10744 29578
rect 10692 29514 10744 29520
rect 10704 28558 10732 29514
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10704 28082 10732 28494
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 11164 26450 11192 26726
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9232 25838 9260 25978
rect 9324 25906 9352 26182
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 10704 25294 10732 25842
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 5092 24274 5120 24822
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 5080 24268 5132 24274
rect 5080 24210 5132 24216
rect 5552 24206 5580 25094
rect 6840 24818 6868 25230
rect 7484 24818 7512 25230
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 6736 24676 6788 24682
rect 6736 24618 6788 24624
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5828 23798 5856 24006
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 6748 23662 6776 24618
rect 6840 24410 6868 24754
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5092 19786 5120 20402
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16794 2728 17070
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2608 15502 2636 16594
rect 3068 16522 3096 17478
rect 3160 16776 3188 17478
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4264 16794 4292 17138
rect 3240 16788 3292 16794
rect 3160 16748 3240 16776
rect 3240 16730 3292 16736
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2608 13462 2636 15438
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2976 15094 3004 15370
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14414 2728 14894
rect 3068 14414 3096 16458
rect 3252 14890 3280 16730
rect 5000 15706 5028 19654
rect 5092 19514 5120 19722
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 6748 19378 6776 23598
rect 7024 22642 7052 24142
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7116 23322 7144 23598
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7208 23118 7236 23666
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7116 22710 7144 23054
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7208 22522 7236 23054
rect 7116 22494 7236 22522
rect 7116 22030 7144 22494
rect 7300 22094 7328 24210
rect 7484 23526 7512 24754
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7852 23594 7880 24074
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7484 22642 7512 23462
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7576 22778 7604 23054
rect 7852 22982 7880 23530
rect 8220 22982 8248 24142
rect 8404 23798 8432 24686
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 8392 23792 8444 23798
rect 8392 23734 8444 23740
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8312 23186 8340 23598
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7208 22066 7328 22094
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7208 21894 7236 22066
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19990 6960 20198
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5092 15502 5120 16458
rect 6380 16454 6408 17614
rect 6472 17066 6500 18294
rect 6656 18290 6684 19314
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6656 17202 6684 18226
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6748 17882 6776 18158
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6932 17338 6960 18158
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6472 16726 6500 17002
rect 6656 16794 6684 17138
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 13938 3096 14350
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12782 2452 13126
rect 2608 12986 2636 13398
rect 2976 13326 3004 13670
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 3068 12442 3096 12854
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3252 12238 3280 13126
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10266 2820 10610
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2792 9602 2820 10202
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2976 9722 3004 10134
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2700 9574 2820 9602
rect 2700 9450 2728 9574
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2792 9178 2820 9454
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 8906 2912 9318
rect 2976 9178 3004 9658
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3068 7886 3096 12174
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 9994 3188 10542
rect 3252 10538 3280 12174
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3344 10062 3372 10678
rect 3804 10674 3832 14214
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 12986 3924 13262
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12986 4016 13194
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4080 12850 4108 13874
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4264 13734 4292 14758
rect 4448 14006 4476 15302
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12434 4108 12786
rect 3988 12406 4108 12434
rect 3988 11082 4016 12406
rect 4264 11082 4292 13670
rect 4540 12850 4568 14962
rect 5092 13870 5120 15438
rect 5552 15434 5580 15914
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5736 15162 5764 16118
rect 6472 16114 6500 16662
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16114 6592 16458
rect 6656 16114 6684 16526
rect 6748 16250 6776 17138
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6564 15502 6592 16050
rect 6656 15570 6684 16050
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6748 15502 6776 16186
rect 6840 16182 6868 17138
rect 7024 17134 7052 19246
rect 7116 18834 7144 19926
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7208 18698 7236 21830
rect 7484 21010 7512 21966
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7300 20466 7328 20878
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19786 7328 20402
rect 7392 19854 7420 20742
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7300 18154 7328 19722
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7116 16658 7144 17614
rect 7484 17202 7512 20946
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20058 7696 20878
rect 7852 20602 7880 22714
rect 8404 22710 8432 23734
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 8496 22506 8524 23122
rect 8680 23050 8708 23190
rect 9324 23118 9352 24142
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9600 23338 9628 23598
rect 9600 23310 9904 23338
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 8668 23044 8720 23050
rect 8668 22986 8720 22992
rect 9324 22710 9352 23054
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 9784 22710 9812 22986
rect 9312 22704 9364 22710
rect 9312 22646 9364 22652
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8496 21894 8524 22442
rect 9220 22432 9272 22438
rect 9220 22374 9272 22380
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7760 19990 7788 20470
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18970 7696 19314
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16454 7144 16594
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 7116 16046 7144 16390
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7668 15570 7696 16390
rect 7760 15706 7788 17138
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 5736 14346 5764 15098
rect 5828 15094 5856 15438
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 6104 14550 6132 15302
rect 6564 14822 6592 15438
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6840 14618 6868 15302
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6104 14414 6132 14486
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 13938 5856 14214
rect 6472 14006 6500 14282
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13326 5120 13806
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 5552 13530 5580 13874
rect 6840 13734 6868 14554
rect 7484 14346 7512 15438
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5264 13388 5316 13394
rect 5644 13376 5672 13466
rect 5316 13348 5672 13376
rect 5264 13330 5316 13336
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4540 11354 4568 12786
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3436 9602 3464 10542
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3160 9586 3464 9602
rect 3148 9580 3464 9586
rect 3200 9574 3464 9580
rect 3148 9522 3200 9528
rect 3436 9518 3464 9574
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3252 8498 3280 9386
rect 3528 8634 3556 9522
rect 3620 8974 3648 10406
rect 3804 9926 3832 10610
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3988 9738 4016 11018
rect 4264 10674 4292 11018
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4264 10130 4292 10474
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3896 9710 4016 9738
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 7002 2544 7346
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 7002 2636 7142
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 3068 6746 3096 7822
rect 3620 7818 3648 8910
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3896 7410 3924 9710
rect 4080 9450 4108 9930
rect 4264 9586 4292 10066
rect 4356 10062 4384 10950
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9722 4384 9998
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3988 8498 4016 8978
rect 4080 8634 4108 9386
rect 4356 8974 4384 9658
rect 4540 9586 4568 10202
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 5092 9450 5120 11086
rect 5828 11082 5856 12718
rect 6932 12434 6960 14214
rect 7116 14006 7144 14282
rect 7852 14278 7880 20198
rect 8036 19854 8064 20402
rect 8404 19854 8432 20402
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 18902 8432 19790
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16794 8248 16934
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 15910 8340 16662
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8116 14408 8168 14414
rect 8168 14368 8248 14396
rect 8116 14350 8168 14356
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7944 14074 7972 14282
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 6932 12406 7052 12434
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 5828 9994 5856 11018
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10606 6684 10746
rect 6932 10742 6960 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3068 6730 3188 6746
rect 2688 6724 2740 6730
rect 3068 6724 3200 6730
rect 3068 6718 3148 6724
rect 2688 6666 2740 6672
rect 3148 6666 3200 6672
rect 2700 6390 2728 6666
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 3160 6322 3188 6666
rect 3896 6390 3924 7346
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2976 5302 3004 6258
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 3160 5234 3188 6258
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5302 4108 7754
rect 4356 6798 4384 8774
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 5828 7478 5856 9930
rect 5920 9654 5948 9998
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5302 4752 5578
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 5092 4690 5120 6734
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 5828 5778 5856 6190
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5234 5856 5714
rect 6656 5710 6684 10542
rect 6748 10266 6776 10678
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 6798 6868 7414
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 7024 6390 7052 12406
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10130 7236 11086
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10742 7328 10950
rect 7576 10742 7604 12582
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9586 7512 9930
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7478 7420 7754
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6458 7328 6598
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 6656 5166 6684 5646
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 7484 4622 7512 9522
rect 7852 6866 7880 10950
rect 8220 10810 8248 14368
rect 8312 13938 8340 15846
rect 8496 15162 8524 21830
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 19786 9076 20334
rect 9232 19990 9260 22374
rect 9324 22030 9352 22646
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 9876 21690 9904 23310
rect 10060 22778 10088 23666
rect 10520 23662 10548 24006
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10244 22438 10272 22918
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 9048 19378 9076 19722
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18290 8616 19110
rect 9048 18426 9076 19314
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18834 9168 19110
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 9232 17270 9260 19926
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 9784 19378 9812 19722
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 9784 18290 9812 18634
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9784 16998 9812 18226
rect 9876 17202 9904 21626
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20466 10272 20742
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10244 19786 10272 20402
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10336 19378 10364 23258
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10428 22642 10456 22918
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10428 20942 10456 22374
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10428 20398 10456 20878
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 19854 10456 20334
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18766 10180 19110
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10336 18170 10364 19314
rect 10152 18142 10364 18170
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9876 16946 9904 17138
rect 10048 16992 10100 16998
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16454 9720 16526
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 13326 8340 13874
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4214 7512 4558
rect 8128 4282 8156 10406
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 7954 8340 8230
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 6934 8248 7822
rect 8404 7342 8432 13806
rect 8496 13394 8524 14486
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 13802 8616 14282
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8588 12918 8616 13194
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8864 12782 8892 14486
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8956 10810 8984 13126
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8864 9722 8892 10678
rect 9048 9994 9076 13330
rect 9140 13326 9168 14554
rect 9324 14550 9352 16050
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 13938 9260 14350
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9140 12986 9168 13262
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10674 9260 10950
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9140 10266 9168 10610
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 9324 8566 9352 14486
rect 9784 14362 9812 16934
rect 9876 16918 9996 16946
rect 10048 16934 10100 16940
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 16658 9904 16730
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9968 15162 9996 16918
rect 10060 16590 10088 16934
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10152 16454 10180 18142
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9968 15026 9996 15098
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9508 14346 9812 14362
rect 9496 14340 9812 14346
rect 9548 14334 9812 14340
rect 9496 14282 9548 14288
rect 10244 14278 10272 18022
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10336 15026 10364 17206
rect 10428 17066 10456 19790
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16658 10456 17002
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 15502 10456 16390
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10520 15026 10548 23598
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 20942 10732 21830
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10704 19786 10732 20878
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 18766 10640 19110
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10612 15570 10640 17070
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10612 14906 10640 15506
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10336 14878 10640 14906
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 13258 9904 13806
rect 10336 13802 10364 14878
rect 10704 14346 10732 14962
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 10336 10810 10364 13738
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 10588 9536 10678
rect 9864 10600 9916 10606
rect 9508 10560 9864 10588
rect 9864 10542 9916 10548
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7886 9904 8230
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 7944 3738 7972 4150
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 1228 800 1256 2314
rect 2516 800 2544 2314
rect 3804 870 3924 898
rect 3804 800 3832 870
rect 1214 0 1270 800
rect 2502 0 2558 800
rect 3790 0 3846 800
rect 3896 762 3924 870
rect 4172 762 4200 2314
rect 5092 800 5120 2314
rect 6380 800 6408 2382
rect 7668 800 7696 2382
rect 8128 2310 8156 4218
rect 8220 3534 8248 6870
rect 8404 6866 8432 7142
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8956 4690 8984 7278
rect 9876 6914 9904 7822
rect 9876 6886 9996 6914
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4146 8984 4626
rect 9324 4282 9352 5238
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9692 4078 9720 4218
rect 9784 4146 9812 4422
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9968 4078 9996 6886
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3602 9996 4014
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 9968 3058 9996 3538
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10152 2582 10180 10406
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10244 7478 10272 7754
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10612 6934 10640 7822
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 5370 10456 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 5370 10548 6734
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10428 4282 10456 5170
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10520 4146 10548 4558
rect 10612 4146 10640 6870
rect 10704 6866 10732 14282
rect 10888 13530 10916 22918
rect 11532 22234 11560 22986
rect 11716 22642 11744 31894
rect 11808 31754 11836 32438
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13360 32224 13412 32230
rect 13360 32166 13412 32172
rect 11900 31754 11928 32166
rect 11796 31748 11848 31754
rect 11900 31726 12020 31754
rect 11796 31690 11848 31696
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11900 28626 11928 29106
rect 11888 28620 11940 28626
rect 11888 28562 11940 28568
rect 11992 24206 12020 31726
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12452 29102 12480 31214
rect 12728 29510 12756 31282
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29646 12940 29990
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12728 29170 12756 29446
rect 12820 29170 12848 29446
rect 12912 29306 12940 29582
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12452 28558 12480 28630
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12360 28082 12388 28358
rect 12544 28082 12572 28562
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12636 28150 12664 28426
rect 12624 28144 12676 28150
rect 12624 28086 12676 28092
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12084 26994 12112 27066
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12084 25974 12112 26930
rect 12360 26042 12388 27338
rect 12452 26994 12480 27950
rect 12544 27538 12572 28018
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12728 27402 12756 29106
rect 12820 28694 12848 29106
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12728 27062 12756 27338
rect 12912 27130 12940 28358
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26738 12480 26930
rect 12624 26784 12676 26790
rect 12452 26710 12572 26738
rect 12624 26726 12676 26732
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12452 26042 12480 26522
rect 12544 26314 12572 26710
rect 12636 26382 12664 26726
rect 12912 26586 12940 27066
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 12360 25906 12388 25978
rect 12544 25974 12572 26250
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12728 25294 12756 25638
rect 13096 25362 13124 25638
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11992 23322 12020 24142
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22234 11744 22578
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11072 20466 11100 22034
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11532 19310 11560 19654
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11072 18290 11100 19246
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11624 17746 11652 22034
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21622 11744 21898
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11808 21554 11836 22510
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11992 21570 12020 22442
rect 12084 22098 12112 23054
rect 12452 22642 12480 24142
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12636 22642 12664 24006
rect 12912 23730 12940 24006
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13188 23662 13216 32166
rect 13372 31890 13400 32166
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 14292 31482 14320 31758
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13280 30938 13308 31214
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 14108 30734 14136 31282
rect 14660 31278 14688 31758
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14292 30258 14320 31078
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13372 28626 13400 29106
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 13280 28082 13308 28494
rect 13372 28218 13400 28562
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 14200 28082 14228 29514
rect 14568 29306 14596 30670
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 14660 29186 14688 31214
rect 14844 30870 14872 31282
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14844 29850 14872 30806
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 14936 30258 14964 30670
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14936 29306 14964 30194
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14924 29300 14976 29306
rect 14924 29242 14976 29248
rect 14568 29158 14688 29186
rect 14568 28558 14596 29158
rect 15028 29102 15056 29582
rect 15108 29572 15160 29578
rect 15108 29514 15160 29520
rect 15120 29238 15148 29514
rect 15108 29232 15160 29238
rect 15108 29174 15160 29180
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15028 28626 15056 29038
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 14016 27538 14044 28018
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14200 27470 14228 28018
rect 14568 28014 14596 28494
rect 15028 28150 15056 28562
rect 15120 28558 15148 29174
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15396 28218 15424 28494
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15016 28144 15068 28150
rect 15016 28086 15068 28092
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14200 27062 14228 27406
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 13360 26580 13412 26586
rect 13360 26522 13412 26528
rect 13372 25974 13400 26522
rect 13464 26466 13492 26998
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 13464 26438 13584 26466
rect 13556 26314 13584 26438
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13464 25906 13492 26250
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13464 24274 13492 25094
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13280 23730 13308 24142
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12452 22166 12480 22578
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12912 22030 12940 22442
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22030 13032 22374
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 11992 21554 12112 21570
rect 11796 21548 11848 21554
rect 11992 21548 12124 21554
rect 11992 21542 12072 21548
rect 11796 21490 11848 21496
rect 12072 21490 12124 21496
rect 11808 18290 11836 21490
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11900 19922 11928 20946
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12084 18698 12112 21490
rect 12912 21146 12940 21966
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 18766 12480 19382
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12084 18358 12112 18634
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 16794 11008 17478
rect 11624 17134 11652 17682
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10980 15502 11008 16730
rect 11164 16522 11192 16934
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 15502 11192 16458
rect 11624 15706 11652 17070
rect 12084 16726 12112 18294
rect 12348 18284 12400 18290
rect 12400 18244 12480 18272
rect 12348 18226 12400 18232
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12176 17610 12204 18158
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 16794 12296 17206
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12452 16658 12480 18244
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11992 14006 12020 14758
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10888 12714 10916 13466
rect 11808 13326 11836 13806
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12918 11836 13262
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 11992 11150 12020 13942
rect 12084 13258 12112 14894
rect 12452 14346 12480 16594
rect 12728 16250 12756 19314
rect 12820 17610 12848 20266
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 13004 17542 13032 18226
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 14074 12480 14282
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11072 10130 11100 11086
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 11164 8906 11192 11018
rect 12084 10062 12112 13194
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12360 10606 12388 11154
rect 12544 11150 12572 15302
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12452 10674 12480 11018
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9654 12112 9998
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11164 7478 11192 8842
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10796 6730 10824 7142
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 4486 11100 5170
rect 11716 4826 11744 7278
rect 12084 6914 12112 9590
rect 12544 9178 12572 10678
rect 12636 10266 12664 11018
rect 12728 10810 12756 15030
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 14074 12848 14350
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13004 12918 13032 17478
rect 13188 17270 13216 23598
rect 13280 22930 13308 23666
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 13280 22902 13492 22930
rect 13464 22642 13492 22902
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13464 22094 13492 22578
rect 14200 22574 14228 23530
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 13372 22066 13492 22094
rect 13372 20398 13400 22066
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 19854 13400 20334
rect 13464 19854 13492 20878
rect 14200 20602 14228 22510
rect 14476 20942 14504 25706
rect 14568 24206 14596 27950
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14660 23662 14688 25774
rect 14752 24818 14780 26386
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14660 23118 14688 23598
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22642 14688 22918
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14200 20398 14228 20538
rect 14384 20534 14412 20742
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 14188 20392 14240 20398
rect 14844 20369 14872 24142
rect 14936 23866 14964 24550
rect 15028 24274 15056 28086
rect 15488 26874 15516 32778
rect 16776 32570 16804 32778
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15948 32026 15976 32370
rect 15844 32020 15896 32026
rect 15844 31962 15896 31968
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15660 31952 15712 31958
rect 15660 31894 15712 31900
rect 15672 31414 15700 31894
rect 15856 31754 15884 31962
rect 15856 31748 15988 31754
rect 15856 31726 15936 31748
rect 15752 31680 15804 31686
rect 15752 31622 15804 31628
rect 15660 31408 15712 31414
rect 15660 31350 15712 31356
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15580 30734 15608 31282
rect 15764 31278 15792 31622
rect 15856 31482 15884 31726
rect 15936 31690 15988 31696
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 15844 31476 15896 31482
rect 15844 31418 15896 31424
rect 16684 31414 16712 31622
rect 16028 31408 16080 31414
rect 16028 31350 16080 31356
rect 16672 31408 16724 31414
rect 16672 31350 16724 31356
rect 15752 31272 15804 31278
rect 15752 31214 15804 31220
rect 15764 30802 15792 31214
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 16040 30734 16068 31350
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 16040 30326 16068 30670
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 15580 28150 15608 29106
rect 16408 28558 16436 29106
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 16396 28552 16448 28558
rect 16396 28494 16448 28500
rect 15568 28144 15620 28150
rect 15568 28086 15620 28092
rect 15764 28082 15792 28494
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15488 26846 15608 26874
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24818 15240 25094
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14936 23186 14964 23802
rect 15028 23798 15056 24210
rect 15304 23866 15332 24754
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15212 23186 15240 23598
rect 15304 23186 15332 23802
rect 15396 23662 15424 25230
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15488 24070 15516 24686
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23730 15516 24006
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15488 23186 15516 23462
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15028 22710 15056 23054
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15304 22234 15332 22578
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15580 20534 15608 26846
rect 15672 26586 15700 26930
rect 15660 26580 15712 26586
rect 15660 26522 15712 26528
rect 15672 25498 15700 26522
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15764 25158 15792 28018
rect 15948 25294 15976 28426
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16040 27606 16068 28086
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16040 27470 16068 27542
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 16408 26994 16436 28494
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15672 22642 15700 24006
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15948 22574 15976 25230
rect 16316 24818 16344 25366
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16408 24206 16436 26930
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15856 20466 15884 21490
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 14924 20392 14976 20398
rect 14188 20334 14240 20340
rect 14830 20360 14886 20369
rect 14096 20324 14148 20330
rect 14924 20334 14976 20340
rect 14830 20295 14886 20304
rect 14096 20266 14148 20272
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 14108 19922 14136 20266
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13280 15638 13308 16050
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 14006 13124 14282
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12820 9450 12848 10950
rect 12912 10742 12940 11086
rect 13004 11014 13032 12650
rect 13096 11150 13124 13126
rect 13280 11150 13308 14826
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12912 7392 12940 10678
rect 12820 7364 12940 7392
rect 11992 6886 12112 6914
rect 12716 6928 12768 6934
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11716 4622 11744 4762
rect 11992 4622 12020 6886
rect 12820 6914 12848 7364
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12768 6886 12848 6914
rect 12716 6870 12768 6876
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5710 12388 6190
rect 12728 5778 12756 6870
rect 12912 6458 12940 7210
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6798 13124 7142
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6458 13032 6598
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4146 11100 4422
rect 12360 4146 12388 5646
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12728 3942 12756 5714
rect 13188 4554 13216 11018
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 5166 13308 10950
rect 13372 6730 13400 19790
rect 13464 15570 13492 19790
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 14752 18766 14780 19246
rect 14936 19174 14964 20334
rect 15672 20058 15700 20402
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14936 18970 14964 19110
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18358 14780 18702
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14384 16114 14412 16526
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 14384 15502 14412 16050
rect 14752 16046 14780 16594
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13938 13768 14350
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 11762 13492 13670
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 14108 13258 14136 13806
rect 14568 13462 14596 15438
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 14384 12238 14412 12582
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14568 11762 14596 13398
rect 14752 12918 14780 15982
rect 15120 15638 15148 19790
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15212 17678 15240 18566
rect 15396 17882 15424 18702
rect 15672 18290 15700 19722
rect 15856 19446 15884 20402
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 16040 19446 16068 19722
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15764 18426 15792 18634
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15856 18358 15884 19382
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15396 17202 15424 17818
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15212 16182 15240 16662
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15396 16454 15424 16526
rect 15948 16454 15976 17070
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15948 15978 15976 16390
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 15026 15700 15438
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15396 13394 15424 13874
rect 15672 13530 15700 14962
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15580 12850 15608 13194
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15212 12238 15240 12786
rect 15764 12238 15792 13262
rect 15948 13190 15976 13874
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12374 15976 13126
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 14752 11762 14780 12174
rect 15212 11830 15240 12174
rect 15764 11830 15792 12174
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15948 11762 15976 12310
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 13464 10742 13492 11698
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5914 13400 6054
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4826 13308 4966
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 14292 4622 14320 5510
rect 14384 4758 14412 5646
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3534 13032 3878
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12360 3194 12388 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10980 2582 11008 2858
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8956 800 8984 2382
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 10244 800 10272 2382
rect 11532 800 11560 2382
rect 12820 800 12848 2382
rect 13188 2378 13216 4490
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 14016 3398 14044 4082
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 14016 2446 14044 3334
rect 14200 2990 14228 4014
rect 14384 4010 14412 4422
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14476 3890 14504 10406
rect 16040 9450 16068 19382
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16224 18426 16252 18906
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 15502 16160 16390
rect 16224 16114 16252 17546
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 12782 16160 15438
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16224 9654 16252 16050
rect 16316 15366 16344 22578
rect 16500 21894 16528 23598
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16408 15570 16436 15982
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16500 15162 16528 21830
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16590 16620 17478
rect 16684 17202 16712 21286
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16592 14958 16620 16050
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12850 16436 13262
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16592 12170 16620 14894
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7410 15240 8230
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15304 6798 15332 8298
rect 15396 7546 15424 8842
rect 16040 8498 16068 9386
rect 16224 8498 16252 9590
rect 16684 8838 16712 11018
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15856 6746 15884 8298
rect 15856 6718 15976 6746
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14936 5710 14964 6190
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14936 5370 14964 5646
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15856 5302 15884 6598
rect 15948 5642 15976 6718
rect 16040 6390 16068 8298
rect 16224 7546 16252 8434
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16316 6662 16344 7754
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16500 6458 16528 8366
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16592 5846 16620 8570
rect 16684 8498 16712 8774
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16776 6914 16804 32506
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 16868 31210 16896 32370
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 17144 31346 17172 31826
rect 17880 31822 17908 32370
rect 18248 32026 18276 32370
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 17316 31816 17368 31822
rect 17868 31816 17920 31822
rect 17316 31758 17368 31764
rect 17696 31776 17868 31804
rect 17328 31482 17356 31758
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17696 31346 17724 31776
rect 17868 31758 17920 31764
rect 18340 31686 18368 32778
rect 19536 32230 19564 33322
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 20640 32026 20668 32914
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21284 32366 21312 32710
rect 22020 32434 22048 32710
rect 22480 32570 22508 33322
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22652 32428 22704 32434
rect 22652 32370 22704 32376
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21088 32292 21140 32298
rect 21088 32234 21140 32240
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 16856 31204 16908 31210
rect 16856 31146 16908 31152
rect 17604 30666 17632 31282
rect 17592 30660 17644 30666
rect 17592 30602 17644 30608
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 19616 29640 19668 29646
rect 19616 29582 19668 29588
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 19536 29170 19564 29446
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19524 29164 19576 29170
rect 19524 29106 19576 29112
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16868 26042 16896 26250
rect 17144 26042 17172 26522
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 17236 25906 17264 27474
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 18248 27130 18276 27406
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18248 26450 18276 27066
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17052 24954 17080 25842
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 17696 24818 17724 25842
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 18248 24818 18276 26250
rect 18340 25702 18368 26930
rect 18432 26790 18460 28426
rect 19352 28150 19380 29106
rect 19628 28558 19656 29582
rect 20180 29306 20208 30194
rect 20364 29646 20392 31282
rect 20548 31278 20576 31894
rect 21100 31890 21128 32234
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 22664 31958 22692 32370
rect 22848 32366 22876 32846
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 22652 31952 22704 31958
rect 22652 31894 22704 31900
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20824 31482 20852 31758
rect 21100 31754 21128 31826
rect 22848 31822 22876 32302
rect 23216 32026 23244 32370
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 22928 31884 22980 31890
rect 22928 31826 22980 31832
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21364 31816 21416 31822
rect 22836 31816 22888 31822
rect 21364 31758 21416 31764
rect 22664 31776 22836 31804
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20548 29714 20576 31214
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20996 30660 21048 30666
rect 20996 30602 21048 30608
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 20364 29152 20392 29582
rect 20548 29238 20576 29650
rect 20536 29232 20588 29238
rect 20536 29174 20588 29180
rect 20640 29170 20668 29990
rect 20824 29714 20852 30194
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20732 29170 20760 29582
rect 20444 29164 20496 29170
rect 20364 29124 20444 29152
rect 20444 29106 20496 29112
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20732 28966 20760 29106
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20732 28558 20760 28902
rect 20824 28626 20852 29650
rect 20916 29578 20944 30194
rect 20904 29572 20956 29578
rect 20904 29514 20956 29520
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20916 28558 20944 29514
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 19628 28218 19656 28494
rect 19904 28218 19932 28494
rect 19616 28212 19668 28218
rect 19616 28154 19668 28160
rect 19892 28212 19944 28218
rect 19892 28154 19944 28160
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 19352 26450 19380 28086
rect 19996 28014 20024 28494
rect 20916 28150 20944 28494
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 21008 27538 21036 30602
rect 21192 28762 21220 31758
rect 21376 31278 21404 31758
rect 22664 31346 22692 31776
rect 22836 31758 22888 31764
rect 22940 31346 22968 31826
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 21364 31272 21416 31278
rect 21364 31214 21416 31220
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21376 29306 21404 31214
rect 21468 30734 21496 31214
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 23032 30938 23060 31282
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23216 30734 23244 31962
rect 23400 31754 23428 32438
rect 24780 32434 24808 32914
rect 25424 32842 25452 33322
rect 28368 33114 28396 33322
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 28356 33108 28408 33114
rect 28356 33050 28408 33056
rect 25412 32836 25464 32842
rect 25412 32778 25464 32784
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 31312 32434 31340 33322
rect 33336 32434 33364 33322
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 28080 32428 28132 32434
rect 28080 32370 28132 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23388 31748 23440 31754
rect 23388 31690 23440 31696
rect 23400 30870 23428 31690
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23492 31346 23520 31622
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23388 30864 23440 30870
rect 23388 30806 23440 30812
rect 23768 30802 23796 31758
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 23756 30796 23808 30802
rect 23756 30738 23808 30744
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 21468 29510 21496 30670
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21364 29300 21416 29306
rect 21364 29242 21416 29248
rect 21652 29238 21680 29514
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 20904 27532 20956 27538
rect 20904 27474 20956 27480
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 20260 27396 20312 27402
rect 20260 27338 20312 27344
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 27130 19840 27270
rect 19800 27124 19852 27130
rect 19800 27066 19852 27072
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17144 23730 17172 24006
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 22642 17172 23666
rect 17328 23186 17356 24686
rect 17696 24154 17724 24754
rect 17960 24200 18012 24206
rect 17696 24148 17960 24154
rect 17696 24142 18012 24148
rect 17696 24126 18000 24142
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 17328 21146 17356 23122
rect 17604 23118 17632 24006
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17696 21554 17724 24126
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18156 22574 18184 22646
rect 18248 22574 18276 23802
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22166 18000 22374
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 17960 22024 18012 22030
rect 18064 21978 18092 22442
rect 18012 21972 18092 21978
rect 17960 21966 18092 21972
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 17972 21950 18092 21966
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 19854 16896 20198
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 17696 19378 17724 21490
rect 18248 21486 18276 21966
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18340 20942 18368 25638
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 18432 23866 18460 25094
rect 19352 24750 19380 26386
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18708 23322 18736 24074
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18708 22710 18736 23258
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 19248 22160 19300 22166
rect 19248 22102 19300 22108
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19168 20942 19196 21354
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 18248 18970 18276 20198
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16868 13938 16896 14962
rect 16960 14074 16988 18702
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 18524 18358 18552 18566
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17052 15910 17080 16458
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16868 13394 16896 13874
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 12238 16896 13330
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 17052 11218 17080 15846
rect 17144 15162 17172 18158
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16590 17264 17138
rect 17420 17134 17448 17614
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17420 16522 17448 17070
rect 17512 16726 17540 17478
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 18248 17270 18276 18022
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17144 11098 17172 15098
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17236 12170 17264 12718
rect 17420 12481 17448 16458
rect 17512 12986 17540 16662
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 15502 17724 16390
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 18248 16182 18276 17206
rect 18708 16522 18736 18566
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16182 18736 16458
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17604 14414 17632 15370
rect 17696 15094 17724 15438
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 13462 17632 14350
rect 17696 13938 17724 15030
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 18248 13190 18276 14962
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17406 12472 17462 12481
rect 17406 12407 17462 12416
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17236 11150 17264 12106
rect 17420 11642 17448 12407
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11762 17540 12174
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17420 11614 17540 11642
rect 17052 11070 17172 11098
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17052 9586 17080 11070
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8974 16896 9318
rect 17236 9178 17264 9590
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17328 9110 17356 9522
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16960 8090 16988 8910
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16960 7410 16988 8026
rect 17420 7478 17448 8910
rect 17512 8498 17540 11614
rect 17604 11150 17632 12786
rect 18064 12306 18092 12786
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 11286 17908 11494
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 18248 10742 18276 13126
rect 18340 11762 18368 13262
rect 18432 12918 18460 14350
rect 18800 13938 18828 20266
rect 19168 15570 19196 20878
rect 19260 20058 19288 22102
rect 19444 22030 19472 23054
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19536 21554 19564 23666
rect 19628 23254 19656 25842
rect 19812 25498 19840 27066
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23594 19748 24074
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19720 23118 19748 23530
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19996 22642 20024 23190
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19524 21548 19576 21554
rect 19352 21508 19524 21536
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19352 19174 19380 21508
rect 19524 21490 19576 21496
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 21010 19472 21286
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19628 19922 19656 21898
rect 19812 21554 19840 22374
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19996 21010 20024 22578
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19444 19718 19472 19790
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19536 19514 19564 19790
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18970 19380 19110
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 18766 19472 19382
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 18426 19472 18702
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 17218 19288 17614
rect 19260 17190 19472 17218
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19260 16250 19288 16458
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19352 15434 19380 16934
rect 19444 16572 19472 17190
rect 19536 16998 19564 18634
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19524 16584 19576 16590
rect 19444 16544 19524 16572
rect 19524 16526 19576 16532
rect 19536 16250 19564 16526
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 14346 19380 15370
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19444 14226 19472 15846
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19352 14198 19472 14226
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18340 11150 18368 11698
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8974 17632 9318
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17696 8634 17724 9114
rect 17788 8974 17816 9522
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17880 8838 17908 9454
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 18432 8634 18460 8842
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16776 6886 16896 6914
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4078 14596 4558
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14384 3862 14504 3890
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 2990 14320 3334
rect 14384 3058 14412 3862
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 3194 14780 3402
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15212 3058 15240 5170
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4214 15332 4966
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15580 4146 15608 4422
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16316 3942 16344 4422
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15672 3194 15700 3470
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14384 2650 14412 2994
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 15488 2446 15516 2926
rect 16316 2446 16344 3878
rect 16684 3602 16712 3878
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16868 3398 16896 6886
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 18248 5302 18276 7414
rect 18340 7002 18368 8502
rect 18616 7886 18644 9386
rect 18708 8974 18736 12106
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18800 7886 18828 8842
rect 19076 8294 19104 13942
rect 19352 12374 19380 14198
rect 19536 13682 19564 14282
rect 19444 13654 19564 13682
rect 19444 12918 19472 13654
rect 19628 13546 19656 19654
rect 19720 18698 19748 20198
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19812 18970 19840 19994
rect 19904 19990 19932 20538
rect 20088 20466 20116 26318
rect 20272 26314 20300 27338
rect 20916 26994 20944 27474
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20168 22704 20220 22710
rect 20168 22646 20220 22652
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19904 18630 19932 19790
rect 20088 19446 20116 20402
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19812 17270 19840 18362
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 20180 16046 20208 22646
rect 20272 21962 20300 26250
rect 20916 25294 20944 26726
rect 21180 26240 21232 26246
rect 21180 26182 21232 26188
rect 21192 25906 21220 26182
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21192 25362 21220 25842
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 20904 25288 20956 25294
rect 21284 25242 21312 28970
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 22388 28218 22416 29106
rect 22756 28422 22784 29106
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 21916 27532 21968 27538
rect 21916 27474 21968 27480
rect 21928 27334 21956 27474
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21376 26382 21404 26930
rect 21640 26852 21692 26858
rect 21640 26794 21692 26800
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 20904 25230 20956 25236
rect 21088 25220 21140 25226
rect 21088 25162 21140 25168
rect 21192 25214 21312 25242
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20640 22710 20668 24142
rect 20824 24070 20852 24754
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20916 24410 20944 24686
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 21100 24274 21128 25162
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16590 20484 16934
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20548 16250 20576 22578
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 19990 20668 20402
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20732 18766 20760 23666
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23118 20852 23598
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20916 22030 20944 23734
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21100 20806 21128 21898
rect 21192 21010 21220 25214
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24206 21312 24618
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21284 21146 21312 24142
rect 21376 23866 21404 24754
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21560 23730 21588 24550
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 21652 22166 21680 26794
rect 21928 25974 21956 27270
rect 22020 26994 22048 27406
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 21916 25968 21968 25974
rect 21916 25910 21968 25916
rect 22388 25906 22416 27270
rect 22756 26314 22784 28358
rect 22940 27062 22968 30670
rect 23216 29782 23244 30670
rect 23204 29776 23256 29782
rect 23204 29718 23256 29724
rect 24504 29170 24532 31350
rect 24596 31346 24624 32370
rect 24780 31686 24808 32370
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 25056 31890 25084 32166
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 25136 31884 25188 31890
rect 25136 31826 25188 31832
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24688 30802 24716 31350
rect 24676 30796 24728 30802
rect 24676 30738 24728 30744
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23216 28218 23244 28970
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23400 27946 23428 28494
rect 23388 27940 23440 27946
rect 23388 27882 23440 27888
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 22572 25158 22600 26250
rect 23492 25838 23520 29106
rect 24688 28490 24716 30194
rect 24780 29646 24808 31622
rect 25148 31482 25176 31826
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 26620 31482 26648 31758
rect 27724 31754 27752 32370
rect 26700 31748 26752 31754
rect 26700 31690 26752 31696
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 26608 31476 26660 31482
rect 26608 31418 26660 31424
rect 26712 31346 26740 31690
rect 27344 31476 27396 31482
rect 27344 31418 27396 31424
rect 27356 31346 27384 31418
rect 24860 31340 24912 31346
rect 25320 31340 25372 31346
rect 24860 31282 24912 31288
rect 25240 31300 25320 31328
rect 24872 29646 24900 31282
rect 25240 30802 25268 31300
rect 25320 31282 25372 31288
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 26700 31340 26752 31346
rect 26700 31282 26752 31288
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25228 30796 25280 30802
rect 25228 30738 25280 30744
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25056 30326 25084 30670
rect 25044 30320 25096 30326
rect 25044 30262 25096 30268
rect 25056 29850 25084 30262
rect 25240 30258 25268 30738
rect 25608 30734 25636 31214
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25148 29850 25176 30194
rect 25044 29844 25096 29850
rect 25044 29786 25096 29792
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 23676 28082 23704 28426
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 23584 25650 23612 25842
rect 23492 25622 23612 25650
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21652 20874 21680 22102
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20824 19786 20852 20266
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14414 19748 14758
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 13938 19748 14350
rect 19904 14278 19932 14554
rect 20272 14550 20300 16050
rect 20824 15502 20852 19722
rect 20916 18970 20944 20538
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 19514 21036 20334
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21100 19378 21128 20742
rect 21376 20534 21404 20810
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21284 19922 21312 20402
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 16114 20944 17478
rect 21192 17354 21220 19314
rect 21836 18834 21864 24346
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21928 23322 21956 23734
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21554 22324 21830
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 22388 20534 22416 21422
rect 22572 20942 22600 25094
rect 23492 24614 23520 25622
rect 24596 25294 24624 26386
rect 24688 25906 24716 27814
rect 24780 26994 24808 29582
rect 24872 27606 24900 29582
rect 25148 28778 25176 29786
rect 25240 29238 25268 30194
rect 25608 30190 25636 30670
rect 25700 30326 25728 31282
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25792 30734 25820 31078
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25688 30320 25740 30326
rect 25688 30262 25740 30268
rect 25792 30258 25820 30670
rect 26148 30660 26200 30666
rect 26148 30602 26200 30608
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 26160 30190 26188 30602
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 25596 30184 25648 30190
rect 25596 30126 25648 30132
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 25780 30116 25832 30122
rect 25780 30058 25832 30064
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 25148 28750 25268 28778
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 25056 27538 25084 28018
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25148 26994 25176 27950
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26586 25176 26930
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 23730 23520 24550
rect 23584 24290 23612 24754
rect 24596 24410 24624 25230
rect 24872 25226 24900 25842
rect 25240 25838 25268 28750
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25320 27532 25372 27538
rect 25320 27474 25372 27480
rect 25332 26382 25360 27474
rect 25424 27062 25452 28018
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 23584 24274 23888 24290
rect 23584 24268 23900 24274
rect 23584 24262 23848 24268
rect 23584 24206 23612 24262
rect 23848 24210 23900 24216
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21836 17882 21864 18770
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21100 17326 21220 17354
rect 21100 17202 21128 17326
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21100 16794 21128 17138
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21192 16454 21220 17206
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16182 21220 16390
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21652 15910 21680 16458
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19536 13518 19656 13546
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19536 12434 19564 13518
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19628 12782 19656 13330
rect 19812 13326 19840 14214
rect 19904 14074 19932 14214
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 20456 14006 20484 14758
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19904 12986 19932 13670
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19812 12442 19840 12786
rect 19800 12436 19852 12442
rect 19536 12406 19656 12434
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19352 9382 19380 12310
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 9110 19380 9318
rect 19628 9178 19656 12406
rect 19800 12378 19852 12384
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19720 12238 19748 12310
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19812 9586 19840 11630
rect 19904 11286 19932 12922
rect 20364 12850 20392 13194
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 11694 20024 12582
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19812 8362 19840 9522
rect 19904 9450 19932 11086
rect 19996 10742 20024 11630
rect 20364 11150 20392 12786
rect 20548 12170 20576 14418
rect 20824 14074 20852 14962
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20916 13734 20944 14962
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14414 21036 14758
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20718 12472 20774 12481
rect 20718 12407 20774 12416
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19996 7886 20024 8910
rect 20548 8566 20576 12106
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11354 20668 12038
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11150 20760 12407
rect 20916 12238 20944 13670
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12306 21128 12582
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20904 12232 20956 12238
rect 21192 12186 21220 14010
rect 21836 12374 21864 16050
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 22388 15638 22416 16050
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21928 12442 21956 15370
rect 22204 15026 22232 15438
rect 22480 15162 22508 16934
rect 22572 15570 22600 17070
rect 22664 16250 22692 22170
rect 23584 22094 23612 24142
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23676 23730 23704 24006
rect 24872 23730 24900 25162
rect 25148 24954 25176 25706
rect 25240 25226 25268 25774
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 23186 24992 23462
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23584 22066 23796 22094
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 22480 14618 22508 15098
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22204 13938 22232 14486
rect 22756 14346 22784 17274
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22296 13938 22324 14010
rect 22756 13954 22784 14282
rect 22480 13938 22784 13954
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22468 13932 22784 13938
rect 22520 13926 22784 13932
rect 22468 13874 22520 13880
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 22284 12844 22336 12850
rect 22336 12804 22416 12832
rect 22284 12786 22336 12792
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 20904 12174 20956 12180
rect 21008 12158 21220 12186
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11354 20944 11698
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 9466 20852 9522
rect 21008 9518 21036 12158
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21100 9586 21128 11290
rect 21376 11150 21404 11562
rect 21560 11150 21588 12174
rect 22388 11898 22416 12804
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22480 11558 22508 12718
rect 22560 12436 22612 12442
rect 22664 12434 22692 13926
rect 22848 13394 22876 16050
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22940 12986 22968 21966
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23216 19922 23244 21422
rect 23584 21146 23612 21422
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19378 23244 19858
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23400 19310 23428 20810
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23768 18766 23796 22066
rect 23860 21350 23888 22510
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24596 22030 24624 22374
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23860 20942 23888 21082
rect 23952 20942 23980 21422
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23940 20936 23992 20942
rect 24032 20936 24084 20942
rect 23940 20878 23992 20884
rect 24030 20904 24032 20913
rect 24084 20904 24086 20913
rect 24030 20839 24086 20848
rect 24780 20058 24808 21966
rect 24872 20602 24900 23054
rect 25148 22982 25176 24890
rect 25332 24818 25360 26318
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25240 24698 25268 24754
rect 25424 24698 25452 26998
rect 25608 26994 25636 27338
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25516 25974 25544 26318
rect 25504 25968 25556 25974
rect 25504 25910 25556 25916
rect 25608 25498 25636 26318
rect 25700 26042 25728 27406
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25240 24670 25452 24698
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25240 23866 25268 24142
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25332 23186 25360 24006
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 25148 21962 25176 22918
rect 25240 22710 25268 22918
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 25240 22098 25268 22646
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24952 20936 25004 20942
rect 24950 20904 24952 20913
rect 25004 20904 25006 20913
rect 24950 20839 25006 20848
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17134 23152 18158
rect 23584 17270 23612 18566
rect 23768 17814 23796 18702
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23572 17264 23624 17270
rect 23572 17206 23624 17212
rect 23768 17202 23796 17750
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 24504 16998 24532 18566
rect 24596 18290 24624 18566
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24688 17746 24716 19654
rect 24964 19446 24992 20742
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18358 24992 18566
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23308 13938 23336 16526
rect 24504 16250 24532 16934
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24596 15910 24624 16526
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 14550 23796 15302
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 23768 12782 23796 14486
rect 23860 14278 23888 15642
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 13870 23888 14214
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23952 12434 23980 15030
rect 24412 14890 24440 15370
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14074 24072 14758
rect 24596 14482 24624 15846
rect 24780 15366 24808 16934
rect 24872 16590 24900 17478
rect 25056 17202 25084 21830
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25148 18766 25176 20878
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25332 18290 25360 22986
rect 25516 20942 25544 24074
rect 25792 22506 25820 30058
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26068 28014 26096 29106
rect 26712 28626 26740 31282
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27620 30660 27672 30666
rect 27620 30602 27672 30608
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27160 29708 27212 29714
rect 27160 29650 27212 29656
rect 27172 29306 27200 29650
rect 27540 29646 27568 30194
rect 27632 29646 27660 30602
rect 27724 30326 27752 30670
rect 28092 30326 28120 32370
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 33140 32224 33192 32230
rect 33140 32166 33192 32172
rect 29092 31272 29144 31278
rect 29092 31214 29144 31220
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 27724 29782 27752 30262
rect 28460 30258 28488 30670
rect 28724 30660 28776 30666
rect 28724 30602 28776 30608
rect 28736 30258 28764 30602
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 27712 29776 27764 29782
rect 27712 29718 27764 29724
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27632 29306 27660 29582
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27172 29170 27200 29242
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 26608 28144 26660 28150
rect 26608 28086 26660 28092
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 26516 28008 26568 28014
rect 26516 27950 26568 27956
rect 25872 27940 25924 27946
rect 25872 27882 25924 27888
rect 25884 27334 25912 27882
rect 26068 27606 26096 27950
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25884 26994 25912 27270
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 26068 25702 26096 27542
rect 26528 27538 26556 27950
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27062 26188 27406
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25884 24206 25912 25638
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25780 22500 25832 22506
rect 25780 22442 25832 22448
rect 25976 22030 26004 24550
rect 26160 22574 26188 26862
rect 26620 26738 26648 28086
rect 26528 26710 26648 26738
rect 26528 26382 26556 26710
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26516 26376 26568 26382
rect 26712 26330 26740 26454
rect 26804 26382 26832 29038
rect 27356 28694 27384 29106
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27344 28688 27396 28694
rect 27344 28630 27396 28636
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 27080 27334 27108 28018
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27080 26586 27108 27270
rect 27264 26994 27292 28358
rect 27356 28150 27384 28630
rect 27344 28144 27396 28150
rect 27344 28086 27396 28092
rect 27448 26994 27476 28970
rect 27540 27470 27568 29242
rect 28092 29170 28120 30058
rect 28920 29782 28948 30670
rect 29012 30394 29040 31078
rect 29104 30802 29132 31214
rect 29092 30796 29144 30802
rect 29092 30738 29144 30744
rect 29104 30394 29132 30738
rect 29000 30388 29052 30394
rect 29000 30330 29052 30336
rect 29092 30388 29144 30394
rect 29092 30330 29144 30336
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29184 30252 29236 30258
rect 29184 30194 29236 30200
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 29012 29714 29040 30194
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29196 29646 29224 30194
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 28368 29306 28396 29582
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 28368 28626 28396 29242
rect 28920 28966 28948 29582
rect 29196 29306 29224 29582
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29656 29102 29684 30194
rect 29644 29096 29696 29102
rect 29644 29038 29696 29044
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28920 28762 28948 28902
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28356 28620 28408 28626
rect 28356 28562 28408 28568
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27724 27470 27752 28018
rect 27908 27606 27936 28494
rect 27896 27600 27948 27606
rect 27896 27542 27948 27548
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27252 26988 27304 26994
rect 27436 26988 27488 26994
rect 27252 26930 27304 26936
rect 27356 26948 27436 26976
rect 27160 26852 27212 26858
rect 27160 26794 27212 26800
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 26568 26324 26740 26330
rect 26516 26318 26740 26324
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 26528 26302 26740 26318
rect 26608 26240 26660 26246
rect 26608 26182 26660 26188
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 26620 25922 26648 26182
rect 26528 25906 26648 25922
rect 26516 25900 26648 25906
rect 26568 25894 26648 25900
rect 26516 25842 26568 25848
rect 26528 25226 26556 25842
rect 26712 25498 26740 26302
rect 26804 25974 26832 26318
rect 26792 25968 26844 25974
rect 26792 25910 26844 25916
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26608 25424 26660 25430
rect 26608 25366 26660 25372
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 26620 24682 26648 25366
rect 26608 24676 26660 24682
rect 26608 24618 26660 24624
rect 26804 24070 26832 25910
rect 26896 25906 26924 26318
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 27080 25158 27108 25774
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27080 24886 27108 25094
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 27172 24750 27200 26794
rect 27264 26042 27292 26930
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27356 25294 27384 26948
rect 27436 26930 27488 26936
rect 27540 26858 27568 27406
rect 28368 26926 28396 28562
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28736 27334 28764 28494
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 29840 26994 29868 27814
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29932 26926 29960 27406
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 29920 26920 29972 26926
rect 29920 26862 29972 26868
rect 27528 26852 27580 26858
rect 27528 26794 27580 26800
rect 28632 26512 28684 26518
rect 28632 26454 28684 26460
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27632 25838 27660 26250
rect 28644 25906 28672 26454
rect 29092 26308 29144 26314
rect 29092 26250 29144 26256
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28276 25498 28304 25774
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 28644 23798 28672 25842
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 28736 23254 28764 24754
rect 28920 24614 28948 25230
rect 29104 24818 29132 26250
rect 29932 26042 29960 26862
rect 29920 26036 29972 26042
rect 29920 25978 29972 25984
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28828 23594 28856 24550
rect 30024 24342 30052 28018
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30116 24750 30144 25230
rect 30104 24744 30156 24750
rect 30104 24686 30156 24692
rect 30012 24336 30064 24342
rect 30012 24278 30064 24284
rect 30116 23866 30144 24686
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 28724 23248 28776 23254
rect 28724 23190 28776 23196
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26976 22432 27028 22438
rect 26976 22374 27028 22380
rect 26988 22098 27016 22374
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 25964 22024 26016 22030
rect 27068 22024 27120 22030
rect 25964 21966 26016 21972
rect 26988 21972 27068 21978
rect 26988 21966 27120 21972
rect 26988 21950 27108 21966
rect 26988 21894 27016 21950
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 27080 21690 27108 21830
rect 27172 21690 27200 22578
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27068 21684 27120 21690
rect 27068 21626 27120 21632
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25884 18970 25912 21014
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 27172 18766 27200 19314
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27264 18834 27292 19110
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25700 18426 25728 18634
rect 26252 18630 26280 18702
rect 27356 18698 27384 21966
rect 27540 21962 27568 23054
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27632 22710 27660 22986
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 28092 22658 28120 23054
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27632 21486 27660 22646
rect 28092 22642 28212 22658
rect 28276 22642 28304 23054
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 28092 22636 28224 22642
rect 28092 22630 28172 22636
rect 28172 22578 28224 22584
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 28000 21554 28028 22442
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27908 20466 27936 21286
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27618 20360 27674 20369
rect 27618 20295 27620 20304
rect 27672 20295 27674 20304
rect 27620 20266 27672 20272
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27712 18896 27764 18902
rect 27712 18838 27764 18844
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27344 18692 27396 18698
rect 27344 18634 27396 18640
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25148 15706 25176 16050
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24780 13938 24808 15030
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25148 14074 25176 14962
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 22664 12406 22784 12434
rect 22560 12378 22612 12384
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20640 9438 20852 9466
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 20640 8838 20668 9438
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8566 20668 8774
rect 21008 8634 21036 8842
rect 21100 8838 21128 9522
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 21100 8498 21128 8774
rect 21192 8634 21220 9386
rect 21284 9178 21312 9590
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21376 8974 21404 9318
rect 21560 9178 21588 11086
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17052 4146 17080 4558
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4146 17540 4422
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16960 3194 16988 3402
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17604 2990 17632 4626
rect 18340 4622 18368 6938
rect 18800 6662 18828 7822
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7478 18920 7686
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 19720 6798 19748 7754
rect 19996 7478 20024 7822
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20548 7546 20576 7754
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 20640 7206 20668 8230
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 19536 6254 19564 6734
rect 20732 6730 20760 8434
rect 21100 7546 21128 8434
rect 21560 7954 21588 9114
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20916 7002 20944 7414
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20732 6458 20760 6666
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 4622 18460 6054
rect 19536 5370 19564 6190
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 20180 4622 20208 5850
rect 20916 4622 20944 6938
rect 21560 6798 21588 7890
rect 21928 6798 21956 11154
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 22480 9178 22508 9522
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22572 8566 22600 12378
rect 22756 12238 22784 12406
rect 23768 12406 23980 12434
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11830 22784 12174
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 22480 7410 22508 8502
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22572 7546 22600 8026
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22756 7410 22784 9046
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22940 7546 22968 7754
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23400 7478 23428 7958
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21284 6390 21312 6598
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 23400 5302 23428 7414
rect 23492 6866 23520 11766
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23676 11286 23704 11698
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 23768 11150 23796 12406
rect 24596 12238 24624 13874
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24688 12238 24716 12378
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 9450 23796 11086
rect 23860 10266 23888 11630
rect 24044 11150 24072 12106
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24596 11830 24624 12038
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24688 11286 24716 12174
rect 24780 12102 24808 12854
rect 25240 12434 25268 18022
rect 25056 12406 25268 12434
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11898 24808 12038
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 8634 23704 8774
rect 23768 8634 23796 9386
rect 24044 8974 24072 11086
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10742 24900 11018
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10266 24624 10542
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 25056 9382 25084 12406
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25148 10062 25176 11766
rect 25332 11558 25360 11834
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 10062 25360 11494
rect 25424 10266 25452 18158
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25700 17338 25728 17614
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25792 15570 25820 17682
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25976 17270 26004 17478
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25976 16794 26004 17206
rect 26160 17202 26188 18566
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 27540 18222 27568 18702
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27724 17678 27752 18838
rect 27908 18766 27936 19314
rect 27896 18760 27948 18766
rect 27896 18702 27948 18708
rect 27908 17746 27936 18702
rect 28000 17882 28028 20402
rect 28184 19446 28212 22578
rect 29748 22574 29776 22918
rect 29736 22568 29788 22574
rect 29736 22510 29788 22516
rect 29920 22094 29972 22098
rect 30208 22094 30236 32166
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 31128 27130 31156 28086
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32220 27396 32272 27402
rect 32220 27338 32272 27344
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 32232 26586 32260 27338
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32220 26580 32272 26586
rect 32220 26522 32272 26528
rect 32600 26382 32628 27270
rect 32692 26382 32720 28018
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 32680 26376 32732 26382
rect 32680 26318 32732 26324
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 30392 24410 30420 25162
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30944 24206 30972 25094
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 30852 22522 30880 24142
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31116 22568 31168 22574
rect 30852 22494 30972 22522
rect 31116 22510 31168 22516
rect 31208 22568 31260 22574
rect 31208 22510 31260 22516
rect 30840 22432 30892 22438
rect 30840 22374 30892 22380
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 30852 22166 30880 22374
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30840 22160 30892 22166
rect 30840 22102 30892 22108
rect 29920 22092 30236 22094
rect 29972 22066 30236 22092
rect 29920 22034 29972 22040
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 30288 21956 30340 21962
rect 30288 21898 30340 21904
rect 28460 21622 28488 21898
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28460 21010 28488 21286
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 29104 20534 29132 21626
rect 29748 21554 29776 21830
rect 30300 21690 30328 21898
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30392 21622 30420 22102
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 30944 20874 30972 22494
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21894 31064 21966
rect 31024 21888 31076 21894
rect 31024 21830 31076 21836
rect 31036 21622 31064 21830
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 31128 21554 31156 22510
rect 31220 22030 31248 22510
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 31128 21078 31156 21490
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 29092 20528 29144 20534
rect 29092 20470 29144 20476
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 26160 16658 26188 17138
rect 26620 17134 26648 17546
rect 26608 17128 26660 17134
rect 26608 17070 26660 17076
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 26068 15978 26096 16118
rect 26160 16114 26188 16390
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 26620 16114 26648 17070
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26056 15972 26108 15978
rect 26056 15914 26108 15920
rect 26068 15858 26096 15914
rect 25976 15830 26096 15858
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25792 15434 25820 15506
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25976 14618 26004 15830
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25792 12646 25820 13806
rect 26068 13326 26096 15642
rect 26160 14414 26188 15846
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14414 26464 14894
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 26620 14074 26648 16050
rect 27724 15502 27752 17614
rect 27816 17338 27844 17614
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27816 15348 27844 16390
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 28000 15706 28028 15982
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 27988 15700 28040 15706
rect 27988 15642 28040 15648
rect 28184 15570 28212 15846
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 27724 15320 27844 15348
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25688 12368 25740 12374
rect 25688 12310 25740 12316
rect 25700 11830 25728 12310
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 25792 11558 25820 12582
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 25976 10810 26004 11154
rect 26068 11150 26096 11494
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25148 9654 25176 9998
rect 25976 9994 26004 10746
rect 26620 10062 26648 10950
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25136 9648 25188 9654
rect 25136 9590 25188 9596
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24044 7886 24072 8298
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24688 7546 24716 8502
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23492 6186 23520 6802
rect 24688 6798 24716 7482
rect 24872 7478 24900 8910
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 8498 24992 8774
rect 25240 8634 25268 9930
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 25148 6798 25176 8298
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23584 6390 23612 6598
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5710 24716 6054
rect 25608 5710 25636 7142
rect 25884 6662 25912 8570
rect 25976 7546 26004 9522
rect 26712 9042 26740 12786
rect 26804 11354 26832 13874
rect 26884 13864 26936 13870
rect 26884 13806 26936 13812
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26056 8900 26108 8906
rect 26056 8842 26108 8848
rect 26068 8498 26096 8842
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25976 5914 26004 7482
rect 26068 7410 26096 8434
rect 26896 8090 26924 13806
rect 26988 13530 27016 14350
rect 27540 14074 27568 14350
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27724 14006 27752 15320
rect 27804 14272 27856 14278
rect 27804 14214 27856 14220
rect 27712 14000 27764 14006
rect 27712 13942 27764 13948
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27632 13802 27660 13874
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27816 12986 27844 14214
rect 28092 14074 28120 15438
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 27988 14000 28040 14006
rect 27908 13960 27988 13988
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 10606 27384 11630
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27356 10266 27384 10542
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 27724 10062 27752 12650
rect 27908 12374 27936 13960
rect 27988 13942 28040 13948
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 28184 13802 28212 13874
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 27896 12368 27948 12374
rect 27896 12310 27948 12316
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26068 7002 26096 7346
rect 27632 7342 27660 8910
rect 27908 8294 27936 11698
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27908 7546 27936 8230
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 24688 5370 24716 5646
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 18248 4214 18276 4422
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 19076 3942 19104 4422
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 18248 3194 18276 3334
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 18248 2514 18276 3130
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19076 2446 19104 3878
rect 19720 3534 19748 4422
rect 20640 3738 20668 4422
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 20640 2446 20668 3674
rect 20732 3194 20760 4082
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20812 3052 20864 3058
rect 20916 3040 20944 4558
rect 21008 3058 21036 4694
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3194 21128 3878
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20864 3012 20944 3040
rect 20996 3052 21048 3058
rect 20812 2994 20864 3000
rect 20996 2994 21048 3000
rect 21100 2446 21128 3130
rect 21192 3058 21220 4626
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21560 4146 21588 4422
rect 22112 4146 22140 4422
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22296 4026 22324 4082
rect 22296 3998 22416 4026
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 22388 3738 22416 3998
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22480 3534 22508 4762
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24412 4214 24440 4558
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24596 4146 24624 4422
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22756 3058 22784 3538
rect 23400 3534 23428 3878
rect 24688 3738 24716 4694
rect 25056 4690 25084 5102
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 23400 2446 23428 3470
rect 25056 2990 25084 3674
rect 25700 3534 25728 4966
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25792 3482 25820 5170
rect 26700 5160 26752 5166
rect 26700 5102 26752 5108
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25976 4214 26004 4558
rect 26608 4548 26660 4554
rect 26608 4490 26660 4496
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 26620 4282 26648 4490
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 25964 4208 26016 4214
rect 25964 4150 26016 4156
rect 25976 3602 26004 4150
rect 26712 4078 26740 5102
rect 27172 4622 27200 6938
rect 28000 6866 28028 12854
rect 28092 12434 28120 13330
rect 28092 12406 28212 12434
rect 28184 12238 28212 12406
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28184 10674 28212 12174
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28276 10266 28304 20198
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28552 18766 28580 19246
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28368 18290 28396 18566
rect 28448 18352 28500 18358
rect 28448 18294 28500 18300
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28368 13802 28396 16458
rect 28460 16454 28488 18294
rect 28552 18154 28580 18702
rect 28540 18148 28592 18154
rect 28540 18090 28592 18096
rect 28644 18034 28672 18702
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28552 18006 28672 18034
rect 28552 17678 28580 18006
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28552 17202 28580 17614
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28736 16522 28764 18226
rect 29012 18222 29040 19314
rect 29104 18834 29132 20470
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 29104 18290 29132 18770
rect 29196 18290 29224 19450
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29288 18766 29316 19246
rect 29276 18760 29328 18766
rect 29276 18702 29328 18708
rect 29380 18698 29408 19314
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29840 18306 29868 18702
rect 29748 18290 29868 18306
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29736 18284 29868 18290
rect 29788 18278 29868 18284
rect 29736 18226 29788 18232
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29012 17882 29040 18158
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17338 28856 17478
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28920 17202 28948 17614
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 29748 16658 29776 18226
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30944 17338 30972 17614
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 30012 17332 30064 17338
rect 30012 17274 30064 17280
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30024 16658 30052 17274
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 28920 16538 28948 16594
rect 28724 16516 28776 16522
rect 28920 16510 29040 16538
rect 28724 16458 28776 16464
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28460 16114 28488 16390
rect 28736 16250 28764 16458
rect 28724 16244 28776 16250
rect 28724 16186 28776 16192
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28356 13796 28408 13802
rect 28356 13738 28408 13744
rect 28368 12850 28396 13738
rect 28460 12986 28488 15438
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28368 11830 28396 12582
rect 28552 12442 28580 14350
rect 28920 13938 28948 16050
rect 29012 15026 29040 16510
rect 29104 16114 29132 16594
rect 30024 16454 30052 16594
rect 30300 16454 30328 17070
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 31128 16794 31156 17546
rect 31312 17202 31340 19314
rect 31404 19242 31432 23122
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31588 20602 31616 21966
rect 31772 21690 31800 23054
rect 31864 22778 31892 23258
rect 31852 22772 31904 22778
rect 31852 22714 31904 22720
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31956 21146 31984 25842
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32324 24818 32352 25638
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32416 24274 32444 26318
rect 32692 26234 32720 26318
rect 32692 26206 32812 26234
rect 32784 25906 32812 26206
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32692 24682 32720 25842
rect 32680 24676 32732 24682
rect 32680 24618 32732 24624
rect 32404 24268 32456 24274
rect 32404 24210 32456 24216
rect 32784 24206 32812 25842
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 33152 23322 33180 32166
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 32680 23180 32732 23186
rect 32680 23122 32732 23128
rect 33140 23180 33192 23186
rect 33140 23122 33192 23128
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32048 22778 32076 23054
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32416 22574 32444 23054
rect 32692 22642 32720 23122
rect 33152 22710 33180 23122
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32416 22030 32444 22510
rect 33152 22098 33180 22646
rect 33336 22574 33364 23054
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33520 22710 33548 22918
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 33508 22704 33560 22710
rect 33508 22646 33560 22652
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33336 22030 33364 22510
rect 33704 22234 33732 22578
rect 33692 22228 33744 22234
rect 33692 22170 33744 22176
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32416 21146 32444 21966
rect 32600 21554 32628 21966
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 32140 20534 32168 20878
rect 32128 20528 32180 20534
rect 32324 20482 32352 20878
rect 32600 20602 32628 21490
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32772 20868 32824 20874
rect 32772 20810 32824 20816
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32128 20470 32180 20476
rect 31944 20392 31996 20398
rect 31944 20334 31996 20340
rect 31956 19854 31984 20334
rect 32140 19922 32168 20470
rect 32232 20454 32352 20482
rect 32784 20466 32812 20810
rect 32496 20460 32548 20466
rect 32128 19916 32180 19922
rect 32128 19858 32180 19864
rect 32232 19854 32260 20454
rect 32496 20402 32548 20408
rect 32772 20460 32824 20466
rect 32772 20402 32824 20408
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32324 19990 32352 20266
rect 32312 19984 32364 19990
rect 32312 19926 32364 19932
rect 32508 19854 32536 20402
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 32496 19848 32548 19854
rect 32496 19790 32548 19796
rect 31956 19378 31984 19790
rect 32232 19446 32260 19790
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 31392 19236 31444 19242
rect 31392 19178 31444 19184
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 32232 17490 32260 19382
rect 32416 19378 32444 19790
rect 32508 19514 32536 19790
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32508 18834 32536 19450
rect 32784 18850 32812 20402
rect 32968 20330 32996 20878
rect 33048 20868 33100 20874
rect 33048 20810 33100 20816
rect 33060 20466 33088 20810
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32956 20324 33008 20330
rect 32956 20266 33008 20272
rect 33060 19514 33088 20402
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 33336 18970 33364 21966
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 32496 18828 32548 18834
rect 32496 18770 32548 18776
rect 32588 18828 32640 18834
rect 32784 18822 32904 18850
rect 32588 18770 32640 18776
rect 32404 18692 32456 18698
rect 32404 18634 32456 18640
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32324 17814 32352 18158
rect 32312 17808 32364 17814
rect 32312 17750 32364 17756
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31312 16726 31340 17138
rect 31300 16720 31352 16726
rect 31300 16662 31352 16668
rect 31312 16590 31340 16662
rect 31404 16658 31432 17138
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30116 16182 30144 16390
rect 30104 16176 30156 16182
rect 30104 16118 30156 16124
rect 30300 16114 30328 16390
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15570 29500 15846
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28540 12436 28592 12442
rect 28540 12378 28592 12384
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28460 11898 28488 12106
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28460 11506 28488 11834
rect 28552 11694 28580 12378
rect 28644 12238 28672 13806
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28736 12306 28764 12786
rect 28920 12714 28948 13670
rect 28908 12708 28960 12714
rect 28908 12650 28960 12656
rect 28920 12434 28948 12650
rect 28920 12406 29224 12434
rect 28724 12300 28776 12306
rect 28724 12242 28776 12248
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28736 11898 28764 12242
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28460 11478 28580 11506
rect 28264 10260 28316 10266
rect 28264 10202 28316 10208
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28460 10062 28488 10202
rect 28552 10130 28580 11478
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 29012 10742 29040 10950
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28540 10124 28592 10130
rect 28540 10066 28592 10072
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28736 9994 28764 10610
rect 29104 10130 29132 10746
rect 29196 10470 29224 12406
rect 29564 11150 29592 15370
rect 30840 15088 30892 15094
rect 30840 15030 30892 15036
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29656 13938 29684 14826
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29748 13938 29776 14282
rect 29932 14074 29960 14962
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 30852 14074 30880 15030
rect 31312 14278 31340 16526
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 31772 14482 31800 15642
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29656 12850 29684 13874
rect 30380 13796 30432 13802
rect 30380 13738 30432 13744
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30208 11762 30236 12718
rect 30392 12170 30420 13738
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 30852 12434 30880 14010
rect 31312 13954 31340 14010
rect 31312 13938 31432 13954
rect 31312 13932 31444 13938
rect 31312 13926 31392 13932
rect 31392 13874 31444 13880
rect 31956 12850 31984 17478
rect 32232 17462 32352 17490
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 32232 16794 32260 17274
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32324 16658 32352 17462
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32416 16590 32444 18634
rect 32508 18290 32536 18770
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32508 17184 32536 18226
rect 32600 17678 32628 18770
rect 32876 18766 32904 18822
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32876 18426 32904 18702
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 32864 18420 32916 18426
rect 32864 18362 32916 18368
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 35072 18216 35124 18222
rect 35072 18158 35124 18164
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32876 17338 32904 18158
rect 35084 17921 35112 18158
rect 35070 17912 35126 17921
rect 35070 17847 35126 17856
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33428 17338 33456 17614
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33416 17332 33468 17338
rect 33416 17274 33468 17280
rect 32588 17196 32640 17202
rect 32508 17156 32588 17184
rect 32588 17138 32640 17144
rect 32600 16998 32628 17138
rect 32588 16992 32640 16998
rect 32588 16934 32640 16940
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 32416 16114 32444 16526
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32312 16040 32364 16046
rect 32312 15982 32364 15988
rect 32324 15706 32352 15982
rect 32312 15700 32364 15706
rect 32312 15642 32364 15648
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 32140 12986 32168 14350
rect 32324 13870 32352 14418
rect 32600 14074 32628 16934
rect 32772 16652 32824 16658
rect 32772 16594 32824 16600
rect 32784 16250 32812 16594
rect 34713 16348 35021 16357
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 13530 32352 13806
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 31944 12844 31996 12850
rect 31944 12786 31996 12792
rect 30852 12406 30972 12434
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 30208 11150 30236 11698
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 29368 10736 29420 10742
rect 29368 10678 29420 10684
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 29092 10124 29144 10130
rect 29092 10066 29144 10072
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 9586 28764 9930
rect 28920 9722 28948 9998
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28184 7546 28212 8434
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 7750 28396 8366
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 27988 6860 28040 6866
rect 27988 6802 28040 6808
rect 28368 6322 28396 7686
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 28736 5302 28764 8774
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 28816 7812 28868 7818
rect 28816 7754 28868 7760
rect 28828 7342 28856 7754
rect 28816 7336 28868 7342
rect 28816 7278 28868 7284
rect 28724 5296 28776 5302
rect 28724 5238 28776 5244
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26700 4072 26752 4078
rect 26700 4014 26752 4020
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26240 3664 26292 3670
rect 26160 3612 26240 3618
rect 26160 3606 26292 3612
rect 25964 3596 26016 3602
rect 25964 3538 26016 3544
rect 26160 3590 26280 3606
rect 26160 3482 26188 3590
rect 26620 3534 26648 3878
rect 25792 3454 26188 3482
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25056 2446 25084 2926
rect 25792 2854 25820 3454
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 26620 2854 26648 3470
rect 26712 3126 26740 4014
rect 26804 3738 26832 4422
rect 27172 4146 27200 4558
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27436 4140 27488 4146
rect 27436 4082 27488 4088
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 26804 2922 26832 3674
rect 27448 3194 27476 4082
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28368 3670 28396 3878
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 26792 2916 26844 2922
rect 26792 2858 26844 2864
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26252 2446 26280 2790
rect 27172 2446 27200 2790
rect 28368 2446 28396 3606
rect 28828 3126 28856 7278
rect 28920 6390 28948 8434
rect 29012 7410 29040 8910
rect 29104 8838 29132 9862
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29196 8090 29224 10406
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29380 7818 29408 10678
rect 29840 9625 29868 11086
rect 30104 11008 30156 11014
rect 30104 10950 30156 10956
rect 30116 10810 30144 10950
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 29826 9616 29882 9625
rect 29826 9551 29882 9560
rect 29840 9042 29868 9551
rect 29828 9036 29880 9042
rect 29828 8978 29880 8984
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29368 7812 29420 7818
rect 29368 7754 29420 7760
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29380 7002 29408 7754
rect 29368 6996 29420 7002
rect 29368 6938 29420 6944
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 28908 6384 28960 6390
rect 28908 6326 28960 6332
rect 29196 5234 29224 6734
rect 29748 5370 29776 8774
rect 29932 7818 29960 10202
rect 30208 9586 30236 11086
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 30196 9580 30248 9586
rect 30196 9522 30248 9528
rect 30208 8974 30236 9522
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 29920 7812 29972 7818
rect 29920 7754 29972 7760
rect 30024 6458 30052 8502
rect 30208 6798 30236 8910
rect 30300 8566 30328 9998
rect 30288 8560 30340 8566
rect 30288 8502 30340 8508
rect 30392 8498 30420 10066
rect 30852 9654 30880 10406
rect 30944 10130 30972 12406
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11898 31248 12038
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31220 11354 31248 11834
rect 31404 11762 31432 12106
rect 32692 11898 32720 15574
rect 32784 15366 32812 16186
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33888 15706 33916 16050
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32772 13728 32824 13734
rect 32876 13682 32904 15438
rect 32956 15428 33008 15434
rect 32956 15370 33008 15376
rect 32968 15162 32996 15370
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 32956 15156 33008 15162
rect 32956 15098 33008 15104
rect 32824 13676 32904 13682
rect 32772 13670 32904 13676
rect 32784 13654 32904 13670
rect 32876 12850 32904 13654
rect 32968 13326 32996 15098
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 33244 12986 33272 14214
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 33232 12980 33284 12986
rect 33232 12922 33284 12928
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 33416 11756 33468 11762
rect 33416 11698 33468 11704
rect 32496 11620 32548 11626
rect 32496 11562 32548 11568
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 31208 11348 31260 11354
rect 31208 11290 31260 11296
rect 32312 11076 32364 11082
rect 32312 11018 32364 11024
rect 32324 10606 32352 11018
rect 32416 10674 32444 11494
rect 32508 11082 32536 11562
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32324 10266 32352 10542
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 33428 10062 33456 11698
rect 33704 10810 33732 11834
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 31220 9489 31248 9930
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 31482 9616 31538 9625
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 31392 9580 31444 9586
rect 31482 9551 31484 9560
rect 31392 9522 31444 9528
rect 31536 9551 31538 9560
rect 31484 9522 31536 9528
rect 31206 9480 31262 9489
rect 31206 9415 31262 9424
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 31220 7886 31248 9415
rect 31312 8498 31340 9522
rect 31404 9450 31432 9522
rect 31942 9480 31998 9489
rect 31392 9444 31444 9450
rect 31942 9415 31944 9424
rect 31392 9386 31444 9392
rect 31996 9415 31998 9424
rect 31944 9386 31996 9392
rect 31404 8634 31432 9386
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31772 8566 31800 9318
rect 33704 9178 33732 9862
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 33888 8974 33916 9862
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 31760 8560 31812 8566
rect 31760 8502 31812 8508
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 32324 8430 32352 8910
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 32312 8424 32364 8430
rect 32312 8366 32364 8372
rect 32324 8090 32352 8366
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30576 7478 30604 7686
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 30564 7472 30616 7478
rect 30564 7414 30616 7420
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 30012 6452 30064 6458
rect 30012 6394 30064 6400
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 29932 3194 29960 5170
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 25688 2372 25740 2378
rect 25688 2314 25740 2320
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 14108 800 14136 2314
rect 15396 800 15424 2314
rect 16684 800 16712 2314
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 17972 870 18092 898
rect 17972 800 18000 870
rect 3896 734 4200 762
rect 5078 0 5134 800
rect 6366 0 6422 800
rect 7654 0 7710 800
rect 8942 0 8998 800
rect 10230 0 10286 800
rect 11518 0 11574 800
rect 12806 0 12862 800
rect 14094 0 14150 800
rect 15382 0 15438 800
rect 16670 0 16726 800
rect 17958 0 18014 800
rect 18064 762 18092 870
rect 18248 762 18276 2314
rect 19352 898 19380 2314
rect 20732 898 20760 2314
rect 22112 898 22140 2314
rect 19260 870 19380 898
rect 20548 870 20760 898
rect 21836 870 22140 898
rect 23124 870 23244 898
rect 19260 800 19288 870
rect 20548 800 20576 870
rect 21836 800 21864 870
rect 23124 800 23152 870
rect 18064 734 18276 762
rect 19246 0 19302 800
rect 20534 0 20590 800
rect 21822 0 21878 800
rect 23110 0 23166 800
rect 23216 762 23244 870
rect 23492 762 23520 2314
rect 24412 800 24440 2314
rect 25700 800 25728 2314
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 26988 800 27016 2314
rect 28276 800 28304 2314
rect 29564 800 29592 2382
rect 30852 800 30880 2382
rect 32140 800 32168 2382
rect 33428 800 33456 2382
rect 34612 2304 34664 2310
rect 34612 2246 34664 2252
rect 34624 1170 34652 2246
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 34624 1142 34744 1170
rect 34716 800 34744 1142
rect 23216 734 23520 762
rect 24398 0 24454 800
rect 25686 0 25742 800
rect 26974 0 27030 800
rect 28262 0 28318 800
rect 29550 0 29606 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
<< via2 >>
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 14830 20304 14886 20360
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 17406 12416 17462 12472
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 20718 12416 20774 12472
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 24030 20884 24032 20904
rect 24032 20884 24084 20904
rect 24084 20884 24086 20904
rect 24030 20848 24086 20884
rect 24950 20884 24952 20904
rect 24952 20884 25004 20904
rect 25004 20884 25006 20904
rect 24950 20848 25006 20884
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 27618 20324 27674 20360
rect 27618 20304 27620 20324
rect 27620 20304 27672 20324
rect 27672 20304 27674 20324
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 35070 17856 35126 17912
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 29826 9560 29882 9616
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 31482 9580 31538 9616
rect 31482 9560 31484 9580
rect 31484 9560 31536 9580
rect 31536 9560 31538 9580
rect 31206 9424 31262 9480
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 31942 9444 31998 9480
rect 31942 9424 31944 9444
rect 31944 9424 31996 9444
rect 31996 9424 31998 9444
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
<< metal3 >>
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 24025 20906 24091 20909
rect 24945 20906 25011 20909
rect 24025 20904 25011 20906
rect 24025 20848 24030 20904
rect 24086 20848 24950 20904
rect 25006 20848 25011 20904
rect 24025 20846 25011 20848
rect 24025 20843 24091 20846
rect 24945 20843 25011 20846
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 14825 20362 14891 20365
rect 27613 20362 27679 20365
rect 14825 20360 27679 20362
rect 14825 20304 14830 20360
rect 14886 20304 27618 20360
rect 27674 20304 27679 20360
rect 14825 20302 27679 20304
rect 14825 20299 14891 20302
rect 27613 20299 27679 20302
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 35065 17914 35131 17917
rect 35200 17914 36000 17944
rect 35065 17912 36000 17914
rect 35065 17856 35070 17912
rect 35126 17856 36000 17912
rect 35065 17854 36000 17856
rect 35065 17851 35131 17854
rect 35200 17824 36000 17854
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 17401 12474 17467 12477
rect 20713 12474 20779 12477
rect 17401 12472 20779 12474
rect 17401 12416 17406 12472
rect 17462 12416 20718 12472
rect 20774 12416 20779 12472
rect 17401 12414 20779 12416
rect 17401 12411 17467 12414
rect 20713 12411 20779 12414
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 29821 9618 29887 9621
rect 31477 9618 31543 9621
rect 29821 9616 31543 9618
rect 29821 9560 29826 9616
rect 29882 9560 31482 9616
rect 31538 9560 31543 9616
rect 29821 9558 31543 9560
rect 29821 9555 29887 9558
rect 31477 9555 31543 9558
rect 31201 9482 31267 9485
rect 31937 9482 32003 9485
rect 31201 9480 32003 9482
rect 31201 9424 31206 9480
rect 31262 9424 31942 9480
rect 31998 9424 32003 9480
rect 31201 9422 32003 9424
rect 31201 9419 31267 9422
rect 31937 9419 32003 9422
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
<< via3 >>
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 33216 5484 33776
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 33760 9704 33776
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 33216 13925 33776
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 33760 18145 33776
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 33216 22366 33776
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 33760 26586 33776
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 26266 22880 26586 23904
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 33216 30807 33776
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30487 28864 30807 29888
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 30487 15808 30807 16832
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 30487 12544 30807 13568
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 33760 35027 33776
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1676037725
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155
timestamp 1676037725
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1676037725
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1676037725
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_211
timestamp 1676037725
transform 1 0 20516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1676037725
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 1676037725
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1676037725
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_267
timestamp 1676037725
transform 1 0 25668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1676037725
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_295
timestamp 1676037725
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp 1676037725
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1676037725
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_322
timestamp 1676037725
transform 1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 1676037725
transform 1 0 32568 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_350
timestamp 1676037725
transform 1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1676037725
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_126
timestamp 1676037725
transform 1 0 12696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1676037725
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp 1676037725
transform 1 0 19780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1676037725
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_289
timestamp 1676037725
transform 1 0 27692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1676037725
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1676037725
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1676037725
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1676037725
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1676037725
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1676037725
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1676037725
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_286
timestamp 1676037725
transform 1 0 27416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1676037725
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1676037725
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1676037725
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_128
timestamp 1676037725
transform 1 0 12880 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_138
timestamp 1676037725
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_174
timestamp 1676037725
transform 1 0 17112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1676037725
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1676037725
transform 1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_251
timestamp 1676037725
transform 1 0 24196 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1676037725
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1676037725
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_299
timestamp 1676037725
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1676037725
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1676037725
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_107
timestamp 1676037725
transform 1 0 10948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1676037725
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_147
timestamp 1676037725
transform 1 0 14628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_155
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp 1676037725
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1676037725
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_212
timestamp 1676037725
transform 1 0 20608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_220
timestamp 1676037725
transform 1 0 21344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1676037725
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_231
timestamp 1676037725
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1676037725
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_261
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_269
timestamp 1676037725
transform 1 0 25852 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_287
timestamp 1676037725
transform 1 0 27508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_299
timestamp 1676037725
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1676037725
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1676037725
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1676037725
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_156
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1676037725
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1676037725
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1676037725
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1676037725
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1676037725
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_312
timestamp 1676037725
transform 1 0 29808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1676037725
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_55
timestamp 1676037725
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_67
timestamp 1676037725
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1676037725
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_147
timestamp 1676037725
transform 1 0 14628 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_155
timestamp 1676037725
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1676037725
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_283
timestamp 1676037725
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_295
timestamp 1676037725
transform 1 0 28244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1676037725
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_68
timestamp 1676037725
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_80
timestamp 1676037725
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1676037725
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1676037725
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_134
timestamp 1676037725
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1676037725
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1676037725
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_260
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_272
timestamp 1676037725
transform 1 0 26128 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_315
timestamp 1676037725
transform 1 0 30084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_327
timestamp 1676037725
transform 1 0 31188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1676037725
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1676037725
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1676037725
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_174
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1676037725
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_225
timestamp 1676037725
transform 1 0 21804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_237
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_271
timestamp 1676037725
transform 1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_283
timestamp 1676037725
transform 1 0 27140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1676037725
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_317
timestamp 1676037725
transform 1 0 30268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_329
timestamp 1676037725
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_341
timestamp 1676037725
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp 1676037725
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1676037725
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_30
timestamp 1676037725
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1676037725
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1676037725
transform 1 0 8372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_138
timestamp 1676037725
transform 1 0 13800 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1676037725
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1676037725
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1676037725
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1676037725
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1676037725
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_295
timestamp 1676037725
transform 1 0 28244 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1676037725
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_61
timestamp 1676037725
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_69
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1676037725
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_99
timestamp 1676037725
transform 1 0 10212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_111
timestamp 1676037725
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1676037725
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1676037725
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_227
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1676037725
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_275
timestamp 1676037725
transform 1 0 26404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1676037725
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_317
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_325
timestamp 1676037725
transform 1 0 31004 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_347
timestamp 1676037725
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1676037725
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1676037725
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_233
timestamp 1676037725
transform 1 0 22540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1676037725
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1676037725
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_312
timestamp 1676037725
transform 1 0 29808 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1676037725
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_355
timestamp 1676037725
transform 1 0 33764 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_49
timestamp 1676037725
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1676037725
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1676037725
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_220
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1676037725
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_261
timestamp 1676037725
transform 1 0 25116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_273
timestamp 1676037725
transform 1 0 26220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_285
timestamp 1676037725
transform 1 0 27324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_297
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1676037725
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_94
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1676037725
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_177
timestamp 1676037725
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_189
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_206
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_245
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_257
timestamp 1676037725
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1676037725
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1676037725
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_290
timestamp 1676037725
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_302
timestamp 1676037725
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_314
timestamp 1676037725
transform 1 0 29992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_326
timestamp 1676037725
transform 1 0 31096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_360
timestamp 1676037725
transform 1 0 34224 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1676037725
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1676037725
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_126
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1676037725
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_267
timestamp 1676037725
transform 1 0 25668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1676037725
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_318
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1676037725
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_347
timestamp 1676037725
transform 1 0 33028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_19
timestamp 1676037725
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_34
timestamp 1676037725
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1676037725
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1676037725
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_100
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_152
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1676037725
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1676037725
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_301
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_313
timestamp 1676037725
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1676037725
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_355
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_363
timestamp 1676037725
transform 1 0 34500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_36
timestamp 1676037725
transform 1 0 4416 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_64
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1676037725
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1676037725
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1676037725
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1676037725
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_184
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_212
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_222
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_234
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_242
timestamp 1676037725
transform 1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_291
timestamp 1676037725
transform 1 0 27876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1676037725
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_317
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1676037725
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1676037725
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_238
timestamp 1676037725
transform 1 0 23000 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_246
timestamp 1676037725
transform 1 0 23736 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1676037725
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_301
timestamp 1676037725
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_313
timestamp 1676037725
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_325
timestamp 1676037725
transform 1 0 31004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1676037725
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_345
timestamp 1676037725
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_357
timestamp 1676037725
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_363
timestamp 1676037725
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1676037725
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1676037725
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_205
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_273
timestamp 1676037725
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_285
timestamp 1676037725
transform 1 0 27324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_291
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1676037725
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_238
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_250
timestamp 1676037725
transform 1 0 24104 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1676037725
transform 1 0 27968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_302
timestamp 1676037725
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_312
timestamp 1676037725
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_324
timestamp 1676037725
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_345
timestamp 1676037725
transform 1 0 32844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_357
timestamp 1676037725
transform 1 0 33948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1676037725
transform 1 0 34500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1676037725
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1676037725
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1676037725
transform 1 0 5152 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_50
timestamp 1676037725
transform 1 0 5704 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_62
timestamp 1676037725
transform 1 0 6808 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_74
timestamp 1676037725
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1676037725
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_171
timestamp 1676037725
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 1676037725
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_228
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1676037725
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1676037725
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1676037725
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_18
timestamp 1676037725
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1676037725
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_65
timestamp 1676037725
transform 1 0 7084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_77
timestamp 1676037725
transform 1 0 8188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_96
timestamp 1676037725
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_146
timestamp 1676037725
transform 1 0 14536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_154
timestamp 1676037725
transform 1 0 15272 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1676037725
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1676037725
transform 1 0 22632 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_242
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_299
timestamp 1676037725
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1676037725
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_316
timestamp 1676037725
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_358
timestamp 1676037725
transform 1 0 34040 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1676037725
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_96
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1676037725
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1676037725
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1676037725
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1676037725
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_330
timestamp 1676037725
transform 1 0 31464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1676037725
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1676037725
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_34
timestamp 1676037725
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1676037725
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1676037725
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_265
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1676037725
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_309
timestamp 1676037725
transform 1 0 29532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1676037725
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1676037725
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_359
timestamp 1676037725
transform 1 0 34132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_363
timestamp 1676037725
transform 1 0 34500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_48
timestamp 1676037725
transform 1 0 5520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1676037725
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1676037725
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1676037725
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_94
timestamp 1676037725
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_110
timestamp 1676037725
transform 1 0 11224 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1676037725
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_155
timestamp 1676037725
transform 1 0 15364 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_234
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_242
timestamp 1676037725
transform 1 0 23368 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_282
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_290
timestamp 1676037725
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_347
timestamp 1676037725
transform 1 0 33028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1676037725
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_62
timestamp 1676037725
transform 1 0 6808 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_70
timestamp 1676037725
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_136
timestamp 1676037725
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_235
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_262
timestamp 1676037725
transform 1 0 25208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_270
timestamp 1676037725
transform 1 0 25944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1676037725
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_310
timestamp 1676037725
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_322
timestamp 1676037725
transform 1 0 30728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_356
timestamp 1676037725
transform 1 0 33856 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_36
timestamp 1676037725
transform 1 0 4416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_54
timestamp 1676037725
transform 1 0 6072 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_100
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_112
timestamp 1676037725
transform 1 0 11408 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1676037725
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1676037725
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1676037725
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_223
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_235
timestamp 1676037725
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1676037725
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_281
timestamp 1676037725
transform 1 0 26956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1676037725
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1676037725
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_319
timestamp 1676037725
transform 1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1676037725
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1676037725
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_37
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1676037725
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 1676037725
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1676037725
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_98
timestamp 1676037725
transform 1 0 10120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_136
timestamp 1676037725
transform 1 0 13616 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1676037725
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1676037725
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_297
timestamp 1676037725
transform 1 0 28428 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_302
timestamp 1676037725
transform 1 0 28888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_318
timestamp 1676037725
transform 1 0 30360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_326
timestamp 1676037725
transform 1 0 31096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_344
timestamp 1676037725
transform 1 0 32752 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_351
timestamp 1676037725
transform 1 0 33396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1676037725
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_60
timestamp 1676037725
transform 1 0 6624 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_72
timestamp 1676037725
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_187
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1676037725
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_225
timestamp 1676037725
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1676037725
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_261
timestamp 1676037725
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_273
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_285
timestamp 1676037725
transform 1 0 27324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1676037725
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1676037725
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_321
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_327
timestamp 1676037725
transform 1 0 31188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_336
timestamp 1676037725
transform 1 0 32016 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1676037725
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_78
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1676037725
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1676037725
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1676037725
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1676037725
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1676037725
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_315
timestamp 1676037725
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1676037725
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_346
timestamp 1676037725
transform 1 0 32936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_358
timestamp 1676037725
transform 1 0 34040 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_362
timestamp 1676037725
transform 1 0 34408 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_104
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1676037725
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_123
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_150
timestamp 1676037725
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_182
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_227
timestamp 1676037725
transform 1 0 21988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1676037725
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1676037725
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_261
timestamp 1676037725
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_276
timestamp 1676037725
transform 1 0 26496 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_316
timestamp 1676037725
transform 1 0 30176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_328
timestamp 1676037725
transform 1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_349
timestamp 1676037725
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1676037725
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1676037725
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1676037725
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1676037725
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_139
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_147
timestamp 1676037725
transform 1 0 14628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_177
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1676037725
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1676037725
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1676037725
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_286
timestamp 1676037725
transform 1 0 27416 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_294
timestamp 1676037725
transform 1 0 28152 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_322
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_331
timestamp 1676037725
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_346
timestamp 1676037725
transform 1 0 32936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 1676037725
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_39
timestamp 1676037725
transform 1 0 4692 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1676037725
transform 1 0 6532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1676037725
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_91
timestamp 1676037725
transform 1 0 9476 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_118
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_130
timestamp 1676037725
transform 1 0 13064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1676037725
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_185
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_207
timestamp 1676037725
transform 1 0 20148 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_234
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1676037725
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_19
timestamp 1676037725
transform 1 0 2852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1676037725
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1676037725
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1676037725
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1676037725
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_202
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_210
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1676037725
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_260
timestamp 1676037725
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_348
timestamp 1676037725
transform 1 0 33120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1676037725
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 1676037725
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_149
timestamp 1676037725
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1676037725
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_234
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_242
timestamp 1676037725
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_261
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_273
timestamp 1676037725
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_285
timestamp 1676037725
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1676037725
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1676037725
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1676037725
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_349
timestamp 1676037725
transform 1 0 33212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1676037725
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1676037725
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1676037725
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_120
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_144
timestamp 1676037725
transform 1 0 14352 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_232
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_259
timestamp 1676037725
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1676037725
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1676037725
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_309
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_315
timestamp 1676037725
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_320
timestamp 1676037725
transform 1 0 30544 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_328
timestamp 1676037725
transform 1 0 31280 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1676037725
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_68
timestamp 1676037725
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_76
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1676037725
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1676037725
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_263
timestamp 1676037725
transform 1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_274
timestamp 1676037725
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1676037725
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 1676037725
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1676037725
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_347
timestamp 1676037725
transform 1 0 33028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1676037725
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1676037725
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1676037725
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1676037725
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1676037725
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_122
timestamp 1676037725
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_140
timestamp 1676037725
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_158
timestamp 1676037725
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_175
timestamp 1676037725
transform 1 0 17204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1676037725
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1676037725
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_242
timestamp 1676037725
transform 1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1676037725
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_307
timestamp 1676037725
transform 1 0 29348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_316
timestamp 1676037725
transform 1 0 30176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_322
timestamp 1676037725
transform 1 0 30728 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1676037725
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_359
timestamp 1676037725
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_36
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_48
timestamp 1676037725
transform 1 0 5520 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_60
timestamp 1676037725
transform 1 0 6624 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_71
timestamp 1676037725
transform 1 0 7636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_120
timestamp 1676037725
transform 1 0 12144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1676037725
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1676037725
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_168
timestamp 1676037725
transform 1 0 16560 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1676037725
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_204
timestamp 1676037725
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_232
timestamp 1676037725
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1676037725
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_276
timestamp 1676037725
transform 1 0 26496 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_284
timestamp 1676037725
transform 1 0 27232 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_296
timestamp 1676037725
transform 1 0 28336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_338
timestamp 1676037725
transform 1 0 32200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1676037725
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1676037725
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1676037725
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1676037725
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1676037725
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_100
timestamp 1676037725
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1676037725
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1676037725
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_236
timestamp 1676037725
transform 1 0 22816 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_248
timestamp 1676037725
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_260
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_266
timestamp 1676037725
transform 1 0 25576 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_319
timestamp 1676037725
transform 1 0 30452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1676037725
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1676037725
transform 1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1676037725
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_51
timestamp 1676037725
transform 1 0 5796 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_59
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_120
timestamp 1676037725
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1676037725
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_150
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_161
timestamp 1676037725
transform 1 0 15916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_176
timestamp 1676037725
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_186
timestamp 1676037725
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1676037725
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1676037725
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_261
timestamp 1676037725
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1676037725
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_326
timestamp 1676037725
transform 1 0 31096 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_338
timestamp 1676037725
transform 1 0 32200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1676037725
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1676037725
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1676037725
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1676037725
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_75
timestamp 1676037725
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_87
timestamp 1676037725
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1676037725
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_145
timestamp 1676037725
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_156
timestamp 1676037725
transform 1 0 15456 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1676037725
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_213
timestamp 1676037725
transform 1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_244
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1676037725
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1676037725
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1676037725
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1676037725
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1676037725
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1676037725
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_36
timestamp 1676037725
transform 1 0 4416 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1676037725
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1676037725
transform 1 0 6624 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_64
timestamp 1676037725
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1676037725
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1676037725
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_127
timestamp 1676037725
transform 1 0 12788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_158
timestamp 1676037725
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1676037725
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1676037725
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1676037725
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1676037725
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_261
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_269
timestamp 1676037725
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1676037725
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_287
timestamp 1676037725
transform 1 0 27508 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1676037725
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1676037725
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1676037725
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_332
timestamp 1676037725
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_344
timestamp 1676037725
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1676037725
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1676037725
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1676037725
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1676037725
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_136
timestamp 1676037725
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1676037725
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_202
timestamp 1676037725
transform 1 0 19688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_210
timestamp 1676037725
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_246
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1676037725
transform 1 0 24748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1676037725
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_290
timestamp 1676037725
transform 1 0 27784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1676037725
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_319
timestamp 1676037725
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1676037725
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1676037725
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_357
timestamp 1676037725
transform 1 0 33948 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_363
timestamp 1676037725
transform 1 0 34500 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_93
timestamp 1676037725
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_105
timestamp 1676037725
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1676037725
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_120
timestamp 1676037725
transform 1 0 12144 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_128
timestamp 1676037725
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1676037725
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_205
timestamp 1676037725
transform 1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1676037725
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1676037725
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_270
timestamp 1676037725
transform 1 0 25944 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_283
timestamp 1676037725
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_293
timestamp 1676037725
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1676037725
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1676037725
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_334
timestamp 1676037725
transform 1 0 31832 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_344
timestamp 1676037725
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1676037725
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_92
timestamp 1676037725
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1676037725
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_121
timestamp 1676037725
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_133
timestamp 1676037725
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_140
timestamp 1676037725
transform 1 0 13984 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1676037725
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1676037725
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_206
timestamp 1676037725
transform 1 0 20056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1676037725
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_236
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_248
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1676037725
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_288
timestamp 1676037725
transform 1 0 27600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_300
timestamp 1676037725
transform 1 0 28704 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_308
timestamp 1676037725
transform 1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1676037725
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_99
timestamp 1676037725
transform 1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_111
timestamp 1676037725
transform 1 0 11316 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_123
timestamp 1676037725
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1676037725
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_152
timestamp 1676037725
transform 1 0 15088 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_160
timestamp 1676037725
transform 1 0 15824 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1676037725
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1676037725
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1676037725
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1676037725
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_328
timestamp 1676037725
transform 1 0 31280 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_340
timestamp 1676037725
transform 1 0 32384 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_352
timestamp 1676037725
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_78
timestamp 1676037725
transform 1 0 8280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_89
timestamp 1676037725
transform 1 0 9292 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_96
timestamp 1676037725
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1676037725
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_143
timestamp 1676037725
transform 1 0 14260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1676037725
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1676037725
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1676037725
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1676037725
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1676037725
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_246
timestamp 1676037725
transform 1 0 23736 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1676037725
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_288
timestamp 1676037725
transform 1 0 27600 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_300
timestamp 1676037725
transform 1 0 28704 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_318
timestamp 1676037725
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1676037725
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_93
timestamp 1676037725
transform 1 0 9660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_105
timestamp 1676037725
transform 1 0 10764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1676037725
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1676037725
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1676037725
transform 1 0 15548 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_170
timestamp 1676037725
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_182
timestamp 1676037725
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_219
timestamp 1676037725
transform 1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_227
timestamp 1676037725
transform 1 0 21988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_271
timestamp 1676037725
transform 1 0 26036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_293
timestamp 1676037725
transform 1 0 28060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_299
timestamp 1676037725
transform 1 0 28612 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1676037725
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_92
timestamp 1676037725
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1676037725
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_136
timestamp 1676037725
transform 1 0 13616 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_144
timestamp 1676037725
transform 1 0 14352 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_151
timestamp 1676037725
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1676037725
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_177
timestamp 1676037725
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_214
timestamp 1676037725
transform 1 0 20792 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1676037725
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_248
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_267
timestamp 1676037725
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1676037725
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1676037725
transform 1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_105
timestamp 1676037725
transform 1 0 10764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_117
timestamp 1676037725
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_125
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 1676037725
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1676037725
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1676037725
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_223
timestamp 1676037725
transform 1 0 21620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_235
timestamp 1676037725
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1676037725
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_262
timestamp 1676037725
transform 1 0 25208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_274
timestamp 1676037725
transform 1 0 26312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_282
timestamp 1676037725
transform 1 0 27048 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_292
timestamp 1676037725
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1676037725
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_316
timestamp 1676037725
transform 1 0 30176 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1676037725
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_340
timestamp 1676037725
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_352
timestamp 1676037725
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_133
timestamp 1676037725
transform 1 0 13340 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_156
timestamp 1676037725
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_187
timestamp 1676037725
transform 1 0 18308 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1676037725
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1676037725
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_294
timestamp 1676037725
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_306
timestamp 1676037725
transform 1 0 29256 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_315
timestamp 1676037725
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1676037725
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1676037725
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1676037725
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_106
timestamp 1676037725
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_118
timestamp 1676037725
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1676037725
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_168
timestamp 1676037725
transform 1 0 16560 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_180
timestamp 1676037725
transform 1 0 17664 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1676037725
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_217
timestamp 1676037725
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1676037725
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_241
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_276
timestamp 1676037725
transform 1 0 26496 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_284
timestamp 1676037725
transform 1 0 27232 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1676037725
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1676037725
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1676037725
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_156
timestamp 1676037725
transform 1 0 15456 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_162
timestamp 1676037725
transform 1 0 16008 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1676037725
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_182
timestamp 1676037725
transform 1 0 17848 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_194
timestamp 1676037725
transform 1 0 18952 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1676037725
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_250
timestamp 1676037725
transform 1 0 24104 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1676037725
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1676037725
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1676037725
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1676037725
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_98
timestamp 1676037725
transform 1 0 10120 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_106
timestamp 1676037725
transform 1 0 10856 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_117
timestamp 1676037725
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_146
timestamp 1676037725
transform 1 0 14536 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_154
timestamp 1676037725
transform 1 0 15272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_162
timestamp 1676037725
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1676037725
transform 1 0 17664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1676037725
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_220
timestamp 1676037725
transform 1 0 21344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_226
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 1676037725
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1676037725
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_292
timestamp 1676037725
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_89
timestamp 1676037725
transform 1 0 9292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_97
timestamp 1676037725
transform 1 0 10028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_124
timestamp 1676037725
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1676037725
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_187
timestamp 1676037725
transform 1 0 18308 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_199
timestamp 1676037725
transform 1 0 19412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_211
timestamp 1676037725
transform 1 0 20516 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_230
timestamp 1676037725
transform 1 0 22264 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_241
timestamp 1676037725
transform 1 0 23276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_257
timestamp 1676037725
transform 1 0 24748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1676037725
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1676037725
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_313
timestamp 1676037725
transform 1 0 29900 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_320
timestamp 1676037725
transform 1 0 30544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1676037725
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_345
timestamp 1676037725
transform 1 0 32844 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_351
timestamp 1676037725
transform 1 0 33396 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_363
timestamp 1676037725
transform 1 0 34500 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_100
timestamp 1676037725
transform 1 0 10304 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_112
timestamp 1676037725
transform 1 0 11408 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_124
timestamp 1676037725
transform 1 0 12512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1676037725
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_159
timestamp 1676037725
transform 1 0 15732 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_172
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1676037725
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_216
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_228
timestamp 1676037725
transform 1 0 22080 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_232
timestamp 1676037725
transform 1 0 22448 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1676037725
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_29
timestamp 1676037725
transform 1 0 3772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_37
timestamp 1676037725
transform 1 0 4508 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1676037725
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_76
timestamp 1676037725
transform 1 0 8096 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_85
timestamp 1676037725
transform 1 0 8924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_97
timestamp 1676037725
transform 1 0 10028 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_103
timestamp 1676037725
transform 1 0 10580 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1676037725
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1676037725
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_147
timestamp 1676037725
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1676037725
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_175
timestamp 1676037725
transform 1 0 17204 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_187
timestamp 1676037725
transform 1 0 18308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_195
timestamp 1676037725
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_197
timestamp 1676037725
transform 1 0 19228 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1676037725
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1676037725
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1676037725
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_236
timestamp 1676037725
transform 1 0 22816 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_248
timestamp 1676037725
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_253
timestamp 1676037725
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_261
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_268
timestamp 1676037725
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_300
timestamp 1676037725
transform 1 0 28704 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1676037725
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_321
timestamp 1676037725
transform 1 0 30636 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_327
timestamp 1676037725
transform 1 0 31188 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1676037725
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_357
timestamp 1676037725
transform 1 0 33948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1676037725
transform 1 0 34408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1676037725
transform -1 0 4232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4416 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5980 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1676037725
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1676037725
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1676037725
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _0473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _0474_
timestamp 1676037725
transform 1 0 9568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0476_
timestamp 1676037725
transform 1 0 26036 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1676037725
transform -1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1676037725
transform -1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1676037725
transform 1 0 28704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0480_
timestamp 1676037725
transform -1 0 33396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0481_
timestamp 1676037725
transform -1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0482__1
timestamp 1676037725
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1676037725
transform -1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1676037725
transform -1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26128 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5336 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10304 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1676037725
transform -1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1676037725
transform 1 0 22080 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1676037725
transform -1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15824 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0503_
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15364 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1676037725
transform -1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0506_
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0507_
timestamp 1676037725
transform -1 0 6348 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0508_
timestamp 1676037725
transform 1 0 7360 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0509_
timestamp 1676037725
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0510_
timestamp 1676037725
transform -1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1676037725
transform 1 0 19780 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0512_
timestamp 1676037725
transform 1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0513_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6624 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0516_
timestamp 1676037725
transform -1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1676037725
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0520_
timestamp 1676037725
transform 1 0 12144 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0522_
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1676037725
transform -1 0 14812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0524_
timestamp 1676037725
transform 1 0 6624 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0527_
timestamp 1676037725
transform 1 0 26404 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_2  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0529_
timestamp 1676037725
transform 1 0 11684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0530_
timestamp 1676037725
transform 1 0 12880 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0532_
timestamp 1676037725
transform 1 0 2576 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp 1676037725
transform -1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3588 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0537_
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0538_
timestamp 1676037725
transform -1 0 4600 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0540_
timestamp 1676037725
transform -1 0 3404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0541_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1676037725
transform -1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0543_
timestamp 1676037725
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0546_
timestamp 1676037725
transform -1 0 15916 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0547_
timestamp 1676037725
transform -1 0 13248 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0548_
timestamp 1676037725
transform -1 0 14260 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0549_
timestamp 1676037725
transform -1 0 25484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27508 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0551_
timestamp 1676037725
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0552_
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27140 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1676037725
transform -1 0 28612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0555_
timestamp 1676037725
transform -1 0 27600 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1676037725
transform -1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26680 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0559_
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_2  _0560_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26312 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_4  _0562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26496 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28704 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0564_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0565_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _0566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27048 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _0567_
timestamp 1676037725
transform 1 0 24656 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1676037725
transform 1 0 24472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0569_
timestamp 1676037725
transform -1 0 25668 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0570_
timestamp 1676037725
transform -1 0 27968 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_8  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0573_
timestamp 1676037725
transform -1 0 27416 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0574_
timestamp 1676037725
transform 1 0 29624 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0575_
timestamp 1676037725
transform -1 0 28336 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_4  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_2  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28980 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_4  _0581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0582_
timestamp 1676037725
transform -1 0 22816 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0583_
timestamp 1676037725
transform -1 0 23276 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27324 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _0585_
timestamp 1676037725
transform -1 0 26036 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29164 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1676037725
transform -1 0 22448 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0589_
timestamp 1676037725
transform -1 0 19504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0590_
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1676037725
transform -1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0592_
timestamp 1676037725
transform 1 0 19780 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1676037725
transform -1 0 23736 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0594_
timestamp 1676037725
transform -1 0 24104 0 1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_2  _0595_
timestamp 1676037725
transform -1 0 21620 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _0596_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1676037725
transform 1 0 20608 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0598_
timestamp 1676037725
transform -1 0 21252 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1676037725
transform -1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23920 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0601_
timestamp 1676037725
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_1  _0603_
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1676037725
transform -1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _0607_
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20608 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1676037725
transform -1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0610_
timestamp 1676037725
transform -1 0 15824 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0611_
timestamp 1676037725
transform -1 0 14996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15180 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0614_
timestamp 1676037725
transform -1 0 19688 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _0615_
timestamp 1676037725
transform -1 0 13800 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _0616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0617_
timestamp 1676037725
transform -1 0 20424 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1676037725
transform -1 0 16376 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16560 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1676037725
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1676037725
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _0623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__a21boi_2  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16008 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0626_
timestamp 1676037725
transform -1 0 15548 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _0627_
timestamp 1676037725
transform -1 0 13432 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0628_
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0630_
timestamp 1676037725
transform -1 0 13800 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1676037725
transform -1 0 10304 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 1676037725
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13984 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _0634_
timestamp 1676037725
transform -1 0 15456 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1676037725
transform -1 0 10212 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0636_
timestamp 1676037725
transform 1 0 11684 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1676037725
transform -1 0 9568 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0639_
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1676037725
transform -1 0 16376 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0641_
timestamp 1676037725
transform -1 0 18308 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0643_
timestamp 1676037725
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _0644_
timestamp 1676037725
transform 1 0 9936 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12512 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp 1676037725
transform 1 0 9476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0649_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1676037725
transform -1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1676037725
transform 1 0 7728 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0652_
timestamp 1676037725
transform 1 0 12880 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0654_
timestamp 1676037725
transform -1 0 13708 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1676037725
transform -1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1676037725
transform -1 0 15916 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1676037725
transform -1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1676037725
transform -1 0 15640 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 1676037725
transform -1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1676037725
transform -1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0662_
timestamp 1676037725
transform 1 0 14720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0663_
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0664_
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1676037725
transform -1 0 8648 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0666_
timestamp 1676037725
transform 1 0 8924 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1676037725
transform 1 0 9292 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1676037725
transform -1 0 9292 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0671_
timestamp 1676037725
transform -1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1676037725
transform -1 0 9568 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0673_
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0674_
timestamp 1676037725
transform -1 0 16376 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0675_
timestamp 1676037725
transform -1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1676037725
transform -1 0 10028 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0678_
timestamp 1676037725
transform -1 0 16652 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0679_
timestamp 1676037725
transform -1 0 16376 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_4  _0680_
timestamp 1676037725
transform 1 0 17664 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0681_
timestamp 1676037725
transform -1 0 32568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1676037725
transform 1 0 31832 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1676037725
transform -1 0 32660 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1676037725
transform -1 0 29624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0688_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _0689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31924 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1676037725
transform -1 0 33212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0692_
timestamp 1676037725
transform -1 0 33120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1676037725
transform -1 0 31832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0694_
timestamp 1676037725
transform -1 0 32660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0695_
timestamp 1676037725
transform -1 0 31648 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0696_
timestamp 1676037725
transform -1 0 31740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0697_
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0698_
timestamp 1676037725
transform -1 0 31556 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32568 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0700_
timestamp 1676037725
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1676037725
transform -1 0 33396 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1676037725
transform -1 0 33672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0703_
timestamp 1676037725
transform -1 0 33212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1676037725
transform 1 0 33120 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0706_
timestamp 1676037725
transform -1 0 32200 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1676037725
transform 1 0 33580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0708_
timestamp 1676037725
transform 1 0 33488 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0709_
timestamp 1676037725
transform -1 0 30176 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ba_1  _0711_
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1676037725
transform -1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_4  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_1  _0715_
timestamp 1676037725
transform -1 0 28152 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 1676037725
transform -1 0 31188 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0719_
timestamp 1676037725
transform 1 0 28428 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1676037725
transform -1 0 27968 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0721_
timestamp 1676037725
transform -1 0 29348 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1676037725
transform -1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1676037725
transform 1 0 29716 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0725_
timestamp 1676037725
transform 1 0 30820 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1676037725
transform -1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1676037725
transform -1 0 27416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _0728_
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0729_
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0730_
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0731_
timestamp 1676037725
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0732_
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0733_
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0735_
timestamp 1676037725
transform 1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0736_
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0738_
timestamp 1676037725
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0739_
timestamp 1676037725
transform -1 0 17204 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0740_
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0741_
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1676037725
transform -1 0 22632 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1676037725
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0744_
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0745_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1676037725
transform 1 0 20516 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0747_
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1676037725
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1676037725
transform -1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0750_
timestamp 1676037725
transform 1 0 24656 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1676037725
transform 1 0 25852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0754_
timestamp 1676037725
transform -1 0 14812 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 1676037725
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0757_
timestamp 1676037725
transform -1 0 3496 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1676037725
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 1676037725
transform -1 0 12880 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0760_
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0761_
timestamp 1676037725
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1676037725
transform 1 0 12052 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0763_
timestamp 1676037725
transform -1 0 30360 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1676037725
transform -1 0 28428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0765_
timestamp 1676037725
transform -1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0767_
timestamp 1676037725
transform -1 0 28980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0768_
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0769_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1676037725
transform -1 0 25300 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0771_
timestamp 1676037725
transform 1 0 25024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1676037725
transform -1 0 28060 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0773_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0774_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0775_
timestamp 1676037725
transform 1 0 12236 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1676037725
transform -1 0 3496 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0777_
timestamp 1676037725
transform 1 0 2668 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0778_
timestamp 1676037725
transform -1 0 4416 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1676037725
transform -1 0 4416 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0780_
timestamp 1676037725
transform -1 0 15640 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0781_
timestamp 1676037725
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1676037725
transform -1 0 17572 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1676037725
transform -1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1676037725
transform -1 0 27784 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1676037725
transform -1 0 28980 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1676037725
transform 1 0 20424 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1676037725
transform -1 0 23000 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1676037725
transform 1 0 27232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0789_
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0790_
timestamp 1676037725
transform 1 0 27968 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0791_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0792_
timestamp 1676037725
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0793_
timestamp 1676037725
transform -1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1676037725
transform 1 0 15088 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0795_
timestamp 1676037725
transform -1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1676037725
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _0797_
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1676037725
transform -1 0 8648 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0799_
timestamp 1676037725
transform -1 0 8648 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _0800_
timestamp 1676037725
transform -1 0 9476 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1676037725
transform -1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0803_
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0806_
timestamp 1676037725
transform -1 0 27876 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0808_
timestamp 1676037725
transform -1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1676037725
transform 1 0 19412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0810_
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0812_
timestamp 1676037725
transform -1 0 21160 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0813_
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _0814_
timestamp 1676037725
transform -1 0 20976 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0816_
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1676037725
transform -1 0 11960 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1676037725
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1676037725
transform 1 0 10212 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 1676037725
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0823_
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0824_
timestamp 1676037725
transform -1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1676037725
transform 1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1676037725
transform 1 0 6348 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0827_
timestamp 1676037725
transform -1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1676037725
transform -1 0 7912 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0830_
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0831_
timestamp 1676037725
transform 1 0 4416 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0832_
timestamp 1676037725
transform -1 0 5796 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0833_
timestamp 1676037725
transform -1 0 4692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1676037725
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0835_
timestamp 1676037725
transform -1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _0836_
timestamp 1676037725
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1676037725
transform 1 0 3128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1676037725
transform -1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0839_
timestamp 1676037725
transform -1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1676037725
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0841_
timestamp 1676037725
transform -1 0 10764 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0842_
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1676037725
transform 1 0 7176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1676037725
transform -1 0 8648 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1676037725
transform -1 0 8556 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0847_
timestamp 1676037725
transform 1 0 6900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1676037725
transform 1 0 4140 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1676037725
transform 1 0 3128 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0850_
timestamp 1676037725
transform 1 0 5060 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1676037725
transform -1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0852_
timestamp 1676037725
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1676037725
transform 1 0 5060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0856_
timestamp 1676037725
transform 1 0 2944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1676037725
transform -1 0 5520 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0858_
timestamp 1676037725
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0862_
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0863_
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1676037725
transform 1 0 6992 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0865_
timestamp 1676037725
transform -1 0 8648 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0866_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0867_
timestamp 1676037725
transform -1 0 9752 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0868_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1676037725
transform -1 0 3496 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0870_
timestamp 1676037725
transform -1 0 3496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0871_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0872_
timestamp 1676037725
transform 1 0 29348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0873_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0874_
timestamp 1676037725
transform 1 0 23552 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0875_
timestamp 1676037725
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0877_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0878_
timestamp 1676037725
transform 1 0 28612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0879_
timestamp 1676037725
transform 1 0 20608 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0880_
timestamp 1676037725
transform 1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0881_
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0882_
timestamp 1676037725
transform -1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0883_
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0884_
timestamp 1676037725
transform -1 0 20976 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0885_
timestamp 1676037725
transform 1 0 14352 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0886_
timestamp 1676037725
transform -1 0 18952 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1676037725
transform -1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1676037725
transform 1 0 25484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0891_
timestamp 1676037725
transform 1 0 11960 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1676037725
transform 1 0 28336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1676037725
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0895_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1676037725
transform 1 0 23552 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1676037725
transform 1 0 17296 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1676037725
transform -1 0 28244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1676037725
transform 1 0 28704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1676037725
transform 1 0 30176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1676037725
transform -1 0 23000 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1676037725
transform 1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1676037725
transform -1 0 31648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0910_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1676037725
transform -1 0 31832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1676037725
transform -1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0913_
timestamp 1676037725
transform -1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1676037725
transform 1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1676037725
transform -1 0 18952 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1676037725
transform 1 0 20792 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1676037725
transform -1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1676037725
transform -1 0 25116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0923_
timestamp 1676037725
transform -1 0 26680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1676037725
transform 1 0 27140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1676037725
transform -1 0 19964 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0926_
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1676037725
transform 1 0 26128 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1676037725
transform -1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0931_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1676037725
transform -1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1676037725
transform -1 0 30176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1676037725
transform -1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1676037725
transform -1 0 31832 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1676037725
transform 1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1676037725
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0941_
timestamp 1676037725
transform 1 0 17664 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1676037725
transform -1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1676037725
transform 1 0 29808 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0946_
timestamp 1676037725
transform 1 0 32200 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1676037725
transform 1 0 30544 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1676037725
transform -1 0 21528 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0950_
timestamp 1676037725
transform 1 0 23276 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1676037725
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 1676037725
transform -1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1676037725
transform -1 0 25116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1676037725
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0956_
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0957_
timestamp 1676037725
transform -1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1676037725
transform -1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0959_
timestamp 1676037725
transform -1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0960_
timestamp 1676037725
transform 1 0 9292 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0961_
timestamp 1676037725
transform 1 0 12144 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0962_
timestamp 1676037725
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0963_
timestamp 1676037725
transform 1 0 2944 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0964_
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0965_
timestamp 1676037725
transform -1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0966_
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0967_
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1676037725
transform -1 0 14536 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0970_
timestamp 1676037725
transform 1 0 12696 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0971_
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1676037725
transform -1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0973_
timestamp 1676037725
transform -1 0 5704 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0974__2
timestamp 1676037725
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975__3
timestamp 1676037725
transform 1 0 15180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976__4
timestamp 1676037725
transform -1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977__5
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978__6
timestamp 1676037725
transform -1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979__7
timestamp 1676037725
transform -1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980__8
timestamp 1676037725
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1676037725
transform 1 0 27324 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1676037725
transform 1 0 27324 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1676037725
transform 1 0 24564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1676037725
transform -1 0 16376 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform -1 0 17020 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1676037725
transform -1 0 29256 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1676037725
transform 1 0 28336 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1676037725
transform 1 0 28612 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1676037725
transform 1 0 19504 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1676037725
transform 1 0 19872 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform -1 0 32844 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1676037725
transform 1 0 32292 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1676037725
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1676037725
transform 1 0 15272 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_4  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1009_
timestamp 1676037725
transform 1 0 1656 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1010_
timestamp 1676037725
transform -1 0 12052 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1011_
timestamp 1676037725
transform -1 0 12144 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1012_
timestamp 1676037725
transform -1 0 13616 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1013_
timestamp 1676037725
transform -1 0 13156 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1676037725
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 10764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1676037725
transform 1 0 7084 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1676037725
transform 1 0 9108 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1676037725
transform 1 0 6532 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1031_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1032_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1033_
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1034_
timestamp 1676037725
transform -1 0 9660 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  _1035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1036_
timestamp 1676037725
transform 1 0 6808 0 -1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _1039_
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1040_
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1676037725
transform -1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1676037725
transform 1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1676037725
transform 1 0 16652 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 17664 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1676037725
transform -1 0 21528 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform -1 0 26036 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 24288 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 26036 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform 1 0 26404 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform -1 0 25484 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1065_
timestamp 1676037725
transform -1 0 31464 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1676037725
transform 1 0 31832 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1069_
timestamp 1676037725
transform 1 0 23184 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1071_
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1072_
timestamp 1676037725
transform 1 0 23092 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1676037725
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1676037725
transform -1 0 18124 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1676037725
transform -1 0 18308 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1676037725
transform 1 0 17848 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1676037725
transform 1 0 29716 0 -1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1676037725
transform 1 0 29808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1676037725
transform 1 0 30084 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1080_
timestamp 1676037725
transform 1 0 30084 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1081_
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1676037725
transform -1 0 21252 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1676037725
transform -1 0 25116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform -1 0 25024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1676037725
transform -1 0 19688 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1676037725
transform 1 0 29992 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1676037725
transform 1 0 21620 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1676037725
transform -1 0 30636 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1676037725
transform 1 0 20148 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0460_
timestamp 1676037725
transform 1 0 20608 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1676037725
transform 1 0 15548 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1676037725
transform 1 0 31188 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1676037725
transform -1 0 33028 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1676037725
transform 1 0 20792 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1676037725
transform -1 0 17480 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1676037725
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1676037725
transform -1 0 22632 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1676037725
transform 1 0 23368 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1676037725
transform -1 0 22632 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1676037725
transform -1 0 14812 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1676037725
transform 1 0 28612 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0460_
timestamp 1676037725
transform -1 0 20056 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1676037725
transform 1 0 31188 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1676037725
transform -1 0 25208 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1676037725
transform -1 0 33028 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1676037725
transform 1 0 18216 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1676037725
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1676037725
transform -1 0 22632 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1676037725
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1676037725
transform -1 0 28612 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1676037725
transform 1 0 18216 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0460_
timestamp 1676037725
transform 1 0 20792 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform -1 0 20056 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 20792 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout29
timestamp 1676037725
transform -1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1676037725
transform -1 0 22816 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout35
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1676037725
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1676037725
transform 1 0 14996 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1676037725
transform 1 0 19688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout40
timestamp 1676037725
transform -1 0 17020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1676037725
transform 1 0 18400 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1676037725
transform -1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout44
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1676037725
transform -1 0 12788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1676037725
transform -1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1676037725
transform -1 0 29808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1676037725
transform 1 0 26128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1676037725
transform -1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1676037725
transform 1 0 26404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1676037725
transform 1 0 13248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout54
timestamp 1676037725
transform -1 0 4784 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout55
timestamp 1676037725
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 10672 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform -1 0 14628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform -1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1676037725
transform -1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform -1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform -1 0 25760 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform -1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform -1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform -1 0 34408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 4784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1676037725
transform -1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1676037725
transform -1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1676037725
transform -1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1676037725
transform 1 0 28336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1676037725
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1676037725
transform -1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_58
timestamp 1676037725
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_59
timestamp 1676037725
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_60
timestamp 1676037725
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_61
timestamp 1676037725
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_62
timestamp 1676037725
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_63
timestamp 1676037725
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_64
timestamp 1676037725
transform -1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_65
timestamp 1676037725
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_66
timestamp 1676037725
transform -1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_67
timestamp 1676037725
transform -1 0 34408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_68
timestamp 1676037725
transform -1 0 34408 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 1766 35200 1822 36000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 7654 35200 7710 36000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 10598 35200 10654 36000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 13542 35200 13598 36000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 16486 35200 16542 36000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 19430 35200 19486 36000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 22374 35200 22430 36000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 25318 35200 25374 36000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 28262 35200 28318 36000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 31206 35200 31262 36000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 34150 35200 34206 36000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 35200 17824 36000 17944 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 4710 35200 4766 36000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 5164 2128 5484 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 13605 2128 13925 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 22046 2128 22366 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 30487 2128 30807 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9384 2128 9704 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
