// This is the unpowered netlist.
module tholin_avalonsemi_5401 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [9:0] io_in;
 output [26:0] io_out;

 wire \CIRCUIT_1957.D0 ;
 wire \CIRCUIT_1957.D1 ;
 wire \CIRCUIT_1957.D2 ;
 wire \CIRCUIT_1957.D3 ;
 wire \CIRCUIT_1957.GATES_10.result ;
 wire \CIRCUIT_1957.GATES_27.result ;
 wire \CIRCUIT_1957.GATES_28.result ;
 wire \CIRCUIT_1957.GATES_30.result ;
 wire \CIRCUIT_1957.GATES_33.input2 ;
 wire \CIRCUIT_1957.GATES_35.result ;
 wire \CIRCUIT_1957.GATES_38.result ;
 wire \CIRCUIT_1957.GATES_39.result ;
 wire \CIRCUIT_1957.GATES_40.result ;
 wire \CIRCUIT_1957.GATES_41.result ;
 wire \CIRCUIT_1957.GATES_42.result ;
 wire \CIRCUIT_1957.GATES_53.result ;
 wire \CIRCUIT_1957.GATES_60.result ;
 wire \CIRCUIT_1957.GATES_9.result ;
 wire \CIRCUIT_1957.MEMORY_62.d ;
 wire \CIRCUIT_1957.MEMORY_62.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_63.d ;
 wire \CIRCUIT_1957.MEMORY_63.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_64.d ;
 wire \CIRCUIT_1957.MEMORY_64.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_65.d ;
 wire \CIRCUIT_1957.MEMORY_65.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_66.d ;
 wire \CIRCUIT_1957.MEMORY_66.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_67.d ;
 wire \CIRCUIT_1957.MEMORY_67.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_68.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_69.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_70.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_71.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_72.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_73.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_74.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_75.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_76.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_77.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_78.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_79.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_80.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_81.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_82.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_83.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_84.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_85.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_86.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_87.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_88.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.CLK1 ;
 wire \CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ;
 wire \CIRCUIT_1957.clock_gen_2_1.GATES_3.result ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A0 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A1 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A2 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A3 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A4 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A5 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A6 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A7 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B0 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B1 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B2 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B3 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A0 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A1 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A2 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A3 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B0 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B1 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B2 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B3 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire clknet_0_clk;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire net68;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net69;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire clknet_0__0460_;
 wire clknet_1_0__leaf__0460_;
 wire clknet_1_1__leaf__0460_;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ;

 sky130_fd_sc_hd__inv_2 _0465_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ));
 sky130_fd_sc_hd__inv_2 _0466_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ));
 sky130_fd_sc_hd__inv_6 _0467_ (.A(net53),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_4 _0468_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ));
 sky130_fd_sc_hd__inv_2 _0469_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _0470_ (.A(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _0471_ (.A(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _0472_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_4 _0473_ (.A(net33),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_4 _0474_ (.A(net28),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _0475_ (.A(net29),
    .Y(_0106_));
 sky130_fd_sc_hd__clkinv_4 _0476_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _0477_ (.A(net32),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .Y(_0110_));
 sky130_fd_sc_hd__clkinv_2 _0480_ (.A(net10),
    .Y(_0111_));
 sky130_fd_sc_hd__clkinv_2 _0481_ (.A(net9),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _0974__2 (.A(clknet_2_0__leaf_clk),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _0483_ (.A(\CIRCUIT_1957.GATES_33.input2 ),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ),
    .Y(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ));
 sky130_fd_sc_hd__or4b_4 _0486_ (.A(net22),
    .B(net21),
    .C(net25),
    .D_N(net24),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_1 _0487_ (.A(_0099_),
    .B(\CIRCUIT_1957.MEMORY_64.s_currentState ),
    .Y(_0116_));
 sky130_fd_sc_hd__and2_2 _0488_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(net53),
    .X(_0117_));
 sky130_fd_sc_hd__or4_1 _0489_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .C(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .D(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .X(_0118_));
 sky130_fd_sc_hd__o22a_1 _0490_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(_0116_),
    .B1(_0118_),
    .B2(net53),
    .X(_0119_));
 sky130_fd_sc_hd__nor3b_4 _0491_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(_0119_),
    .C_N(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0120_));
 sky130_fd_sc_hd__mux2_1 _0492_ (.A0(\CIRCUIT_1957.MEMORY_75.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_83.s_currentState ),
    .S(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0493_ (.A0(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .A1(_0121_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0494_ (.A0(_0122_),
    .A1(net20),
    .S(_0115_),
    .X(_0060_));
 sky130_fd_sc_hd__or3b_1 _0495_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .B(_0120_),
    .C_N(\CIRCUIT_1957.MEMORY_74.s_currentState ),
    .X(_0123_));
 sky130_fd_sc_hd__o21ai_1 _0496_ (.A1(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_82.s_currentState ),
    .B1(_0120_),
    .Y(_0124_));
 sky130_fd_sc_hd__a21oi_1 _0497_ (.A1(_0123_),
    .A2(_0124_),
    .B1(_0115_),
    .Y(_0125_));
 sky130_fd_sc_hd__a21o_1 _0498_ (.A1(net19),
    .A2(_0115_),
    .B1(_0125_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0499_ (.A0(\CIRCUIT_1957.MEMORY_73.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_81.s_currentState ),
    .S(_0120_),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_1 _0500_ (.A(\CIRCUIT_1957.MEMORY_75.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_74.s_currentState ),
    .Y(_0127_));
 sky130_fd_sc_hd__or4bb_4 _0501_ (.A(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .B(_0127_),
    .C_N(\CIRCUIT_1957.MEMORY_72.s_currentState ),
    .D_N(\CIRCUIT_1957.MEMORY_73.s_currentState ),
    .X(_0128_));
 sky130_fd_sc_hd__nand2_4 _0502_ (.A(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_4 _0503_ (.A(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .Y(_0130_));
 sky130_fd_sc_hd__nor2_2 _0504_ (.A(_0129_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2_2 _0506_ (.A(_0128_),
    .B(_0131_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_1 _0507_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0134_));
 sky130_fd_sc_hd__or3b_1 _0508_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0099_),
    .C_N(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2_1 _0509_ (.A(net42),
    .B(net44),
    .Y(_0136_));
 sky130_fd_sc_hd__mux2_1 _0510_ (.A0(_0126_),
    .A1(_0136_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0511_ (.A0(_0137_),
    .A1(net18),
    .S(_0115_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0512_ (.A0(\CIRCUIT_1957.MEMORY_72.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_80.s_currentState ),
    .S(_0120_),
    .X(_0138_));
 sky130_fd_sc_hd__nand2_1 _0513_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__o21a_1 _0515_ (.A1(_0134_),
    .A2(_0140_),
    .B1(_0117_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0516_ (.A0(_0138_),
    .A1(_0141_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0517_ (.A0(_0142_),
    .A1(net17),
    .S(_0115_),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_2 _0518_ (.A0(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_87.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_79.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0120_),
    .X(net27));
 sky130_fd_sc_hd__mux2_1 _0519_ (.A0(net27),
    .A1(net16),
    .S(_0115_),
    .X(_0056_));
 sky130_fd_sc_hd__mux4_2 _0520_ (.A0(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_86.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_78.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0120_),
    .X(net26));
 sky130_fd_sc_hd__mux2_1 _0521_ (.A0(net26),
    .A1(net15),
    .S(_0115_),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_2 _0522_ (.A0(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_85.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_77.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0120_),
    .X(net23));
 sky130_fd_sc_hd__mux2_1 _0523_ (.A0(net23),
    .A1(net14),
    .S(_0115_),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_2 _0524_ (.A0(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_84.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_76.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0120_),
    .X(net12));
 sky130_fd_sc_hd__mux2_1 _0525_ (.A0(net12),
    .A1(net13),
    .S(_0115_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_2 _0526_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0002_));
 sky130_fd_sc_hd__or4b_4 _0527_ (.A(net22),
    .B(net25),
    .C(net24),
    .D_N(net21),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_2 _0528_ (.A0(net5),
    .A1(net1),
    .S(_0143_),
    .X(\CIRCUIT_1957.D0 ));
 sky130_fd_sc_hd__mux2_2 _0529_ (.A0(net6),
    .A1(net2),
    .S(_0143_),
    .X(\CIRCUIT_1957.D1 ));
 sky130_fd_sc_hd__mux2_2 _0530_ (.A0(net7),
    .A1(net3),
    .S(_0143_),
    .X(\CIRCUIT_1957.D2 ));
 sky130_fd_sc_hd__mux2_4 _0531_ (.A0(net8),
    .A1(net4),
    .S(_0143_),
    .X(\CIRCUIT_1957.D3 ));
 sky130_fd_sc_hd__nand2_2 _0532_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(_0144_),
    .Y(\CIRCUIT_1957.clock_gen_2_1.CLK1 ));
 sky130_fd_sc_hd__and3b_2 _0534_ (.A_N(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .C(_0117_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _0535_ (.A(_0144_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__a31o_1 _0536_ (.A1(_0113_),
    .A2(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .A3(_0146_),
    .B1(net54),
    .X(_0147_));
 sky130_fd_sc_hd__a21o_1 _0537_ (.A1(\CIRCUIT_1957.GATES_33.input2 ),
    .A2(_0146_),
    .B1(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .X(_0148_));
 sky130_fd_sc_hd__a21o_1 _0538_ (.A1(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ),
    .A2(_0148_),
    .B1(_0147_),
    .X(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(_0114_),
    .A1(\CIRCUIT_1957.GATES_33.input2 ),
    .S(_0146_),
    .X(_0149_));
 sky130_fd_sc_hd__and3b_2 _0540_ (.A_N(net54),
    .B(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ),
    .C(_0149_),
    .X(\CIRCUIT_1957.GATES_33.input2 ));
 sky130_fd_sc_hd__a41o_1 _0541_ (.A1(_0113_),
    .A2(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ),
    .A3(_0144_),
    .A4(_0145_),
    .B1(_0147_),
    .X(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ));
 sky130_fd_sc_hd__nand2_1 _0542_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _0543_ (.A(_0145_),
    .B(_0150_),
    .Y(\CIRCUIT_1957.GATES_53.result ));
 sky130_fd_sc_hd__or4_4 _0544_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(net53),
    .C(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .D(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _0545_ (.A(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__nor2_2 _0546_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .Y(_0153_));
 sky130_fd_sc_hd__and2_2 _0547_ (.A(net31),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__nand2_2 _0548_ (.A(net31),
    .B(_0153_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_2 _0549_ (.A(net28),
    .B(net30),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2b_1 _0550_ (.A_N(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .B(net32),
    .Y(_0157_));
 sky130_fd_sc_hd__o21a_1 _0551_ (.A1(_0104_),
    .A2(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a31o_1 _0552_ (.A1(net33),
    .A2(_0156_),
    .A3(_0157_),
    .B1(_0109_),
    .X(_0159_));
 sky130_fd_sc_hd__a211o_1 _0553_ (.A1(net33),
    .A2(_0156_),
    .B1(_0109_),
    .C1(net31),
    .X(_0160_));
 sky130_fd_sc_hd__nor2_1 _0554_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .Y(_0161_));
 sky130_fd_sc_hd__nand2_2 _0555_ (.A(_0160_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__nor2_1 _0556_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .B(net32),
    .Y(_0163_));
 sky130_fd_sc_hd__and2b_1 _0557_ (.A_N(_0163_),
    .B(_0156_),
    .X(_0164_));
 sky130_fd_sc_hd__and3b_1 _0558_ (.A_N(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .B(net31),
    .C(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_2 _0559_ (.A(net32),
    .B(_0159_),
    .Y(_0166_));
 sky130_fd_sc_hd__o311a_2 _0560_ (.A1(net28),
    .A2(_0163_),
    .A3(_0165_),
    .B1(_0106_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .X(_0167_));
 sky130_fd_sc_hd__a211oi_4 _0561_ (.A1(net30),
    .A2(_0107_),
    .B1(_0167_),
    .C1(net28),
    .Y(_0168_));
 sky130_fd_sc_hd__a32o_4 _0562_ (.A1(_0162_),
    .A2(_0166_),
    .A3(_0168_),
    .B1(_0167_),
    .B2(_0105_),
    .X(_0169_));
 sky130_fd_sc_hd__and3_1 _0563_ (.A(net33),
    .B(_0110_),
    .C(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__a21oi_2 _0564_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .A2(_0169_),
    .B1(_0110_),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_2 _0565_ (.A(_0170_),
    .B(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__a311oi_4 _0566_ (.A1(_0162_),
    .A2(_0166_),
    .A3(_0168_),
    .B1(_0164_),
    .C1(_0107_),
    .Y(_0173_));
 sky130_fd_sc_hd__and2_2 _0567_ (.A(_0105_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _0568_ (.A(_0105_),
    .B(_0173_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_2 _0569_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .B(_0107_),
    .Y(_0176_));
 sky130_fd_sc_hd__a21o_1 _0570_ (.A1(_0160_),
    .A2(_0166_),
    .B1(_0161_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_8 _0571_ (.A0(_0159_),
    .A1(_0177_),
    .S(_0169_),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_4 _0572_ (.A(net30),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__nor2_1 _0573_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .Y(_0180_));
 sky130_fd_sc_hd__nor2_2 _0574_ (.A(net32),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__and2_2 _0575_ (.A(net32),
    .B(_0180_),
    .X(_0182_));
 sky130_fd_sc_hd__o21ba_1 _0576_ (.A1(_0170_),
    .A2(_0171_),
    .B1_N(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__o2bb2a_2 _0577_ (.A1_N(net30),
    .A2_N(_0178_),
    .B1(_0181_),
    .B2(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__o31ai_4 _0578_ (.A1(_0174_),
    .A2(_0179_),
    .A3(_0184_),
    .B1(_0176_),
    .Y(_0185_));
 sky130_fd_sc_hd__o31a_2 _0579_ (.A1(_0181_),
    .A2(_0182_),
    .A3(_0185_),
    .B1(_0172_),
    .X(_0186_));
 sky130_fd_sc_hd__nor4_4 _0580_ (.A(_0172_),
    .B(_0181_),
    .C(_0182_),
    .D(_0185_),
    .Y(_0187_));
 sky130_fd_sc_hd__o311a_4 _0581_ (.A1(_0174_),
    .A2(_0179_),
    .A3(_0184_),
    .B1(_0176_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .X(_0188_));
 sky130_fd_sc_hd__and2b_1 _0582_ (.A_N(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .B(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__nor2_2 _0583_ (.A(_0186_),
    .B(_0187_),
    .Y(_0190_));
 sky130_fd_sc_hd__or3_4 _0584_ (.A(_0181_),
    .B(_0183_),
    .C(_0185_),
    .X(_0191_));
 sky130_fd_sc_hd__o311a_2 _0585_ (.A1(_0174_),
    .A2(_0179_),
    .A3(_0184_),
    .B1(_0176_),
    .C1(net30),
    .X(_0192_));
 sky130_fd_sc_hd__xor2_4 _0586_ (.A(_0178_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__xnor2_4 _0587_ (.A(_0191_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_1 _0589_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .Y(_0196_));
 sky130_fd_sc_hd__nand2_2 _0590_ (.A(net32),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_2 _0592_ (.A(net31),
    .B(_0196_),
    .Y(_0199_));
 sky130_fd_sc_hd__and2b_1 _0593_ (.A_N(_0188_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .X(_0200_));
 sky130_fd_sc_hd__xor2_4 _0594_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .B(_0188_),
    .X(_0201_));
 sky130_fd_sc_hd__a21oi_2 _0595_ (.A1(_0197_),
    .A2(_0201_),
    .B1(_0199_),
    .Y(_0202_));
 sky130_fd_sc_hd__o311a_2 _0596_ (.A1(_0189_),
    .A2(_0199_),
    .A3(_0200_),
    .B1(_0197_),
    .C1(_0106_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _0597_ (.A(net30),
    .B(_0202_),
    .X(_0204_));
 sky130_fd_sc_hd__a211o_1 _0598_ (.A1(_0197_),
    .A2(_0201_),
    .B1(_0199_),
    .C1(_0106_),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _0599_ (.A1(_0190_),
    .A2(_0205_),
    .B1(_0203_),
    .Y(_0206_));
 sky130_fd_sc_hd__or3_1 _0600_ (.A(net30),
    .B(_0186_),
    .C(_0187_),
    .X(_0207_));
 sky130_fd_sc_hd__o21a_1 _0601_ (.A1(_0186_),
    .A2(_0187_),
    .B1(net30),
    .X(_0208_));
 sky130_fd_sc_hd__a221o_4 _0602_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .A2(_0194_),
    .B1(_0202_),
    .B2(_0207_),
    .C1(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__or3b_1 _0603_ (.A(_0179_),
    .B(_0184_),
    .C_N(_0173_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(_0105_),
    .A1(_0175_),
    .S(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__o21a_4 _0605_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .A2(_0194_),
    .B1(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _0606_ (.A(_0209_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__a211oi_4 _0607_ (.A1(_0209_),
    .A2(_0212_),
    .B1(_0203_),
    .C1(_0204_),
    .Y(_0214_));
 sky130_fd_sc_hd__xnor2_2 _0608_ (.A(_0190_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _0609_ (.A(net28),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor2_2 _0610_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .Y(_0217_));
 sky130_fd_sc_hd__and2_2 _0611_ (.A(net31),
    .B(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__or2_4 _0612_ (.A(net31),
    .B(_0217_),
    .X(_0219_));
 sky130_fd_sc_hd__a21oi_4 _0613_ (.A1(_0209_),
    .A2(_0212_),
    .B1(_0104_),
    .Y(_0220_));
 sky130_fd_sc_hd__xnor2_4 _0614_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__o21ai_1 _0615_ (.A1(_0218_),
    .A2(_0221_),
    .B1(_0219_),
    .Y(_0222_));
 sky130_fd_sc_hd__a211o_2 _0616_ (.A1(_0209_),
    .A2(_0212_),
    .B1(_0198_),
    .C1(_0199_),
    .X(_0223_));
 sky130_fd_sc_hd__xor2_4 _0617_ (.A(_0201_),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _0618_ (.A(net29),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__o221ai_4 _0619_ (.A1(_0218_),
    .A2(_0221_),
    .B1(_0224_),
    .B2(net29),
    .C1(_0219_),
    .Y(_0226_));
 sky130_fd_sc_hd__xnor2_1 _0620_ (.A(_0105_),
    .B(_0206_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _0621_ (.A(_0195_),
    .B(_0211_),
    .Y(_0228_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(_0195_),
    .A1(_0228_),
    .S(_0227_),
    .X(_0229_));
 sky130_fd_sc_hd__o21bai_1 _0623_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .A2(_0215_),
    .B1_N(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a31o_4 _0624_ (.A1(_0216_),
    .A2(_0225_),
    .A3(_0226_),
    .B1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__a21boi_2 _0625_ (.A1(net33),
    .A2(_0231_),
    .B1_N(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .Y(_0232_));
 sky130_fd_sc_hd__a21oi_4 _0626_ (.A1(_0217_),
    .A2(_0231_),
    .B1(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__or2_4 _0627_ (.A(net31),
    .B(_0153_),
    .X(_0234_));
 sky130_fd_sc_hd__xnor2_1 _0628_ (.A(net29),
    .B(_0222_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(_0231_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__xnor2_2 _0630_ (.A(_0224_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _0632_ (.A(net28),
    .B(_0237_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3b_4 _0633_ (.A_N(_0218_),
    .B(_0219_),
    .C(_0231_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_4 _0634_ (.A(_0221_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _0635_ (.A(net29),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__o221ai_4 _0636_ (.A1(_0154_),
    .A2(_0233_),
    .B1(_0241_),
    .B2(net29),
    .C1(_0234_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _0637_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__and3_1 _0638_ (.A(_0105_),
    .B(_0225_),
    .C(_0226_),
    .X(_0245_));
 sky130_fd_sc_hd__a21oi_1 _0639_ (.A1(_0225_),
    .A2(_0226_),
    .B1(_0105_),
    .Y(_0246_));
 sky130_fd_sc_hd__nor2_1 _0640_ (.A(_0245_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _0641_ (.A(_0215_),
    .B(_0229_),
    .Y(_0248_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(_0215_),
    .A1(_0248_),
    .S(_0247_),
    .X(_0249_));
 sky130_fd_sc_hd__o21ai_1 _0643_ (.A1(net28),
    .A2(_0237_),
    .B1(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__a31o_4 _0644_ (.A1(_0239_),
    .A2(_0242_),
    .A3(_0243_),
    .B1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__o211ai_4 _0645_ (.A1(_0154_),
    .A2(_0233_),
    .B1(_0234_),
    .C1(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21o_1 _0646_ (.A1(net29),
    .A2(_0251_),
    .B1(_0241_),
    .X(_0253_));
 sky130_fd_sc_hd__nand3_1 _0647_ (.A(net29),
    .B(_0241_),
    .C(_0251_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand3_2 _0648_ (.A(_0252_),
    .B(_0253_),
    .C(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21o_1 _0649_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0252_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _0650_ (.A(_0255_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__a21o_1 _0651_ (.A1(_0255_),
    .A2(_0256_),
    .B1(_0105_),
    .X(_0258_));
 sky130_fd_sc_hd__a31o_1 _0652_ (.A1(_0155_),
    .A2(_0234_),
    .A3(_0251_),
    .B1(_0233_),
    .X(_0259_));
 sky130_fd_sc_hd__nand4_4 _0653_ (.A(_0155_),
    .B(_0233_),
    .C(_0234_),
    .D(_0251_),
    .Y(_0260_));
 sky130_fd_sc_hd__and3_1 _0654_ (.A(net29),
    .B(_0259_),
    .C(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _0655_ (.A(_0104_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .Y(_0262_));
 sky130_fd_sc_hd__and2_1 _0656_ (.A(net31),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__inv_2 _0657_ (.A(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__or2_1 _0658_ (.A(net31),
    .B(_0262_),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _0659_ (.A(net33),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .C(_0251_),
    .X(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0660_ (.A1(net33),
    .A2(_0251_),
    .B1(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_1 _0661_ (.A(_0266_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__o31a_2 _0662_ (.A1(_0263_),
    .A2(_0266_),
    .A3(_0267_),
    .B1(_0265_),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_1 _0663_ (.A1(_0259_),
    .A2(_0260_),
    .B1(net29),
    .X(_0270_));
 sky130_fd_sc_hd__a21oi_2 _0664_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0261_),
    .Y(_0271_));
 sky130_fd_sc_hd__nor2_1 _0665_ (.A(_0238_),
    .B(_0249_),
    .Y(_0272_));
 sky130_fd_sc_hd__xnor2_1 _0666_ (.A(_0105_),
    .B(_0244_),
    .Y(_0273_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(_0238_),
    .A1(_0272_),
    .S(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__a31o_1 _0668_ (.A1(_0105_),
    .A2(_0255_),
    .A3(_0256_),
    .B1(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_4 _0669_ (.A1(_0258_),
    .A2(_0271_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__and2b_1 _0670_ (.A_N(_0271_),
    .B(_0275_),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _0671_ (.A1(net28),
    .A2(_0276_),
    .B1(_0257_),
    .Y(_0278_));
 sky130_fd_sc_hd__a31o_1 _0672_ (.A1(net28),
    .A2(_0257_),
    .A3(_0274_),
    .B1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__or2_4 _0673_ (.A(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .X(_0280_));
 sky130_fd_sc_hd__or2_4 _0674_ (.A(_0129_),
    .B(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _0675_ (.A1(_0277_),
    .A2(_0279_),
    .B1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__o21a_1 _0676_ (.A1(_0277_),
    .A2(_0279_),
    .B1(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2b_4 _0677_ (.A_N(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .Y(_0284_));
 sky130_fd_sc_hd__nor2_4 _0678_ (.A(_0129_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2b_4 _0679_ (.A_N(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .Y(_0286_));
 sky130_fd_sc_hd__or2_4 _0680_ (.A(_0130_),
    .B(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_2 _0681_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .Y(_0288_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0289_));
 sky130_fd_sc_hd__and2_1 _0683_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0290_));
 sky130_fd_sc_hd__and3_1 _0684_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .C(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__and4_2 _0685_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .C(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .D(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__a31o_2 _0687_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A3(_0290_),
    .B1(_0292_),
    .X(_0294_));
 sky130_fd_sc_hd__a21oi_2 _0688_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .A2(_0294_),
    .B1(_0291_),
    .Y(_0295_));
 sky130_fd_sc_hd__a22oi_2 _0689_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .Y(_0296_));
 sky130_fd_sc_hd__and4_1 _0690_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .C(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .D(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .X(_0297_));
 sky130_fd_sc_hd__nor2_1 _0691_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or3_4 _0692_ (.A(_0295_),
    .B(_0296_),
    .C(_0297_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .Y(_0300_));
 sky130_fd_sc_hd__a21oi_2 _0694_ (.A1(_0288_),
    .A2(_0299_),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21oi_2 _0695_ (.A1(_0299_),
    .A2(_0300_),
    .B1(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2b_1 _0696_ (.A_N(_0298_),
    .B(_0295_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _0697_ (.A(_0299_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_2 _0698_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0305_));
 sky130_fd_sc_hd__xor2_1 _0699_ (.A(_0288_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a21oi_1 _0700_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B1(_0290_),
    .Y(_0307_));
 sky130_fd_sc_hd__nor2_1 _0701_ (.A(_0291_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__and2_1 _0702_ (.A(_0294_),
    .B(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o21a_1 _0703_ (.A1(_0289_),
    .A2(_0309_),
    .B1(_0295_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _0704_ (.A(_0306_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a2bb2o_2 _0705_ (.A1_N(_0288_),
    .A2_N(_0305_),
    .B1(_0306_),
    .B2(_0310_),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_2 _0706_ (.A(_0304_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nor2_1 _0707_ (.A(_0306_),
    .B(_0310_),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_4 _0708_ (.A(_0311_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_2 _0709_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .Y(_0316_));
 sky130_fd_sc_hd__a22oi_4 _0710_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0317_));
 sky130_fd_sc_hd__o21ba_1 _0711_ (.A1(_0305_),
    .A2(_0316_),
    .B1_N(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_1 _0712_ (.A(_0294_),
    .B(_0308_),
    .Y(_0319_));
 sky130_fd_sc_hd__or2_2 _0713_ (.A(_0309_),
    .B(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__o22a_4 _0714_ (.A1(_0305_),
    .A2(_0316_),
    .B1(_0317_),
    .B2(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__xor2_1 _0715_ (.A(_0318_),
    .B(_0320_),
    .X(_0322_));
 sky130_fd_sc_hd__a22oi_1 _0716_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_1 _0717_ (.A(_0290_),
    .B(_0292_),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_1 _0718_ (.A(_0294_),
    .B(_0323_),
    .X(_0325_));
 sky130_fd_sc_hd__a21o_1 _0719_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0316_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_4 _0720_ (.A(_0322_),
    .B(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_4 _0721_ (.A(_0315_),
    .B(_0321_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _0722_ (.A(_0327_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__o21bai_2 _0723_ (.A1(_0315_),
    .A2(_0321_),
    .B1_N(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__and2_1 _0724_ (.A(_0313_),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__a31o_1 _0725_ (.A1(_0299_),
    .A2(_0303_),
    .A3(_0312_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a21oi_1 _0726_ (.A1(_0302_),
    .A2(_0332_),
    .B1(_0301_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _0727_ (.A(_0322_),
    .B(_0326_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2b_4 _0728_ (.A_N(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_4 _0729_ (.A(_0286_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2b_4 _0730_ (.A_N(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .Y(_0337_));
 sky130_fd_sc_hd__nor2_4 _0731_ (.A(_0284_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__or2_4 _0732_ (.A(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .X(_0339_));
 sky130_fd_sc_hd__nor2_4 _0733_ (.A(_0130_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__a22o_1 _0734_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ),
    .A2(_0338_),
    .B1(_0340_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_4 _0735_ (.A(_0280_),
    .B(_0339_),
    .Y(_0342_));
 sky130_fd_sc_hd__nor2_2 _0736_ (.A(_0284_),
    .B(_0339_),
    .Y(_0343_));
 sky130_fd_sc_hd__a221o_1 _0737_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ),
    .A2(_0342_),
    .B1(_0343_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ),
    .C1(_0341_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_4 _0738_ (.A(_0280_),
    .B(_0337_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_2 _0739_ (.A(_0335_),
    .B(_0339_),
    .Y(_0346_));
 sky130_fd_sc_hd__nor2_4 _0740_ (.A(_0130_),
    .B(_0337_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_2 _0741_ (.A(_0335_),
    .B(_0337_),
    .Y(_0348_));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ),
    .A2(_0347_),
    .B1(_0348_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ),
    .X(_0349_));
 sky130_fd_sc_hd__a221o_1 _0743_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ),
    .A2(_0345_),
    .B1(_0346_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ),
    .C1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__nor2_2 _0744_ (.A(_0284_),
    .B(_0286_),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_4 _0745_ (.A(_0280_),
    .B(_0286_),
    .Y(_0352_));
 sky130_fd_sc_hd__a22o_1 _0746_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ),
    .A2(_0351_),
    .B1(_0352_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ),
    .X(_0353_));
 sky130_fd_sc_hd__or2_4 _0747_ (.A(_0129_),
    .B(_0335_),
    .X(_0354_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _0749_ (.A(net33),
    .B(_0107_),
    .Y(_0356_));
 sky130_fd_sc_hd__a41o_1 _0750_ (.A1(_0108_),
    .A2(_0156_),
    .A3(_0355_),
    .A4(_0356_),
    .B1(_0353_),
    .X(_0357_));
 sky130_fd_sc_hd__or3_1 _0751_ (.A(_0344_),
    .B(_0350_),
    .C(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__a31o_1 _0752_ (.A1(_0327_),
    .A2(_0334_),
    .A3(_0336_),
    .B1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__a2bb2o_1 _0753_ (.A1_N(_0287_),
    .A2_N(_0333_),
    .B1(_0213_),
    .B2(_0285_),
    .X(_0360_));
 sky130_fd_sc_hd__or3_1 _0754_ (.A(_0283_),
    .B(_0359_),
    .C(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_4 _0755_ (.A1(_0128_),
    .A2(\CIRCUIT_1957.D3 ),
    .B1(_0361_),
    .B2(net43),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_1 _0756_ (.A(_0099_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__xnor2_2 _0757_ (.A(_0099_),
    .B(_0362_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0152_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__xnor2_1 _0759_ (.A(_0106_),
    .B(_0269_),
    .Y(_0366_));
 sky130_fd_sc_hd__and4_1 _0760_ (.A(_0259_),
    .B(_0260_),
    .C(_0276_),
    .D(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__a22oi_1 _0761_ (.A1(_0259_),
    .A2(_0260_),
    .B1(_0276_),
    .B2(_0366_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21ba_1 _0762_ (.A1(_0367_),
    .A2(_0368_),
    .B1_N(_0281_),
    .X(_0369_));
 sky130_fd_sc_hd__xnor2_1 _0763_ (.A(_0302_),
    .B(_0332_),
    .Y(_0370_));
 sky130_fd_sc_hd__nor2_1 _0764_ (.A(_0287_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand3_1 _0765_ (.A(_0316_),
    .B(_0324_),
    .C(_0325_),
    .Y(_0372_));
 sky130_fd_sc_hd__a22o_1 _0766_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ),
    .A2(_0338_),
    .B1(_0342_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ),
    .X(_0373_));
 sky130_fd_sc_hd__a221o_1 _0767_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ),
    .A2(_0340_),
    .B1(_0343_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ),
    .C1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _0768_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ),
    .A2(_0345_),
    .B1(_0346_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ),
    .X(_0375_));
 sky130_fd_sc_hd__a221o_1 _0769_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ),
    .A2(_0351_),
    .B1(_0352_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ),
    .C1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a31o_1 _0770_ (.A1(_0156_),
    .A2(_0158_),
    .A3(_0355_),
    .B1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__a221o_1 _0771_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ),
    .A2(_0347_),
    .B1(_0348_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ),
    .C1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__a31o_1 _0772_ (.A1(_0326_),
    .A2(_0336_),
    .A3(_0372_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__or3_2 _0773_ (.A(_0371_),
    .B(_0374_),
    .C(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__a211o_1 _0774_ (.A1(_0231_),
    .A2(_0285_),
    .B1(_0369_),
    .C1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__a22o_4 _0775_ (.A1(_0128_),
    .A2(\CIRCUIT_1957.D2 ),
    .B1(_0381_),
    .B2(net43),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__xnor2_4 _0777_ (.A(_0099_),
    .B(_0382_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_2 _0778_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .B(_0151_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _0779_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .B(_0151_),
    .C(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__a31o_1 _0780_ (.A1(_0264_),
    .A2(_0265_),
    .A3(_0276_),
    .B1(_0268_),
    .X(_0387_));
 sky130_fd_sc_hd__a41o_1 _0781_ (.A1(_0264_),
    .A2(_0265_),
    .A3(_0268_),
    .A4(_0276_),
    .B1(_0281_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _0782_ (.A(_0262_),
    .B(_0276_),
    .Y(_0389_));
 sky130_fd_sc_hd__and2b_1 _0783_ (.A_N(_0388_),
    .B(_0387_),
    .X(_0390_));
 sky130_fd_sc_hd__xnor2_1 _0784_ (.A(_0313_),
    .B(_0330_),
    .Y(_0391_));
 sky130_fd_sc_hd__a22o_1 _0785_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .X(_0392_));
 sky130_fd_sc_hd__a22o_1 _0786_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ),
    .A2(_0345_),
    .B1(_0346_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ),
    .A2(_0342_),
    .B1(_0348_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ),
    .X(_0394_));
 sky130_fd_sc_hd__a221o_1 _0788_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ),
    .A2(_0340_),
    .B1(_0347_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ),
    .C1(_0393_),
    .X(_0395_));
 sky130_fd_sc_hd__a221o_1 _0789_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ),
    .A2(_0343_),
    .B1(_0352_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ),
    .C1(_0394_),
    .X(_0396_));
 sky130_fd_sc_hd__a31o_1 _0790_ (.A1(_0293_),
    .A2(_0336_),
    .A3(_0392_),
    .B1(_0395_),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _0791_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ),
    .A2(_0338_),
    .B1(_0351_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ),
    .C1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__a2bb2o_1 _0792_ (.A1_N(_0287_),
    .A2_N(_0391_),
    .B1(_0355_),
    .B2(_0169_),
    .X(_0399_));
 sky130_fd_sc_hd__or3_1 _0793_ (.A(_0396_),
    .B(_0398_),
    .C(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__a21o_1 _0794_ (.A1(_0251_),
    .A2(_0285_),
    .B1(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__o21ai_1 _0795_ (.A1(_0390_),
    .A2(_0401_),
    .B1(net43),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _0796_ (.A(_0128_),
    .B(\CIRCUIT_1957.D1 ),
    .Y(_0403_));
 sky130_fd_sc_hd__o311a_4 _0797_ (.A1(_0111_),
    .A2(_0128_),
    .A3(_0132_),
    .B1(_0402_),
    .C1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__xnor2_4 _0799_ (.A(net53),
    .B(_0404_),
    .Y(_0406_));
 sky130_fd_sc_hd__and2_2 _0800_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .B(_0151_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__a21bo_1 _0802_ (.A1(net33),
    .A2(_0276_),
    .B1_N(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .X(_0409_));
 sky130_fd_sc_hd__a21oi_2 _0803_ (.A1(_0389_),
    .A2(_0409_),
    .B1(_0281_),
    .Y(_0410_));
 sky130_fd_sc_hd__nor2_1 _0804_ (.A(_0185_),
    .B(_0354_),
    .Y(_0411_));
 sky130_fd_sc_hd__or2_2 _0805_ (.A(_0287_),
    .B(_0329_),
    .X(_0412_));
 sky130_fd_sc_hd__a21oi_4 _0806_ (.A1(_0327_),
    .A2(_0328_),
    .B1(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__a32o_1 _0807_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A3(_0336_),
    .B1(_0345_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ),
    .X(_0414_));
 sky130_fd_sc_hd__a221o_1 _0808_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ),
    .A2(_0338_),
    .B1(_0343_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ),
    .C1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ),
    .A2(_0342_),
    .B1(_0346_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ),
    .X(_0416_));
 sky130_fd_sc_hd__a221o_1 _0810_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ),
    .A2(_0340_),
    .B1(_0352_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ),
    .C1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a211o_1 _0811_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ),
    .A2(_0348_),
    .B1(_0415_),
    .C1(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__a221o_1 _0812_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ),
    .A2(_0347_),
    .B1(_0351_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a211o_1 _0813_ (.A1(_0276_),
    .A2(_0285_),
    .B1(_0411_),
    .C1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__o31ai_4 _0814_ (.A1(_0410_),
    .A2(_0413_),
    .A3(_0420_),
    .B1(net43),
    .Y(_0421_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(_0128_),
    .B(\CIRCUIT_1957.D0 ),
    .Y(_0422_));
 sky130_fd_sc_hd__o31a_2 _0816_ (.A1(_0112_),
    .A2(_0128_),
    .A3(_0132_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _0817_ (.A(_0421_),
    .B(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a21o_1 _0819_ (.A1(_0421_),
    .A2(_0423_),
    .B1(net53),
    .X(_0426_));
 sky130_fd_sc_hd__nand3_2 _0820_ (.A(net53),
    .B(_0421_),
    .C(_0423_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .B(_0151_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_1 _0822_ (.A1(_0426_),
    .A2(_0427_),
    .B1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand3_1 _0823_ (.A(_0426_),
    .B(_0427_),
    .C(_0428_),
    .Y(_0430_));
 sky130_fd_sc_hd__and2b_1 _0824_ (.A_N(_0429_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__and2b_1 _0825_ (.A_N(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__mux2_2 _0827_ (.A0(\CIRCUIT_1957.MEMORY_64.s_currentState ),
    .A1(net53),
    .S(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__a21o_1 _0828_ (.A1(_0430_),
    .A2(_0434_),
    .B1(_0429_),
    .X(_0435_));
 sky130_fd_sc_hd__xor2_2 _0829_ (.A(_0406_),
    .B(_0407_),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_2 _0830_ (.A(_0435_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__xor2_2 _0831_ (.A(_0384_),
    .B(_0385_),
    .X(_0438_));
 sky130_fd_sc_hd__a21oi_2 _0832_ (.A1(_0408_),
    .A2(_0437_),
    .B1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__xor2_1 _0833_ (.A(_0152_),
    .B(_0364_),
    .X(_0440_));
 sky130_fd_sc_hd__o21ai_1 _0834_ (.A1(_0386_),
    .A2(_0439_),
    .B1(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a21o_4 _0835_ (.A1(_0139_),
    .A2(_0151_),
    .B1(_0117_),
    .X(_0442_));
 sky130_fd_sc_hd__clkinv_2 _0836_ (.A(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__a21oi_1 _0837_ (.A1(_0365_),
    .A2(_0441_),
    .B1(_0443_),
    .Y(\CIRCUIT_1957.MEMORY_64.d ));
 sky130_fd_sc_hd__o21ai_1 _0838_ (.A1(_0431_),
    .A2(_0434_),
    .B1(_0442_),
    .Y(_0444_));
 sky130_fd_sc_hd__a21oi_1 _0839_ (.A1(_0431_),
    .A2(_0434_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _0840_ (.A(_0426_),
    .B(_0428_),
    .Y(_0446_));
 sky130_fd_sc_hd__or3b_1 _0841_ (.A(_0424_),
    .B(_0101_),
    .C_N(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .X(_0447_));
 sky130_fd_sc_hd__a41o_1 _0842_ (.A1(_0427_),
    .A2(_0443_),
    .A3(_0446_),
    .A4(_0447_),
    .B1(_0445_),
    .X(\CIRCUIT_1957.MEMORY_65.d ));
 sky130_fd_sc_hd__a21o_1 _0843_ (.A1(_0099_),
    .A2(_0405_),
    .B1(_0407_),
    .X(_0448_));
 sky130_fd_sc_hd__a31o_1 _0844_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A3(_0405_),
    .B1(_0442_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _0845_ (.A1(net53),
    .A2(_0404_),
    .B1(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_1 _0846_ (.A(_0435_),
    .B(_0436_),
    .X(_0451_));
 sky130_fd_sc_hd__a32o_1 _0847_ (.A1(_0437_),
    .A2(_0442_),
    .A3(_0451_),
    .B1(_0450_),
    .B2(_0448_),
    .X(\CIRCUIT_1957.MEMORY_66.d ));
 sky130_fd_sc_hd__a31o_1 _0848_ (.A1(_0408_),
    .A2(_0437_),
    .A3(_0438_),
    .B1(_0443_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_1 _0849_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ),
    .A2(_0383_),
    .B1(_0385_),
    .Y(_0453_));
 sky130_fd_sc_hd__a31o_1 _0850_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A3(_0382_),
    .B1(_0442_),
    .X(_0454_));
 sky130_fd_sc_hd__a21oi_1 _0851_ (.A1(net53),
    .A2(_0383_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__a2bb2o_1 _0852_ (.A1_N(_0439_),
    .A2_N(_0452_),
    .B1(_0453_),
    .B2(_0455_),
    .X(\CIRCUIT_1957.MEMORY_67.d ));
 sky130_fd_sc_hd__a21oi_1 _0853_ (.A1(_0099_),
    .A2(_0362_),
    .B1(_0152_),
    .Y(_0456_));
 sky130_fd_sc_hd__a311o_1 _0854_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A3(_0362_),
    .B1(_0442_),
    .C1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__o31a_1 _0855_ (.A1(_0386_),
    .A2(_0439_),
    .A3(_0440_),
    .B1(_0442_),
    .X(_0458_));
 sky130_fd_sc_hd__a2bb2o_1 _0856_ (.A1_N(_0363_),
    .A2_N(_0457_),
    .B1(_0458_),
    .B2(_0441_),
    .X(\CIRCUIT_1957.MEMORY_63.d ));
 sky130_fd_sc_hd__and3_1 _0857_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0099_),
    .C(_0134_),
    .X(\CIRCUIT_1957.MEMORY_62.d ));
 sky130_fd_sc_hd__o21a_1 _0858_ (.A1(_0145_),
    .A2(_0150_),
    .B1(\CIRCUIT_1957.MEMORY_88.s_currentState ),
    .X(\CIRCUIT_1957.GATES_60.result ));
 sky130_fd_sc_hd__and3_1 _0859_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .C(_0145_),
    .X(_0459_));
 sky130_fd_sc_hd__and3_1 _0860_ (.A(_0113_),
    .B(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .C(_0459_),
    .X(\CIRCUIT_1957.GATES_42.result ));
 sky130_fd_sc_hd__and3_2 _0861_ (.A(_0117_),
    .B(_0140_),
    .C(_0144_),
    .X(\CIRCUIT_1957.GATES_41.result ));
 sky130_fd_sc_hd__and2_2 _0862_ (.A(\CIRCUIT_1957.GATES_33.input2 ),
    .B(_0459_),
    .X(\CIRCUIT_1957.GATES_40.result ));
 sky130_fd_sc_hd__and3_2 _0863_ (.A(_0113_),
    .B(_0114_),
    .C(_0459_),
    .X(\CIRCUIT_1957.GATES_39.result ));
 sky130_fd_sc_hd__and3_1 _0864_ (.A(_0117_),
    .B(_0134_),
    .C(_0144_),
    .X(\CIRCUIT_1957.GATES_38.result ));
 sky130_fd_sc_hd__mux2_2 _0865_ (.A0(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A1(_0362_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(\CIRCUIT_1957.GATES_35.result ));
 sky130_fd_sc_hd__mux2_4 _0866_ (.A0(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A1(_0382_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(\CIRCUIT_1957.GATES_30.result ));
 sky130_fd_sc_hd__mux2_4 _0867_ (.A0(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A1(_0405_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(\CIRCUIT_1957.GATES_28.result ));
 sky130_fd_sc_hd__mux2_2 _0868_ (.A0(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .A1(_0425_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(\CIRCUIT_1957.GATES_27.result ));
 sky130_fd_sc_hd__and3_1 _0869_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .C(_0432_),
    .X(\CIRCUIT_1957.GATES_10.result ));
 sky130_fd_sc_hd__a31o_2 _0870_ (.A1(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .A2(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .A3(_0443_),
    .B1(\CIRCUIT_1957.GATES_10.result ),
    .X(\CIRCUIT_1957.GATES_9.result ));
 sky130_fd_sc_hd__nand2_2 _0871_ (.A(clknet_2_3__leaf_clk),
    .B(net43),
    .Y(_0460_));
 sky130_fd_sc_hd__and3_2 _0872_ (.A(clknet_2_2__leaf_clk),
    .B(net42),
    .C(_0338_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__and3_2 _0873_ (.A(clknet_2_3__leaf_clk),
    .B(net42),
    .C(_0348_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__and3_2 _0874_ (.A(clknet_2_3__leaf_clk),
    .B(net42),
    .C(_0347_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__and3_2 _0875_ (.A(clknet_2_3__leaf_clk),
    .B(net42),
    .C(_0336_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__nor2_2 _0876_ (.A(_0287_),
    .B(clknet_1_1__leaf__0460_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__nor2_2 _0877_ (.A(_0281_),
    .B(clknet_1_0__leaf__0460_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__and3_2 _0878_ (.A(clknet_2_3__leaf_clk),
    .B(net43),
    .C(_0285_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__nor2_2 _0879_ (.A(_0354_),
    .B(clknet_1_0__leaf__0460_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__and3_2 _0880_ (.A(clknet_2_3__leaf_clk),
    .B(net42),
    .C(_0342_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__and3_2 _0881_ (.A(clknet_2_3__leaf_clk),
    .B(net42),
    .C(_0343_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__and3_2 _0882_ (.A(clknet_2_2__leaf_clk),
    .B(net42),
    .C(_0346_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__and3_2 _0883_ (.A(clknet_2_2__leaf_clk),
    .B(net42),
    .C(_0340_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__and3_2 _0884_ (.A(clknet_2_2__leaf_clk),
    .B(net42),
    .C(_0345_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__and3_2 _0885_ (.A(clknet_2_3__leaf_clk),
    .B(net43),
    .C(_0352_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__and3_2 _0886_ (.A(clknet_2_3__leaf_clk),
    .B(net43),
    .C(_0351_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(_0103_),
    .B(net46),
    .Y(_0461_));
 sky130_fd_sc_hd__a21o_1 _0888_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ),
    .A2(net49),
    .B1(net40),
    .X(_0027_));
 sky130_fd_sc_hd__nor2_2 _0889_ (.A(_0102_),
    .B(net44),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _0890_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ),
    .A2(net49),
    .B1(net38),
    .X(_0028_));
 sky130_fd_sc_hd__nor2_2 _0891_ (.A(_0101_),
    .B(net46),
    .Y(_0463_));
 sky130_fd_sc_hd__a21o_1 _0892_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ),
    .A2(net48),
    .B1(net36),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_2 _0893_ (.A(_0100_),
    .B(net46),
    .Y(_0464_));
 sky130_fd_sc_hd__a21o_1 _0894_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ),
    .A2(net49),
    .B1(net34),
    .X(_0030_));
 sky130_fd_sc_hd__a21o_1 _0895_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ),
    .A2(net48),
    .B1(net40),
    .X(_0031_));
 sky130_fd_sc_hd__a21o_1 _0896_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ),
    .A2(net49),
    .B1(net38),
    .X(_0032_));
 sky130_fd_sc_hd__a21o_1 _0897_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ),
    .A2(net44),
    .B1(net36),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _0898_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ),
    .A2(net44),
    .B1(net34),
    .X(_0034_));
 sky130_fd_sc_hd__a21o_1 _0899_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ),
    .A2(net44),
    .B1(net40),
    .X(_0035_));
 sky130_fd_sc_hd__a21o_1 _0900_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ),
    .A2(net44),
    .B1(net38),
    .X(_0036_));
 sky130_fd_sc_hd__a21o_1 _0901_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ),
    .A2(net48),
    .B1(net36),
    .X(_0037_));
 sky130_fd_sc_hd__a21o_1 _0902_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ),
    .A2(net48),
    .B1(net34),
    .X(_0038_));
 sky130_fd_sc_hd__a21o_1 _0903_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ),
    .A2(net48),
    .B1(net40),
    .X(_0039_));
 sky130_fd_sc_hd__a21o_1 _0904_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ),
    .A2(net48),
    .B1(net38),
    .X(_0040_));
 sky130_fd_sc_hd__a21o_1 _0905_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ),
    .A2(net44),
    .B1(net36),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _0906_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ),
    .A2(net45),
    .B1(net34),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _0907_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ),
    .A2(net45),
    .B1(net40),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ),
    .A2(net45),
    .B1(net38),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _0909_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ),
    .A2(net48),
    .B1(net36),
    .X(_0045_));
 sky130_fd_sc_hd__a21o_1 _0910_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ),
    .A2(net48),
    .B1(net34),
    .X(_0046_));
 sky130_fd_sc_hd__a21o_1 _0911_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ),
    .A2(net48),
    .B1(net40),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_1 _0912_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ),
    .A2(net48),
    .B1(net38),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _0913_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ),
    .A2(net44),
    .B1(net36),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _0914_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ),
    .A2(net44),
    .B1(net34),
    .X(_0050_));
 sky130_fd_sc_hd__a21o_1 _0915_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ),
    .A2(net46),
    .B1(net40),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _0916_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ),
    .A2(net46),
    .B1(net38),
    .X(_0052_));
 sky130_fd_sc_hd__a21o_1 _0917_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ),
    .A2(net47),
    .B1(net37),
    .X(_0061_));
 sky130_fd_sc_hd__a21o_1 _0918_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ),
    .A2(net47),
    .B1(net35),
    .X(_0062_));
 sky130_fd_sc_hd__a21o_1 _0919_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ),
    .A2(net47),
    .B1(net41),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_1 _0920_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ),
    .A2(net47),
    .B1(net39),
    .X(_0064_));
 sky130_fd_sc_hd__or2_1 _0921_ (.A(net25),
    .B(net56),
    .X(_0065_));
 sky130_fd_sc_hd__and2b_1 _0922_ (.A_N(net56),
    .B(net21),
    .X(_0066_));
 sky130_fd_sc_hd__and2b_1 _0923_ (.A_N(net56),
    .B(net22),
    .X(_0067_));
 sky130_fd_sc_hd__and2b_1 _0924_ (.A_N(net56),
    .B(net24),
    .X(_0068_));
 sky130_fd_sc_hd__a21o_1 _0925_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ),
    .A2(net45),
    .B1(net36),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _0926_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ),
    .A2(net44),
    .B1(net34),
    .X(_0070_));
 sky130_fd_sc_hd__a21o_1 _0927_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ),
    .A2(net45),
    .B1(net40),
    .X(_0071_));
 sky130_fd_sc_hd__a21o_1 _0928_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ),
    .A2(net45),
    .B1(net38),
    .X(_0072_));
 sky130_fd_sc_hd__a21o_1 _0929_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ),
    .A2(net49),
    .B1(net36),
    .X(_0073_));
 sky130_fd_sc_hd__a21o_1 _0930_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ),
    .A2(net49),
    .B1(net34),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _0931_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ),
    .A2(net49),
    .B1(net40),
    .X(_0075_));
 sky130_fd_sc_hd__a21o_1 _0932_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ),
    .A2(net49),
    .B1(net38),
    .X(_0076_));
 sky130_fd_sc_hd__a21o_1 _0933_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .A2(net50),
    .B1(net36),
    .X(_0077_));
 sky130_fd_sc_hd__a21o_1 _0934_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(net50),
    .B1(net34),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_1 _0935_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .A2(net50),
    .B1(net40),
    .X(_0079_));
 sky130_fd_sc_hd__a21o_1 _0936_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .A2(net50),
    .B1(net38),
    .X(_0080_));
 sky130_fd_sc_hd__a21o_1 _0937_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(net51),
    .B1(net37),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .A2(net51),
    .B1(net35),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _0939_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .A2(net51),
    .B1(net41),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _0940_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .A2(net51),
    .B1(net39),
    .X(_0084_));
 sky130_fd_sc_hd__a21o_1 _0941_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .A2(net46),
    .B1(net37),
    .X(_0085_));
 sky130_fd_sc_hd__a21o_1 _0942_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .A2(net46),
    .B1(net35),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_1 _0943_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .A2(net46),
    .B1(net41),
    .X(_0087_));
 sky130_fd_sc_hd__a21o_1 _0944_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .A2(net47),
    .B1(net39),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _0945_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .A2(net51),
    .B1(net37),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_1 _0946_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .A2(net51),
    .B1(net35),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_1 _0947_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .A2(net51),
    .B1(net41),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_1 _0948_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .A2(net51),
    .B1(net39),
    .X(_0092_));
 sky130_fd_sc_hd__a21o_1 _0949_ (.A1(net33),
    .A2(net46),
    .B1(net37),
    .X(_0093_));
 sky130_fd_sc_hd__a21o_1 _0950_ (.A1(net32),
    .A2(net46),
    .B1(net35),
    .X(_0094_));
 sky130_fd_sc_hd__a21o_1 _0951_ (.A1(net30),
    .A2(net47),
    .B1(net41),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _0952_ (.A1(net28),
    .A2(net47),
    .B1(net39),
    .X(_0096_));
 sky130_fd_sc_hd__a21o_1 _0953_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ),
    .A2(net49),
    .B1(net36),
    .X(_0097_));
 sky130_fd_sc_hd__a21o_1 _0954_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ),
    .A2(net49),
    .B1(net34),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_2 _0955_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .X(\CIRCUIT_1957.clock_gen_2_1.GATES_3.result ));
 sky130_fd_sc_hd__nand2_2 _0956_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_2 _0957_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0958_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_2 _0959_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_2 _0960_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_2 _0961_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_2 _0962_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_2 _0963_ (.A(net54),
    .B(clknet_2_1__leaf_clk),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_2 _0964_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_2 _0965_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_2 _0966_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_2 _0967_ (.A(net54),
    .B(clknet_2_0__leaf_clk),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2_2 _0968_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_2 _0969_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_2 _0970_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_2 _0971_ (.A(net54),
    .B(clknet_2_1__leaf_clk),
    .Y(_0016_));
 sky130_fd_sc_hd__nand2_2 _0972_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_2 _0973_ (.A(net55),
    .B(clknet_2_1__leaf_clk),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0975__3 (.A(clknet_2_0__leaf_clk),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _0976__4 (.A(clknet_2_2__leaf_clk),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _0977__5 (.A(clknet_2_2__leaf_clk),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _0978__6 (.A(clknet_2_2__leaf_clk),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _0979__7 (.A(clknet_2_2__leaf_clk),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _0980__8 (.A(clknet_2_2__leaf_clk),
    .Y(net76));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0027_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0028_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0029_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0030_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0031_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0032_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0033_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0034_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0035_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0036_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0037_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0038_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0039_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0040_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0041_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0042_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0043_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0044_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0045_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0046_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0047_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0048_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0049_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0050_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0051_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0052_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ));
 sky130_fd_sc_hd__dfstp_4 _1007_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.GATES_3.result ),
    .D(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .SET_B(_0000_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1008_ (.CLK(clknet_2_0__leaf_clk),
    .D(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ),
    .RESET_B(_0001_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1009_ (.CLK(_0003_),
    .D(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ),
    .RESET_B(_0002_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1010_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D0 ),
    .RESET_B(_0004_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1011_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D1 ),
    .RESET_B(_0005_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1012_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D2 ),
    .RESET_B(_0006_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1013_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D3 ),
    .RESET_B(_0007_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1014_ (.CLK(clknet_2_1__leaf_clk),
    .D(\CIRCUIT_1957.GATES_53.result ),
    .RESET_B(_0008_),
    .Q(\CIRCUIT_1957.MEMORY_88.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_87.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_86.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_85.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_84.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_83.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_82.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_81.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_80.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_79.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_78.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_77.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_76.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1027_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .RESET_B(_0009_),
    .Q(\CIRCUIT_1957.MEMORY_75.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1028_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .RESET_B(_0010_),
    .Q(\CIRCUIT_1957.MEMORY_74.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1029_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .RESET_B(_0011_),
    .Q(\CIRCUIT_1957.MEMORY_73.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1030_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .RESET_B(_0012_),
    .Q(\CIRCUIT_1957.MEMORY_72.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1031_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .RESET_B(_0013_),
    .Q(\CIRCUIT_1957.MEMORY_71.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1032_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .RESET_B(_0014_),
    .Q(\CIRCUIT_1957.MEMORY_70.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1033_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .RESET_B(_0015_),
    .Q(\CIRCUIT_1957.MEMORY_69.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1034_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .RESET_B(_0016_),
    .Q(\CIRCUIT_1957.MEMORY_68.s_currentState ));
 sky130_fd_sc_hd__dfxtp_4 _1035_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_67.d ),
    .Q(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__dfxtp_4 _1036_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_66.d ),
    .Q(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _1037_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_65.d ),
    .Q(\CIRCUIT_1957.MEMORY_65.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1038_ (.CLK(\CIRCUIT_1957.GATES_10.result ),
    .D(\CIRCUIT_1957.MEMORY_64.d ),
    .RESET_B(_0017_),
    .Q(\CIRCUIT_1957.MEMORY_64.s_currentState ));
 sky130_fd_sc_hd__dfxtp_4 _1039_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_63.d ),
    .Q(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1040_ (.CLK(\CIRCUIT_1957.GATES_60.result ),
    .D(\CIRCUIT_1957.MEMORY_62.d ),
    .RESET_B(_0018_),
    .Q(\CIRCUIT_1957.MEMORY_62.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(net69),
    .D(_0053_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(net70),
    .D(_0054_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(net71),
    .D(_0055_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(net72),
    .D(_0056_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(net73),
    .D(_0057_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(net74),
    .D(_0058_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(net75),
    .D(_0059_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(net76),
    .D(_0060_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0061_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0062_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0063_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0064_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0065_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0066_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0067_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0068_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0069_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0070_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0071_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0072_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0073_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0074_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0075_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0076_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ));
 sky130_fd_sc_hd__dfxtp_4 _1065_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0077_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ));
 sky130_fd_sc_hd__dfxtp_4 _1066_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0078_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ));
 sky130_fd_sc_hd__dfxtp_2 _1067_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0079_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ));
 sky130_fd_sc_hd__dfxtp_4 _1068_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0080_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ));
 sky130_fd_sc_hd__dfxtp_4 _1069_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0081_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ));
 sky130_fd_sc_hd__dfxtp_2 _1070_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0082_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ));
 sky130_fd_sc_hd__dfxtp_4 _1071_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0083_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ));
 sky130_fd_sc_hd__dfxtp_4 _1072_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0084_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0085_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A0 ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0086_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A1 ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0087_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A2 ));
 sky130_fd_sc_hd__dfxtp_4 _1076_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0088_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A3 ));
 sky130_fd_sc_hd__dfxtp_4 _1077_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0089_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A4 ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0090_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A5 ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0091_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A6 ));
 sky130_fd_sc_hd__dfxtp_2 _1080_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0092_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A7 ));
 sky130_fd_sc_hd__dfxtp_4 _1081_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0093_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B0 ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0094_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B1 ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0095_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B2 ));
 sky130_fd_sc_hd__dfxtp_4 _1084_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0096_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B3 ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0097_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0098_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_68 (.HI(net68));
 sky130_fd_sc_hd__inv_2 _0482__1 (.A(clknet_2_0__leaf_clk),
    .Y(net69));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_67 (.HI(net67));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_in[8]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_in[9]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output17 (.A(net17),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_6 fanout28 (.A(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .X(net28));
 sky130_fd_sc_hd__buf_6 fanout29 (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .X(net31));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .X(net32));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(_0464_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(_0464_),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(_0463_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(_0463_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(_0462_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(_0462_),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(_0461_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(_0461_),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(_0133_),
    .X(net42));
 sky130_fd_sc_hd__buf_6 fanout43 (.A(_0133_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net52),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net52),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(net52),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net52),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__buf_4 fanout49 (.A(net51),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(_0135_),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ),
    .X(net53));
 sky130_fd_sc_hd__buf_6 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__buf_8 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 fanout56 (.A(net11),
    .X(net56));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_57 (.LO(net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0460_ (.A(_0460_),
    .X(clknet_0__0460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0460_ (.A(clknet_0__0460_),
    .X(clknet_1_0__leaf__0460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0460_ (.A(clknet_0__0460_),
    .X(clknet_1_1__leaf__0460_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_362 ();
 assign io_oeb = net67;
 assign io_out[22] = net63;
 assign io_out[23] = net64;
 assign io_out[24] = net65;
 assign io_out[25] = net66;
 assign io_out[26] = net68;
 assign io_out[4] = net57;
 assign io_out[5] = net58;
 assign io_out[6] = net59;
 assign io_out[7] = net60;
 assign io_out[8] = net61;
 assign io_out[9] = net62;
endmodule

