magic
tech sky130B
magscale 1 2
timestamp 1676595702
<< obsli1 >>
rect 1104 2159 10856 15793
<< obsm1 >>
rect 566 2128 11394 15824
<< metal2 >>
rect 2934 17200 3046 18000
rect 8914 17200 9026 18000
rect 542 0 654 800
rect 1738 0 1850 800
rect 2934 0 3046 800
rect 4130 0 4242 800
rect 5326 0 5438 800
rect 6522 0 6634 800
rect 7718 0 7830 800
rect 8914 0 9026 800
rect 10110 0 10222 800
rect 11306 0 11418 800
<< obsm2 >>
rect 572 17144 2878 17354
rect 3102 17144 8858 17354
rect 9082 17144 11388 17354
rect 572 856 11388 17144
rect 710 800 1682 856
rect 1906 800 2878 856
rect 3102 800 4074 856
rect 4298 800 5270 856
rect 5494 800 6466 856
rect 6690 800 7662 856
rect 7886 800 8858 856
rect 9082 800 10054 856
rect 10278 800 11250 856
<< metal3 >>
rect 0 15860 800 16100
rect 0 12324 800 12564
rect 0 8788 800 9028
rect 0 5252 800 5492
rect 0 1716 800 1956
<< obsm3 >>
rect 880 15780 11014 16013
rect 800 12644 11014 15780
rect 880 12244 11014 12644
rect 800 9108 11014 12244
rect 880 8708 11014 9108
rect 800 5572 11014 8708
rect 880 5172 11014 5572
rect 800 2036 11014 5172
rect 880 1803 11014 2036
<< metal4 >>
rect 2163 2128 2483 15824
rect 3382 2128 3702 15824
rect 4601 2128 4921 15824
rect 5820 2128 6140 15824
rect 7039 2128 7359 15824
rect 8258 2128 8578 15824
rect 9477 2128 9797 15824
rect 10696 2128 11016 15824
<< labels >>
rlabel metal2 s 2934 17200 3046 18000 6 clk
port 1 nsew signal input
rlabel metal3 s 0 1716 800 1956 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 5252 800 5492 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 0 12324 800 12564 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 0 15860 800 16100 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 11306 0 11418 800 6 io_oeb
port 7 nsew signal output
rlabel metal2 s 542 0 654 800 6 io_out[0]
port 8 nsew signal output
rlabel metal2 s 1738 0 1850 800 6 io_out[1]
port 9 nsew signal output
rlabel metal2 s 2934 0 3046 800 6 io_out[2]
port 10 nsew signal output
rlabel metal2 s 4130 0 4242 800 6 io_out[3]
port 11 nsew signal output
rlabel metal2 s 5326 0 5438 800 6 io_out[4]
port 12 nsew signal output
rlabel metal2 s 6522 0 6634 800 6 io_out[5]
port 13 nsew signal output
rlabel metal2 s 7718 0 7830 800 6 io_out[6]
port 14 nsew signal output
rlabel metal2 s 8914 0 9026 800 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 10110 0 10222 800 6 io_out[8]
port 16 nsew signal output
rlabel metal2 s 8914 17200 9026 18000 6 rst
port 17 nsew signal input
rlabel metal4 s 2163 2128 2483 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 3382 2128 3702 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 5820 2128 6140 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 8258 2128 8578 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 10696 2128 11016 15824 6 vssd1
port 19 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 479998
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MC14500/runs/23_02_17_02_00/results/signoff/wrapped_MC14500.magic.gds
string GDS_START 203710
<< end >>

