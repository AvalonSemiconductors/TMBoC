magic
tech sky130B
magscale 1 2
timestamp 1683538728
<< viali >>
rect 1593 15453 1627 15487
rect 1777 15317 1811 15351
rect 1593 15113 1627 15147
rect 1685 14297 1719 14331
rect 2053 14297 2087 14331
rect 1593 14025 1627 14059
rect 1685 12121 1719 12155
rect 2053 12121 2087 12155
rect 1593 11849 1627 11883
rect 5549 11849 5583 11883
rect 5641 11849 5675 11883
rect 5273 11781 5307 11815
rect 2237 11713 2271 11747
rect 2421 11713 2455 11747
rect 5457 11713 5491 11747
rect 5825 11713 5859 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 2329 11509 2363 11543
rect 6561 11509 6595 11543
rect 6009 11305 6043 11339
rect 7021 11237 7055 11271
rect 2973 11169 3007 11203
rect 4077 11169 4111 11203
rect 6561 11169 6595 11203
rect 1593 11101 1627 11135
rect 2053 11101 2087 11135
rect 2697 11101 2731 11135
rect 2789 11101 2823 11135
rect 4169 11101 4203 11135
rect 5365 11101 5399 11135
rect 5457 11101 5491 11135
rect 5733 11101 5767 11135
rect 5917 11101 5951 11135
rect 6653 11101 6687 11135
rect 4721 11033 4755 11067
rect 4445 10965 4479 10999
rect 3525 10693 3559 10727
rect 1777 10625 1811 10659
rect 1961 10625 1995 10659
rect 2053 10625 2087 10659
rect 2197 10625 2231 10659
rect 3249 10625 3283 10659
rect 3342 10625 3376 10659
rect 3617 10625 3651 10659
rect 3714 10625 3748 10659
rect 4445 10625 4479 10659
rect 4629 10625 4663 10659
rect 4905 10625 4939 10659
rect 6561 10625 6595 10659
rect 6653 10625 6687 10659
rect 2329 10489 2363 10523
rect 3893 10489 3927 10523
rect 4537 10421 4571 10455
rect 6745 10421 6779 10455
rect 6929 10421 6963 10455
rect 4445 10081 4479 10115
rect 1593 10013 1627 10047
rect 2973 10013 3007 10047
rect 3065 10013 3099 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4537 10013 4571 10047
rect 1869 9945 1903 9979
rect 3433 9877 3467 9911
rect 1593 9673 1627 9707
rect 7481 9061 7515 9095
rect 5917 8993 5951 9027
rect 6469 8993 6503 9027
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6377 8925 6411 8959
rect 6561 8925 6595 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 8585 8925 8619 8959
rect 1593 8789 1627 8823
rect 8493 8789 8527 8823
rect 1869 8517 1903 8551
rect 2881 8517 2915 8551
rect 1593 8449 1627 8483
rect 2513 8449 2547 8483
rect 2789 8449 2823 8483
rect 3801 8449 3835 8483
rect 4077 8449 4111 8483
rect 3893 8381 3927 8415
rect 3985 8381 4019 8415
rect 4261 8313 4295 8347
rect 1777 7905 1811 7939
rect 2329 7905 2363 7939
rect 4353 7905 4387 7939
rect 5273 7905 5307 7939
rect 1593 7837 1627 7871
rect 1961 7837 1995 7871
rect 2421 7837 2455 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 2973 7769 3007 7803
rect 5457 7769 5491 7803
rect 5641 7769 5675 7803
rect 4813 7497 4847 7531
rect 2145 7429 2179 7463
rect 3893 7429 3927 7463
rect 3985 7429 4019 7463
rect 5457 7429 5491 7463
rect 5641 7429 5675 7463
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 2237 7361 2271 7395
rect 2881 7361 2915 7395
rect 3065 7361 3099 7395
rect 3709 7361 3743 7395
rect 4077 7361 4111 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5365 7361 5399 7395
rect 7205 7361 7239 7395
rect 6561 7293 6595 7327
rect 7113 7293 7147 7327
rect 2421 7225 2455 7259
rect 2973 7225 3007 7259
rect 4261 7157 4295 7191
rect 5365 7157 5399 7191
rect 6377 6885 6411 6919
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 6101 6749 6135 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 6193 6681 6227 6715
rect 5181 6613 5215 6647
rect 6929 6613 6963 6647
rect 5089 6409 5123 6443
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7941 6273 7975 6307
rect 8033 6205 8067 6239
rect 7113 6137 7147 6171
rect 1593 6069 1627 6103
rect 2145 6069 2179 6103
rect 5457 6069 5491 6103
rect 7481 6069 7515 6103
rect 7941 6069 7975 6103
rect 8309 6069 8343 6103
rect 5365 5865 5399 5899
rect 2237 5729 2271 5763
rect 1685 5661 1719 5695
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 5181 5593 5215 5627
rect 5381 5593 5415 5627
rect 2973 5525 3007 5559
rect 5549 5525 5583 5559
rect 1961 5321 1995 5355
rect 2789 5321 2823 5355
rect 1777 5185 1811 5219
rect 1961 5185 1995 5219
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 3157 4981 3191 5015
rect 4537 4709 4571 4743
rect 5641 4709 5675 4743
rect 6009 4641 6043 4675
rect 1593 4573 1627 4607
rect 1777 4573 1811 4607
rect 1961 4573 1995 4607
rect 2789 4573 2823 4607
rect 3433 4573 3467 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 7573 4573 7607 4607
rect 1869 4505 1903 4539
rect 4537 4505 4571 4539
rect 2145 4437 2179 4471
rect 2697 4437 2731 4471
rect 3341 4437 3375 4471
rect 5549 4437 5583 4471
rect 7481 4437 7515 4471
rect 1685 4233 1719 4267
rect 4645 4233 4679 4267
rect 5641 4233 5675 4267
rect 2329 4165 2363 4199
rect 4445 4165 4479 4199
rect 1869 4097 1903 4131
rect 2605 4097 2639 4131
rect 3617 4097 3651 4131
rect 5549 4097 5583 4131
rect 5825 4097 5859 4131
rect 6745 4097 6779 4131
rect 6929 4097 6963 4131
rect 7389 4097 7423 4131
rect 7481 4097 7515 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8585 4097 8619 4131
rect 2513 4029 2547 4063
rect 3249 4029 3283 4063
rect 3801 4029 3835 4063
rect 6009 4029 6043 4063
rect 2789 3961 2823 3995
rect 3341 3961 3375 3995
rect 2605 3893 2639 3927
rect 4629 3893 4663 3927
rect 4813 3893 4847 3927
rect 6837 3893 6871 3927
rect 8769 3893 8803 3927
rect 2329 3689 2363 3723
rect 4169 3689 4203 3723
rect 3985 3621 4019 3655
rect 2421 3553 2455 3587
rect 5641 3553 5675 3587
rect 6101 3553 6135 3587
rect 7481 3553 7515 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 2145 3485 2179 3519
rect 3249 3485 3283 3519
rect 3433 3485 3467 3519
rect 4905 3485 4939 3519
rect 5089 3485 5123 3519
rect 5733 3485 5767 3519
rect 7389 3485 7423 3519
rect 9321 3485 9355 3519
rect 4137 3417 4171 3451
rect 4353 3417 4387 3451
rect 1961 3349 1995 3383
rect 3341 3349 3375 3383
rect 4997 3349 5031 3383
rect 7757 3349 7791 3383
rect 2513 3145 2547 3179
rect 2053 3009 2087 3043
rect 2513 3009 2547 3043
rect 2697 3009 2731 3043
rect 3157 3009 3191 3043
rect 9873 3009 9907 3043
rect 1777 2941 1811 2975
rect 3249 2941 3283 2975
rect 10149 2941 10183 2975
rect 1777 2601 1811 2635
rect 3249 2465 3283 2499
rect 1593 2397 1627 2431
rect 2329 2397 2363 2431
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 6745 2397 6779 2431
rect 8125 2397 8159 2431
rect 9689 2397 9723 2431
rect 2605 2329 2639 2363
rect 4261 2329 4295 2363
rect 5549 2329 5583 2363
rect 7021 2329 7055 2363
rect 8401 2329 8435 2363
rect 9965 2329 9999 2363
<< metal1 >>
rect 1104 15802 10856 15824
rect 1104 15750 2169 15802
rect 2221 15750 2233 15802
rect 2285 15750 2297 15802
rect 2349 15750 2361 15802
rect 2413 15750 2425 15802
rect 2477 15750 4607 15802
rect 4659 15750 4671 15802
rect 4723 15750 4735 15802
rect 4787 15750 4799 15802
rect 4851 15750 4863 15802
rect 4915 15750 7045 15802
rect 7097 15750 7109 15802
rect 7161 15750 7173 15802
rect 7225 15750 7237 15802
rect 7289 15750 7301 15802
rect 7353 15750 9483 15802
rect 9535 15750 9547 15802
rect 9599 15750 9611 15802
rect 9663 15750 9675 15802
rect 9727 15750 9739 15802
rect 9791 15750 10856 15802
rect 1104 15728 10856 15750
rect 934 15444 940 15496
rect 992 15484 998 15496
rect 1578 15484 1584 15496
rect 992 15456 1584 15484
rect 992 15444 998 15456
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 1765 15351 1823 15357
rect 1765 15317 1777 15351
rect 1811 15348 1823 15351
rect 5442 15348 5448 15360
rect 1811 15320 5448 15348
rect 1811 15317 1823 15320
rect 1765 15311 1823 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 1104 15258 11016 15280
rect 1104 15206 3388 15258
rect 3440 15206 3452 15258
rect 3504 15206 3516 15258
rect 3568 15206 3580 15258
rect 3632 15206 3644 15258
rect 3696 15206 5826 15258
rect 5878 15206 5890 15258
rect 5942 15206 5954 15258
rect 6006 15206 6018 15258
rect 6070 15206 6082 15258
rect 6134 15206 8264 15258
rect 8316 15206 8328 15258
rect 8380 15206 8392 15258
rect 8444 15206 8456 15258
rect 8508 15206 8520 15258
rect 8572 15206 10702 15258
rect 10754 15206 10766 15258
rect 10818 15206 10830 15258
rect 10882 15206 10894 15258
rect 10946 15206 10958 15258
rect 11010 15206 11016 15258
rect 1104 15184 11016 15206
rect 1578 15104 1584 15156
rect 1636 15104 1642 15156
rect 1104 14714 10856 14736
rect 1104 14662 2169 14714
rect 2221 14662 2233 14714
rect 2285 14662 2297 14714
rect 2349 14662 2361 14714
rect 2413 14662 2425 14714
rect 2477 14662 4607 14714
rect 4659 14662 4671 14714
rect 4723 14662 4735 14714
rect 4787 14662 4799 14714
rect 4851 14662 4863 14714
rect 4915 14662 7045 14714
rect 7097 14662 7109 14714
rect 7161 14662 7173 14714
rect 7225 14662 7237 14714
rect 7289 14662 7301 14714
rect 7353 14662 9483 14714
rect 9535 14662 9547 14714
rect 9599 14662 9611 14714
rect 9663 14662 9675 14714
rect 9727 14662 9739 14714
rect 9791 14662 10856 14714
rect 1104 14640 10856 14662
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1673 14331 1731 14337
rect 1673 14328 1685 14331
rect 992 14300 1685 14328
rect 992 14288 998 14300
rect 1673 14297 1685 14300
rect 1719 14297 1731 14331
rect 1673 14291 1731 14297
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14328 2099 14331
rect 2682 14328 2688 14340
rect 2087 14300 2688 14328
rect 2087 14297 2099 14300
rect 2041 14291 2099 14297
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 1104 14170 11016 14192
rect 1104 14118 3388 14170
rect 3440 14118 3452 14170
rect 3504 14118 3516 14170
rect 3568 14118 3580 14170
rect 3632 14118 3644 14170
rect 3696 14118 5826 14170
rect 5878 14118 5890 14170
rect 5942 14118 5954 14170
rect 6006 14118 6018 14170
rect 6070 14118 6082 14170
rect 6134 14118 8264 14170
rect 8316 14118 8328 14170
rect 8380 14118 8392 14170
rect 8444 14118 8456 14170
rect 8508 14118 8520 14170
rect 8572 14118 10702 14170
rect 10754 14118 10766 14170
rect 10818 14118 10830 14170
rect 10882 14118 10894 14170
rect 10946 14118 10958 14170
rect 11010 14118 11016 14170
rect 1104 14096 11016 14118
rect 934 14016 940 14068
rect 992 14056 998 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 992 14028 1593 14056
rect 992 14016 998 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 1104 13626 10856 13648
rect 1104 13574 2169 13626
rect 2221 13574 2233 13626
rect 2285 13574 2297 13626
rect 2349 13574 2361 13626
rect 2413 13574 2425 13626
rect 2477 13574 4607 13626
rect 4659 13574 4671 13626
rect 4723 13574 4735 13626
rect 4787 13574 4799 13626
rect 4851 13574 4863 13626
rect 4915 13574 7045 13626
rect 7097 13574 7109 13626
rect 7161 13574 7173 13626
rect 7225 13574 7237 13626
rect 7289 13574 7301 13626
rect 7353 13574 9483 13626
rect 9535 13574 9547 13626
rect 9599 13574 9611 13626
rect 9663 13574 9675 13626
rect 9727 13574 9739 13626
rect 9791 13574 10856 13626
rect 1104 13552 10856 13574
rect 1104 13082 11016 13104
rect 1104 13030 3388 13082
rect 3440 13030 3452 13082
rect 3504 13030 3516 13082
rect 3568 13030 3580 13082
rect 3632 13030 3644 13082
rect 3696 13030 5826 13082
rect 5878 13030 5890 13082
rect 5942 13030 5954 13082
rect 6006 13030 6018 13082
rect 6070 13030 6082 13082
rect 6134 13030 8264 13082
rect 8316 13030 8328 13082
rect 8380 13030 8392 13082
rect 8444 13030 8456 13082
rect 8508 13030 8520 13082
rect 8572 13030 10702 13082
rect 10754 13030 10766 13082
rect 10818 13030 10830 13082
rect 10882 13030 10894 13082
rect 10946 13030 10958 13082
rect 11010 13030 11016 13082
rect 1104 13008 11016 13030
rect 1104 12538 10856 12560
rect 1104 12486 2169 12538
rect 2221 12486 2233 12538
rect 2285 12486 2297 12538
rect 2349 12486 2361 12538
rect 2413 12486 2425 12538
rect 2477 12486 4607 12538
rect 4659 12486 4671 12538
rect 4723 12486 4735 12538
rect 4787 12486 4799 12538
rect 4851 12486 4863 12538
rect 4915 12486 7045 12538
rect 7097 12486 7109 12538
rect 7161 12486 7173 12538
rect 7225 12486 7237 12538
rect 7289 12486 7301 12538
rect 7353 12486 9483 12538
rect 9535 12486 9547 12538
rect 9599 12486 9611 12538
rect 9663 12486 9675 12538
rect 9727 12486 9739 12538
rect 9791 12486 10856 12538
rect 1104 12464 10856 12486
rect 934 12112 940 12164
rect 992 12152 998 12164
rect 1673 12155 1731 12161
rect 1673 12152 1685 12155
rect 992 12124 1685 12152
rect 992 12112 998 12124
rect 1673 12121 1685 12124
rect 1719 12121 1731 12155
rect 1673 12115 1731 12121
rect 2038 12112 2044 12164
rect 2096 12112 2102 12164
rect 1104 11994 11016 12016
rect 1104 11942 3388 11994
rect 3440 11942 3452 11994
rect 3504 11942 3516 11994
rect 3568 11942 3580 11994
rect 3632 11942 3644 11994
rect 3696 11942 5826 11994
rect 5878 11942 5890 11994
rect 5942 11942 5954 11994
rect 6006 11942 6018 11994
rect 6070 11942 6082 11994
rect 6134 11942 8264 11994
rect 8316 11942 8328 11994
rect 8380 11942 8392 11994
rect 8444 11942 8456 11994
rect 8508 11942 8520 11994
rect 8572 11942 10702 11994
rect 10754 11942 10766 11994
rect 10818 11942 10830 11994
rect 10882 11942 10894 11994
rect 10946 11942 10958 11994
rect 11010 11942 11016 11994
rect 1104 11920 11016 11942
rect 934 11840 940 11892
rect 992 11880 998 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 992 11852 1593 11880
rect 992 11840 998 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5500 11852 5549 11880
rect 5500 11840 5506 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 5537 11843 5595 11849
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 5261 11815 5319 11821
rect 5261 11812 5273 11815
rect 2740 11784 5273 11812
rect 2740 11772 2746 11784
rect 5261 11781 5273 11784
rect 5307 11812 5319 11815
rect 5902 11812 5908 11824
rect 5307 11784 5908 11812
rect 5307 11781 5319 11784
rect 5261 11775 5319 11781
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2096 11716 2237 11744
rect 2096 11704 2102 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6454 11744 6460 11756
rect 5859 11716 6460 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6454 11704 6460 11716
rect 6512 11744 6518 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6512 11716 6561 11744
rect 6512 11704 6518 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11540 2375 11543
rect 3234 11540 3240 11552
rect 2363 11512 3240 11540
rect 2363 11509 2375 11512
rect 2317 11503 2375 11509
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 6546 11500 6552 11552
rect 6604 11500 6610 11552
rect 1104 11450 10856 11472
rect 1104 11398 2169 11450
rect 2221 11398 2233 11450
rect 2285 11398 2297 11450
rect 2349 11398 2361 11450
rect 2413 11398 2425 11450
rect 2477 11398 4607 11450
rect 4659 11398 4671 11450
rect 4723 11398 4735 11450
rect 4787 11398 4799 11450
rect 4851 11398 4863 11450
rect 4915 11398 7045 11450
rect 7097 11398 7109 11450
rect 7161 11398 7173 11450
rect 7225 11398 7237 11450
rect 7289 11398 7301 11450
rect 7353 11398 9483 11450
rect 9535 11398 9547 11450
rect 9599 11398 9611 11450
rect 9663 11398 9675 11450
rect 9727 11398 9739 11450
rect 9791 11398 10856 11450
rect 1104 11376 10856 11398
rect 5997 11339 6055 11345
rect 5997 11305 6009 11339
rect 6043 11336 6055 11339
rect 6730 11336 6736 11348
rect 6043 11308 6736 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7926 11268 7932 11280
rect 7055 11240 7932 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 2958 11160 2964 11212
rect 3016 11160 3022 11212
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4246 11200 4252 11212
rect 4111 11172 4252 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5626 11200 5632 11212
rect 5276 11172 5632 11200
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1581 11135 1639 11141
rect 1581 11132 1593 11135
rect 1544 11104 1593 11132
rect 1544 11092 1550 11104
rect 1581 11101 1593 11104
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2038 11092 2044 11144
rect 2096 11092 2102 11144
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 2823 11104 4169 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 4157 11101 4169 11104
rect 4203 11132 4215 11135
rect 5276 11132 5304 11172
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 5684 11172 5764 11200
rect 5684 11160 5690 11172
rect 4203 11104 5304 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 2498 11064 2504 11076
rect 1912 11036 2504 11064
rect 1912 11024 1918 11036
rect 2498 11024 2504 11036
rect 2556 11064 2562 11076
rect 2792 11064 2820 11095
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 5442 11092 5448 11144
rect 5500 11092 5506 11144
rect 5736 11141 5764 11172
rect 6546 11160 6552 11212
rect 6604 11160 6610 11212
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 2556 11036 2820 11064
rect 2556 11024 2562 11036
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 4709 11067 4767 11073
rect 4709 11064 4721 11067
rect 3016 11036 4721 11064
rect 3016 11024 3022 11036
rect 4709 11033 4721 11036
rect 4755 11064 4767 11067
rect 4890 11064 4896 11076
rect 4755 11036 4896 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5368 11064 5396 11092
rect 6546 11064 6552 11076
rect 5368 11036 6552 11064
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 6656 11008 6684 11095
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10996 4491 10999
rect 6638 10996 6644 11008
rect 4479 10968 6644 10996
rect 4479 10965 4491 10968
rect 4433 10959 4491 10965
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 1104 10906 11016 10928
rect 1104 10854 3388 10906
rect 3440 10854 3452 10906
rect 3504 10854 3516 10906
rect 3568 10854 3580 10906
rect 3632 10854 3644 10906
rect 3696 10854 5826 10906
rect 5878 10854 5890 10906
rect 5942 10854 5954 10906
rect 6006 10854 6018 10906
rect 6070 10854 6082 10906
rect 6134 10854 8264 10906
rect 8316 10854 8328 10906
rect 8380 10854 8392 10906
rect 8444 10854 8456 10906
rect 8508 10854 8520 10906
rect 8572 10854 10702 10906
rect 10754 10854 10766 10906
rect 10818 10854 10830 10906
rect 10882 10854 10894 10906
rect 10946 10854 10958 10906
rect 11010 10854 11016 10906
rect 1104 10832 11016 10854
rect 3513 10727 3571 10733
rect 1780 10696 3464 10724
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1780 10665 1808 10696
rect 1765 10659 1823 10665
rect 1765 10656 1777 10659
rect 1544 10628 1777 10656
rect 1544 10616 1550 10628
rect 1765 10625 1777 10628
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1912 10628 1961 10656
rect 1912 10616 1918 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2038 10616 2044 10668
rect 2096 10616 2102 10668
rect 2185 10659 2243 10665
rect 2185 10625 2197 10659
rect 2231 10656 2243 10659
rect 2682 10656 2688 10668
rect 2231 10628 2688 10656
rect 2231 10625 2243 10628
rect 2185 10619 2243 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3330 10659 3388 10665
rect 3330 10625 3342 10659
rect 3376 10625 3388 10659
rect 3436 10656 3464 10696
rect 3513 10693 3525 10727
rect 3559 10724 3571 10727
rect 3559 10696 4016 10724
rect 3559 10693 3571 10696
rect 3513 10687 3571 10693
rect 3988 10668 4016 10696
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3436 10628 3617 10656
rect 3330 10619 3388 10625
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 3702 10659 3760 10665
rect 3702 10625 3714 10659
rect 3748 10656 3760 10659
rect 3748 10628 3832 10656
rect 3748 10625 3760 10628
rect 3702 10619 3760 10625
rect 3050 10588 3056 10600
rect 2332 10560 3056 10588
rect 2332 10529 2360 10560
rect 3050 10548 3056 10560
rect 3108 10588 3114 10600
rect 3344 10588 3372 10619
rect 3108 10560 3372 10588
rect 3804 10588 3832 10628
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 4246 10656 4252 10668
rect 4028 10628 4252 10656
rect 4028 10616 4034 10628
rect 4246 10616 4252 10628
rect 4304 10656 4310 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4304 10628 4445 10656
rect 4304 10616 4310 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4580 10628 4629 10656
rect 4580 10616 4586 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4890 10616 4896 10668
rect 4948 10616 4954 10668
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6512 10628 6561 10656
rect 6512 10616 6518 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 5534 10588 5540 10600
rect 3804 10560 5540 10588
rect 3108 10548 3114 10560
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 2682 10480 2688 10532
rect 2740 10520 2746 10532
rect 3804 10520 3832 10560
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 2740 10492 3832 10520
rect 3881 10523 3939 10529
rect 2740 10480 2746 10492
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 5442 10520 5448 10532
rect 3927 10492 5448 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 4120 10424 4537 10452
rect 4120 10412 4126 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 4525 10415 4583 10421
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 6914 10412 6920 10464
rect 6972 10412 6978 10464
rect 1104 10362 10856 10384
rect 1104 10310 2169 10362
rect 2221 10310 2233 10362
rect 2285 10310 2297 10362
rect 2349 10310 2361 10362
rect 2413 10310 2425 10362
rect 2477 10310 4607 10362
rect 4659 10310 4671 10362
rect 4723 10310 4735 10362
rect 4787 10310 4799 10362
rect 4851 10310 4863 10362
rect 4915 10310 7045 10362
rect 7097 10310 7109 10362
rect 7161 10310 7173 10362
rect 7225 10310 7237 10362
rect 7289 10310 7301 10362
rect 7353 10310 9483 10362
rect 9535 10310 9547 10362
rect 9599 10310 9611 10362
rect 9663 10310 9675 10362
rect 9727 10310 9739 10362
rect 9791 10310 10856 10362
rect 1104 10288 10856 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 4522 10248 4528 10260
rect 3108 10220 4528 10248
rect 3108 10208 3114 10220
rect 3234 10140 3240 10192
rect 3292 10140 3298 10192
rect 3252 10112 3280 10140
rect 3252 10084 4200 10112
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 1578 10044 1584 10056
rect 992 10016 1584 10044
rect 992 10004 998 10016
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3970 10044 3976 10056
rect 3283 10016 3976 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 1486 9936 1492 9988
rect 1544 9976 1550 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1544 9948 1869 9976
rect 1544 9936 1550 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 3252 9976 3280 10007
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4172 10053 4200 10084
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4264 10044 4292 10220
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5626 10112 5632 10124
rect 4479 10084 5632 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4264 10016 4537 10044
rect 4157 10007 4215 10013
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 1857 9939 1915 9945
rect 2976 9948 3280 9976
rect 2976 9920 3004 9948
rect 2958 9868 2964 9920
rect 3016 9868 3022 9920
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3878 9908 3884 9920
rect 3467 9880 3884 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 1578 9664 1584 9716
rect 1636 9664 1642 9716
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 7374 9092 7380 9104
rect 5920 9064 7380 9092
rect 5920 9033 5948 9064
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 7469 9095 7527 9101
rect 7469 9061 7481 9095
rect 7515 9092 7527 9095
rect 7515 9064 8616 9092
rect 7515 9061 7527 9064
rect 7469 9055 7527 9061
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6503 8996 7604 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 6380 8888 6408 8919
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6972 8928 7021 8956
rect 6972 8916 6978 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7374 8956 7380 8968
rect 7239 8928 7380 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 1912 8860 6408 8888
rect 7024 8888 7052 8919
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7576 8965 7604 8996
rect 8588 8965 8616 9064
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8956 7619 8959
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7607 8928 8033 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8846 8956 8852 8968
rect 8619 8928 8852 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8220 8888 8248 8919
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 7024 8860 8248 8888
rect 1912 8848 1918 8860
rect 934 8780 940 8832
rect 992 8820 998 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 992 8792 1593 8820
rect 992 8780 998 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 8662 8820 8668 8832
rect 8527 8792 8668 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 4982 8616 4988 8628
rect 2884 8588 4988 8616
rect 1854 8508 1860 8560
rect 1912 8508 1918 8560
rect 2884 8557 2912 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8517 2927 8551
rect 4430 8548 4436 8560
rect 2869 8511 2927 8517
rect 3804 8520 4436 8548
rect 934 8440 940 8492
rect 992 8480 998 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 992 8452 1593 8480
rect 992 8440 998 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 3804 8489 3832 8520
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 2648 8452 2789 8480
rect 2648 8440 2654 8452
rect 2777 8449 2789 8452
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 3896 8344 3924 8375
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4080 8412 4108 8443
rect 4080 8384 4200 8412
rect 4062 8344 4068 8356
rect 3896 8316 4068 8344
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4172 8276 4200 8384
rect 4249 8347 4307 8353
rect 4249 8313 4261 8347
rect 4295 8344 4307 8347
rect 5258 8344 5264 8356
rect 4295 8316 5264 8344
rect 4295 8313 4307 8316
rect 4249 8307 4307 8313
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 3936 8248 4200 8276
rect 3936 8236 3942 8248
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 4062 8032 4068 8084
rect 4120 8032 4126 8084
rect 4080 8004 4108 8032
rect 4080 7976 4292 8004
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 1765 7939 1823 7945
rect 1765 7936 1777 7939
rect 1544 7908 1777 7936
rect 1544 7896 1550 7908
rect 1765 7905 1777 7908
rect 1811 7905 1823 7939
rect 1765 7899 1823 7905
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2682 7936 2688 7948
rect 2363 7908 2688 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2590 7868 2596 7880
rect 2455 7840 2596 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 1670 7760 1676 7812
rect 1728 7800 1734 7812
rect 2424 7800 2452 7831
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 4120 7840 4169 7868
rect 4120 7828 4126 7840
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 1728 7772 2452 7800
rect 1728 7760 1734 7772
rect 2958 7760 2964 7812
rect 3016 7760 3022 7812
rect 3786 7760 3792 7812
rect 3844 7800 3850 7812
rect 4264 7800 4292 7976
rect 4338 7896 4344 7948
rect 4396 7896 4402 7948
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 4540 7908 5273 7936
rect 4540 7880 4568 7908
rect 5261 7905 5273 7908
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4816 7800 4844 7831
rect 3844 7772 4844 7800
rect 3844 7760 3850 7772
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 5040 7772 5457 7800
rect 5040 7760 5046 7772
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 5445 7763 5503 7769
rect 5629 7803 5687 7809
rect 5629 7769 5641 7803
rect 5675 7769 5687 7803
rect 5629 7763 5687 7769
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 5644 7732 5672 7763
rect 4764 7704 5672 7732
rect 4764 7692 4770 7704
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4488 7500 4813 7528
rect 4488 7488 4494 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2133 7463 2191 7469
rect 2133 7460 2145 7463
rect 1636 7432 2145 7460
rect 1636 7420 1642 7432
rect 2133 7429 2145 7432
rect 2179 7460 2191 7463
rect 2179 7432 3096 7460
rect 2179 7429 2191 7432
rect 2133 7423 2191 7429
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1728 7364 1869 7392
rect 1728 7352 1734 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2038 7352 2044 7404
rect 2096 7352 2102 7404
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 2498 7392 2504 7404
rect 2271 7364 2504 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3068 7401 3096 7432
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 3973 7463 4031 7469
rect 3973 7429 3985 7463
rect 4019 7460 4031 7463
rect 4522 7460 4528 7472
rect 4019 7432 4528 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 4632 7432 4936 7460
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3786 7392 3792 7404
rect 3743 7364 3792 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4430 7352 4436 7404
rect 4488 7392 4494 7404
rect 4632 7392 4660 7432
rect 4488 7364 4660 7392
rect 4488 7352 4494 7364
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4908 7401 4936 7432
rect 5442 7420 5448 7472
rect 5500 7420 5506 7472
rect 5626 7420 5632 7472
rect 5684 7420 5690 7472
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 4982 7392 4988 7404
rect 4939 7364 4988 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 4080 7324 4108 7352
rect 2424 7296 4108 7324
rect 2424 7265 2452 7296
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7225 2467 7259
rect 2409 7219 2467 7225
rect 2961 7259 3019 7265
rect 2961 7225 2973 7259
rect 3007 7256 3019 7259
rect 4724 7256 4752 7352
rect 5368 7324 5396 7355
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6880 7364 7205 7392
rect 6880 7352 6886 7364
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 7374 7392 7380 7404
rect 7239 7364 7380 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 6362 7324 6368 7336
rect 5368 7296 6368 7324
rect 6362 7284 6368 7296
rect 6420 7324 6426 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 6420 7296 6561 7324
rect 6420 7284 6426 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 6549 7287 6607 7293
rect 6886 7296 7113 7324
rect 6886 7268 6914 7296
rect 7101 7293 7113 7296
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 6886 7256 6920 7268
rect 3007 7228 6920 7256
rect 3007 7225 3019 7228
rect 2961 7219 3019 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 4246 7148 4252 7200
rect 4304 7148 4310 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 5040 7160 5365 7188
rect 5040 7148 5046 7160
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 5353 7151 5411 7157
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2866 6984 2872 6996
rect 2096 6956 2872 6984
rect 2096 6944 2102 6956
rect 2866 6944 2872 6956
rect 2924 6984 2930 6996
rect 6546 6984 6552 6996
rect 2924 6956 6552 6984
rect 2924 6944 2930 6956
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6365 6919 6423 6925
rect 6365 6885 6377 6919
rect 6411 6914 6423 6919
rect 6411 6886 6445 6914
rect 6411 6885 6423 6886
rect 6365 6879 6423 6885
rect 6380 6848 6408 6879
rect 7098 6848 7104 6860
rect 5368 6820 6224 6848
rect 6380 6820 7104 6848
rect 5368 6789 5396 6820
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5684 6752 6101 6780
rect 5684 6740 5690 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6196 6780 6224 6820
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 6362 6780 6368 6792
rect 6196 6752 6368 6780
rect 6089 6743 6147 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6972 6752 7021 6780
rect 6972 6740 6978 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 5552 6712 5580 6740
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5552 6684 6193 6712
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 6181 6675 6239 6681
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 5132 6616 5181 6644
rect 5132 6604 5138 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7006 6644 7012 6656
rect 6963 6616 7012 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 5074 6400 5080 6452
rect 5132 6400 5138 6452
rect 4982 6264 4988 6316
rect 5040 6264 5046 6316
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6304 7343 6307
rect 7926 6304 7932 6316
rect 7331 6276 7932 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 7024 6236 7052 6264
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7024 6208 8033 6236
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7156 6140 7972 6168
rect 7156 6128 7162 6140
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 992 6072 1593 6100
rect 992 6060 998 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2133 6103 2191 6109
rect 2133 6100 2145 6103
rect 1912 6072 2145 6100
rect 1912 6060 1918 6072
rect 2133 6069 2145 6072
rect 2179 6069 2191 6103
rect 2133 6063 2191 6069
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5626 6100 5632 6112
rect 5491 6072 5632 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7469 6103 7527 6109
rect 7469 6069 7481 6103
rect 7515 6100 7527 6103
rect 7558 6100 7564 6112
rect 7515 6072 7564 6100
rect 7515 6069 7527 6072
rect 7469 6063 7527 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7944 6109 7972 6140
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8754 6100 8760 6112
rect 8343 6072 8760 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5040 5868 5365 5896
rect 5040 5856 5046 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2682 5760 2688 5772
rect 2271 5732 2688 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2682 5720 2688 5732
rect 2740 5760 2746 5772
rect 2740 5732 3188 5760
rect 2740 5720 2746 5732
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 992 5664 1685 5692
rect 992 5652 998 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3050 5692 3056 5704
rect 3007 5664 3056 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3160 5701 3188 5732
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 5074 5584 5080 5636
rect 5132 5624 5138 5636
rect 5169 5627 5227 5633
rect 5169 5624 5181 5627
rect 5132 5596 5181 5624
rect 5132 5584 5138 5596
rect 5169 5593 5181 5596
rect 5215 5593 5227 5627
rect 5169 5587 5227 5593
rect 5258 5584 5264 5636
rect 5316 5624 5322 5636
rect 5369 5627 5427 5633
rect 5369 5624 5381 5627
rect 5316 5596 5381 5624
rect 5316 5584 5322 5596
rect 5369 5593 5381 5596
rect 5415 5593 5427 5627
rect 5369 5587 5427 5593
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 2961 5559 3019 5565
rect 2961 5556 2973 5559
rect 2924 5528 2973 5556
rect 2924 5516 2930 5528
rect 2961 5525 2973 5528
rect 3007 5525 3019 5559
rect 2961 5519 3019 5525
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2498 5352 2504 5364
rect 1995 5324 2504 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2498 5312 2504 5324
rect 2556 5352 2562 5364
rect 2777 5355 2835 5361
rect 2777 5352 2789 5355
rect 2556 5324 2789 5352
rect 2556 5312 2562 5324
rect 2777 5321 2789 5324
rect 2823 5321 2835 5355
rect 2777 5315 2835 5321
rect 2866 5284 2872 5296
rect 2700 5256 2872 5284
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1762 5216 1768 5228
rect 1636 5188 1768 5216
rect 1636 5176 1642 5188
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 2700 5225 2728 5256
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2958 5176 2964 5228
rect 3016 5176 3022 5228
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 3050 5148 3056 5160
rect 1544 5120 3056 5148
rect 1544 5108 1550 5120
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3786 5012 3792 5024
rect 3191 4984 3792 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 4522 4700 4528 4752
rect 4580 4700 4586 4752
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5592 4644 6009 4672
rect 5592 4632 5598 4644
rect 5997 4641 6009 4644
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1544 4576 1593 4604
rect 1544 4564 1550 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 1946 4564 1952 4616
rect 2004 4564 2010 4616
rect 2774 4564 2780 4616
rect 2832 4564 2838 4616
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3108 4576 3433 4604
rect 3108 4564 3114 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 7558 4564 7564 4616
rect 7616 4564 7622 4616
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 1857 4539 1915 4545
rect 1857 4536 1869 4539
rect 1728 4508 1869 4536
rect 1728 4496 1734 4508
rect 1857 4505 1869 4508
rect 1903 4505 1915 4539
rect 1857 4499 1915 4505
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4525 4539 4583 4545
rect 4525 4536 4537 4539
rect 4120 4508 4537 4536
rect 4120 4496 4126 4508
rect 4525 4505 4537 4508
rect 4571 4505 4583 4539
rect 4525 4499 4583 4505
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 2133 4471 2191 4477
rect 2133 4468 2145 4471
rect 2096 4440 2145 4468
rect 2096 4428 2102 4440
rect 2133 4437 2145 4440
rect 2179 4437 2191 4471
rect 2133 4431 2191 4437
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 2648 4440 2697 4468
rect 2648 4428 2654 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 2685 4431 2743 4437
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3329 4471 3387 4477
rect 3329 4468 3341 4471
rect 2832 4440 3341 4468
rect 2832 4428 2838 4440
rect 3329 4437 3341 4440
rect 3375 4437 3387 4471
rect 3329 4431 3387 4437
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5718 4468 5724 4480
rect 5583 4440 5724 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7248 4440 7481 4468
rect 7248 4428 7254 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7469 4431 7527 4437
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1762 4264 1768 4276
rect 1719 4236 1768 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1762 4224 1768 4236
rect 1820 4224 1826 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4633 4267 4691 4273
rect 4633 4264 4645 4267
rect 4304 4236 4645 4264
rect 4304 4224 4310 4236
rect 4633 4233 4645 4236
rect 4679 4233 4691 4267
rect 4633 4227 4691 4233
rect 5626 4224 5632 4276
rect 5684 4224 5690 4276
rect 2317 4199 2375 4205
rect 2317 4165 2329 4199
rect 2363 4196 2375 4199
rect 2498 4196 2504 4208
rect 2363 4168 2504 4196
rect 2363 4165 2375 4168
rect 2317 4159 2375 4165
rect 2498 4156 2504 4168
rect 2556 4196 2562 4208
rect 2682 4196 2688 4208
rect 2556 4168 2688 4196
rect 2556 4156 2562 4168
rect 2682 4156 2688 4168
rect 2740 4156 2746 4208
rect 3326 4156 3332 4208
rect 3384 4196 3390 4208
rect 4062 4196 4068 4208
rect 3384 4168 4068 4196
rect 3384 4156 3390 4168
rect 4062 4156 4068 4168
rect 4120 4196 4126 4208
rect 4433 4199 4491 4205
rect 4433 4196 4445 4199
rect 4120 4168 4445 4196
rect 4120 4156 4126 4168
rect 4433 4165 4445 4168
rect 4479 4165 4491 4199
rect 7190 4196 7196 4208
rect 4433 4159 4491 4165
rect 6840 4168 7196 4196
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 1854 4128 1860 4140
rect 992 4100 1860 4128
rect 992 4088 998 4100
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2774 4128 2780 4140
rect 2639 4100 2780 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3160 4100 3617 4128
rect 2498 4020 2504 4072
rect 2556 4020 2562 4072
rect 3160 4060 3188 4100
rect 3605 4097 3617 4100
rect 3651 4128 3663 4131
rect 4154 4128 4160 4140
rect 3651 4100 4160 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5092 4100 5549 4128
rect 2792 4032 3188 4060
rect 3237 4063 3295 4069
rect 2792 4001 2820 4032
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3283 4032 3740 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 2777 3995 2835 4001
rect 2777 3961 2789 3995
rect 2823 3961 2835 3995
rect 2777 3955 2835 3961
rect 3326 3952 3332 4004
rect 3384 3952 3390 4004
rect 3712 3992 3740 4032
rect 3786 4020 3792 4072
rect 3844 4020 3850 4072
rect 4430 3992 4436 4004
rect 3712 3964 4436 3992
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 5092 3936 5120 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5684 4100 5825 4128
rect 5684 4088 5690 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 6840 4128 6868 4168
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 7300 4168 7512 4196
rect 6779 4100 6868 4128
rect 6917 4131 6975 4137
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7300 4128 7328 4168
rect 7484 4137 7512 4168
rect 6963 4100 7328 4128
rect 7377 4131 7435 4137
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 7392 4060 7420 4091
rect 6043 4032 7420 4060
rect 7484 4060 7512 4091
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7616 4100 7665 4128
rect 7616 4088 7622 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 8294 4128 8300 4140
rect 7883 4100 8300 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8846 4128 8852 4140
rect 8619 4100 8852 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8404 4060 8432 4091
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 8662 4060 8668 4072
rect 7484 4032 7604 4060
rect 8404 4032 8668 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 7392 3992 7420 4032
rect 7466 3992 7472 4004
rect 7392 3964 7472 3992
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 7576 3992 7604 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 8754 4020 8760 4072
rect 8812 4020 8818 4072
rect 8772 3992 8800 4020
rect 7576 3964 8800 3992
rect 2590 3884 2596 3936
rect 2648 3884 2654 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4396 3896 4629 3924
rect 4396 3884 4402 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3924 4859 3927
rect 5074 3924 5080 3936
rect 4847 3896 5080 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3924 6883 3927
rect 7374 3924 7380 3936
rect 6871 3896 7380 3924
rect 6871 3893 6883 3896
rect 6825 3887 6883 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2682 3720 2688 3732
rect 2363 3692 2688 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 4154 3680 4160 3732
rect 4212 3680 4218 3732
rect 3973 3655 4031 3661
rect 3973 3621 3985 3655
rect 4019 3621 4031 3655
rect 3973 3615 4031 3621
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 2498 3584 2504 3596
rect 2455 3556 2504 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 2096 3488 2145 3516
rect 2096 3476 2102 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3988 3516 4016 3615
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3584 6147 3587
rect 6730 3584 6736 3596
rect 6135 3556 6736 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 3467 3488 4016 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4580 3488 4905 3516
rect 4580 3476 4586 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5644 3516 5672 3547
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7466 3544 7472 3596
rect 7524 3544 7530 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8352 3556 9229 3584
rect 8352 3544 8358 3556
rect 9217 3553 9229 3556
rect 9263 3553 9275 3587
rect 9217 3547 9275 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9858 3584 9864 3596
rect 9723 3556 9864 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 5132 3488 5672 3516
rect 5132 3476 5138 3488
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 8720 3488 9321 3516
rect 8720 3476 8726 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4125 3451 4183 3457
rect 4125 3448 4137 3451
rect 3844 3420 4137 3448
rect 3844 3408 3850 3420
rect 4125 3417 4137 3420
rect 4171 3417 4183 3451
rect 4125 3411 4183 3417
rect 4341 3451 4399 3457
rect 4341 3417 4353 3451
rect 4387 3448 4399 3451
rect 4430 3448 4436 3460
rect 4387 3420 4436 3448
rect 4387 3417 4399 3420
rect 4341 3411 4399 3417
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 1946 3340 1952 3392
rect 2004 3340 2010 3392
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 3970 3380 3976 3392
rect 3375 3352 3976 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5258 3380 5264 3392
rect 5031 3352 5264 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 8110 3380 8116 3392
rect 7791 3352 8116 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 2498 3136 2504 3188
rect 2556 3136 2562 3188
rect 1486 3068 1492 3120
rect 1544 3108 1550 3120
rect 2516 3108 2544 3136
rect 1544 3080 2452 3108
rect 2516 3080 3188 3108
rect 1544 3068 1550 3080
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2424 3040 2452 3080
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2424 3012 2513 3040
rect 2041 3003 2099 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 1762 2932 1768 2984
rect 1820 2932 1826 2984
rect 2056 2972 2084 3003
rect 2682 3000 2688 3052
rect 2740 3000 2746 3052
rect 3160 3049 3188 3080
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 8812 3012 9873 3040
rect 8812 3000 8818 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 2056 2944 3249 2972
rect 3237 2941 3249 2944
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 11054 2972 11060 2984
rect 10183 2944 11060 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 1765 2635 1823 2641
rect 1765 2632 1777 2635
rect 1728 2604 1777 2632
rect 1728 2592 1734 2604
rect 1765 2601 1777 2604
rect 1811 2632 1823 2635
rect 2682 2632 2688 2644
rect 1811 2604 2688 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 1596 2468 3249 2496
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1596 2437 1624 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 992 2400 1593 2428
rect 992 2388 998 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2004 2400 2329 2428
rect 2004 2388 2010 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9858 2428 9864 2440
rect 9723 2400 9864 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 2222 2320 2228 2372
rect 2280 2360 2286 2372
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 2280 2332 2605 2360
rect 2280 2320 2286 2332
rect 2593 2329 2605 2332
rect 2639 2329 2651 2363
rect 2593 2323 2651 2329
rect 4246 2320 4252 2372
rect 4304 2320 4310 2372
rect 5534 2320 5540 2372
rect 5592 2320 5598 2372
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 6972 2332 7021 2360
rect 6972 2320 6978 2332
rect 7009 2329 7021 2332
rect 7055 2329 7067 2363
rect 7009 2323 7067 2329
rect 8389 2363 8447 2369
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 8662 2360 8668 2372
rect 8435 2332 8668 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 9640 2332 9965 2360
rect 9640 2320 9646 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 9953 2323 10011 2329
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 750 892 756 944
rect 808 932 814 944
rect 1762 932 1768 944
rect 808 904 1768 932
rect 808 892 814 904
rect 1762 892 1768 904
rect 1820 892 1826 944
rect 3694 892 3700 944
rect 3752 932 3758 944
rect 4246 932 4252 944
rect 3752 904 4252 932
rect 3752 892 3758 904
rect 4246 892 4252 904
rect 4304 892 4310 944
rect 8110 892 8116 944
rect 8168 932 8174 944
rect 8662 932 8668 944
rect 8168 904 8668 932
rect 8168 892 8174 904
rect 8662 892 8668 904
rect 8720 892 8726 944
<< via1 >>
rect 2169 15750 2221 15802
rect 2233 15750 2285 15802
rect 2297 15750 2349 15802
rect 2361 15750 2413 15802
rect 2425 15750 2477 15802
rect 4607 15750 4659 15802
rect 4671 15750 4723 15802
rect 4735 15750 4787 15802
rect 4799 15750 4851 15802
rect 4863 15750 4915 15802
rect 7045 15750 7097 15802
rect 7109 15750 7161 15802
rect 7173 15750 7225 15802
rect 7237 15750 7289 15802
rect 7301 15750 7353 15802
rect 9483 15750 9535 15802
rect 9547 15750 9599 15802
rect 9611 15750 9663 15802
rect 9675 15750 9727 15802
rect 9739 15750 9791 15802
rect 940 15444 992 15496
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 5448 15308 5500 15360
rect 3388 15206 3440 15258
rect 3452 15206 3504 15258
rect 3516 15206 3568 15258
rect 3580 15206 3632 15258
rect 3644 15206 3696 15258
rect 5826 15206 5878 15258
rect 5890 15206 5942 15258
rect 5954 15206 6006 15258
rect 6018 15206 6070 15258
rect 6082 15206 6134 15258
rect 8264 15206 8316 15258
rect 8328 15206 8380 15258
rect 8392 15206 8444 15258
rect 8456 15206 8508 15258
rect 8520 15206 8572 15258
rect 10702 15206 10754 15258
rect 10766 15206 10818 15258
rect 10830 15206 10882 15258
rect 10894 15206 10946 15258
rect 10958 15206 11010 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2169 14662 2221 14714
rect 2233 14662 2285 14714
rect 2297 14662 2349 14714
rect 2361 14662 2413 14714
rect 2425 14662 2477 14714
rect 4607 14662 4659 14714
rect 4671 14662 4723 14714
rect 4735 14662 4787 14714
rect 4799 14662 4851 14714
rect 4863 14662 4915 14714
rect 7045 14662 7097 14714
rect 7109 14662 7161 14714
rect 7173 14662 7225 14714
rect 7237 14662 7289 14714
rect 7301 14662 7353 14714
rect 9483 14662 9535 14714
rect 9547 14662 9599 14714
rect 9611 14662 9663 14714
rect 9675 14662 9727 14714
rect 9739 14662 9791 14714
rect 940 14288 992 14340
rect 2688 14288 2740 14340
rect 3388 14118 3440 14170
rect 3452 14118 3504 14170
rect 3516 14118 3568 14170
rect 3580 14118 3632 14170
rect 3644 14118 3696 14170
rect 5826 14118 5878 14170
rect 5890 14118 5942 14170
rect 5954 14118 6006 14170
rect 6018 14118 6070 14170
rect 6082 14118 6134 14170
rect 8264 14118 8316 14170
rect 8328 14118 8380 14170
rect 8392 14118 8444 14170
rect 8456 14118 8508 14170
rect 8520 14118 8572 14170
rect 10702 14118 10754 14170
rect 10766 14118 10818 14170
rect 10830 14118 10882 14170
rect 10894 14118 10946 14170
rect 10958 14118 11010 14170
rect 940 14016 992 14068
rect 2169 13574 2221 13626
rect 2233 13574 2285 13626
rect 2297 13574 2349 13626
rect 2361 13574 2413 13626
rect 2425 13574 2477 13626
rect 4607 13574 4659 13626
rect 4671 13574 4723 13626
rect 4735 13574 4787 13626
rect 4799 13574 4851 13626
rect 4863 13574 4915 13626
rect 7045 13574 7097 13626
rect 7109 13574 7161 13626
rect 7173 13574 7225 13626
rect 7237 13574 7289 13626
rect 7301 13574 7353 13626
rect 9483 13574 9535 13626
rect 9547 13574 9599 13626
rect 9611 13574 9663 13626
rect 9675 13574 9727 13626
rect 9739 13574 9791 13626
rect 3388 13030 3440 13082
rect 3452 13030 3504 13082
rect 3516 13030 3568 13082
rect 3580 13030 3632 13082
rect 3644 13030 3696 13082
rect 5826 13030 5878 13082
rect 5890 13030 5942 13082
rect 5954 13030 6006 13082
rect 6018 13030 6070 13082
rect 6082 13030 6134 13082
rect 8264 13030 8316 13082
rect 8328 13030 8380 13082
rect 8392 13030 8444 13082
rect 8456 13030 8508 13082
rect 8520 13030 8572 13082
rect 10702 13030 10754 13082
rect 10766 13030 10818 13082
rect 10830 13030 10882 13082
rect 10894 13030 10946 13082
rect 10958 13030 11010 13082
rect 2169 12486 2221 12538
rect 2233 12486 2285 12538
rect 2297 12486 2349 12538
rect 2361 12486 2413 12538
rect 2425 12486 2477 12538
rect 4607 12486 4659 12538
rect 4671 12486 4723 12538
rect 4735 12486 4787 12538
rect 4799 12486 4851 12538
rect 4863 12486 4915 12538
rect 7045 12486 7097 12538
rect 7109 12486 7161 12538
rect 7173 12486 7225 12538
rect 7237 12486 7289 12538
rect 7301 12486 7353 12538
rect 9483 12486 9535 12538
rect 9547 12486 9599 12538
rect 9611 12486 9663 12538
rect 9675 12486 9727 12538
rect 9739 12486 9791 12538
rect 940 12112 992 12164
rect 2044 12155 2096 12164
rect 2044 12121 2053 12155
rect 2053 12121 2087 12155
rect 2087 12121 2096 12155
rect 2044 12112 2096 12121
rect 3388 11942 3440 11994
rect 3452 11942 3504 11994
rect 3516 11942 3568 11994
rect 3580 11942 3632 11994
rect 3644 11942 3696 11994
rect 5826 11942 5878 11994
rect 5890 11942 5942 11994
rect 5954 11942 6006 11994
rect 6018 11942 6070 11994
rect 6082 11942 6134 11994
rect 8264 11942 8316 11994
rect 8328 11942 8380 11994
rect 8392 11942 8444 11994
rect 8456 11942 8508 11994
rect 8520 11942 8572 11994
rect 10702 11942 10754 11994
rect 10766 11942 10818 11994
rect 10830 11942 10882 11994
rect 10894 11942 10946 11994
rect 10958 11942 11010 11994
rect 940 11840 992 11892
rect 5448 11840 5500 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 2688 11772 2740 11824
rect 5908 11772 5960 11824
rect 2044 11704 2096 11756
rect 2504 11704 2556 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 6460 11704 6512 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 3240 11500 3292 11552
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 2169 11398 2221 11450
rect 2233 11398 2285 11450
rect 2297 11398 2349 11450
rect 2361 11398 2413 11450
rect 2425 11398 2477 11450
rect 4607 11398 4659 11450
rect 4671 11398 4723 11450
rect 4735 11398 4787 11450
rect 4799 11398 4851 11450
rect 4863 11398 4915 11450
rect 7045 11398 7097 11450
rect 7109 11398 7161 11450
rect 7173 11398 7225 11450
rect 7237 11398 7289 11450
rect 7301 11398 7353 11450
rect 9483 11398 9535 11450
rect 9547 11398 9599 11450
rect 9611 11398 9663 11450
rect 9675 11398 9727 11450
rect 9739 11398 9791 11450
rect 6736 11296 6788 11348
rect 7932 11228 7984 11280
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 4252 11160 4304 11212
rect 1492 11092 1544 11144
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 5632 11160 5684 11212
rect 1860 11024 1912 11076
rect 2504 11024 2556 11076
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 2964 11024 3016 11076
rect 4896 11024 4948 11076
rect 6552 11024 6604 11076
rect 6644 10956 6696 11008
rect 3388 10854 3440 10906
rect 3452 10854 3504 10906
rect 3516 10854 3568 10906
rect 3580 10854 3632 10906
rect 3644 10854 3696 10906
rect 5826 10854 5878 10906
rect 5890 10854 5942 10906
rect 5954 10854 6006 10906
rect 6018 10854 6070 10906
rect 6082 10854 6134 10906
rect 8264 10854 8316 10906
rect 8328 10854 8380 10906
rect 8392 10854 8444 10906
rect 8456 10854 8508 10906
rect 8520 10854 8572 10906
rect 10702 10854 10754 10906
rect 10766 10854 10818 10906
rect 10830 10854 10882 10906
rect 10894 10854 10946 10906
rect 10958 10854 11010 10906
rect 1492 10616 1544 10668
rect 1860 10616 1912 10668
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2688 10616 2740 10668
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 3056 10548 3108 10600
rect 3976 10616 4028 10668
rect 4252 10616 4304 10668
rect 4528 10616 4580 10668
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 6460 10616 6512 10668
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 2688 10480 2740 10532
rect 5540 10548 5592 10600
rect 5448 10480 5500 10532
rect 4068 10412 4120 10464
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 2169 10310 2221 10362
rect 2233 10310 2285 10362
rect 2297 10310 2349 10362
rect 2361 10310 2413 10362
rect 2425 10310 2477 10362
rect 4607 10310 4659 10362
rect 4671 10310 4723 10362
rect 4735 10310 4787 10362
rect 4799 10310 4851 10362
rect 4863 10310 4915 10362
rect 7045 10310 7097 10362
rect 7109 10310 7161 10362
rect 7173 10310 7225 10362
rect 7237 10310 7289 10362
rect 7301 10310 7353 10362
rect 9483 10310 9535 10362
rect 9547 10310 9599 10362
rect 9611 10310 9663 10362
rect 9675 10310 9727 10362
rect 9739 10310 9791 10362
rect 3056 10208 3108 10260
rect 3240 10140 3292 10192
rect 940 10004 992 10056
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3976 10047 4028 10056
rect 1492 9936 1544 9988
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4528 10208 4580 10260
rect 5632 10072 5684 10124
rect 2964 9868 3016 9920
rect 3884 9868 3936 9920
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 7380 9052 7432 9104
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 1860 8848 1912 8900
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6920 8916 6972 8968
rect 7380 8916 7432 8968
rect 8852 8916 8904 8968
rect 940 8780 992 8832
rect 8668 8780 8720 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 1860 8551 1912 8560
rect 1860 8517 1869 8551
rect 1869 8517 1903 8551
rect 1903 8517 1912 8551
rect 1860 8508 1912 8517
rect 4988 8576 5040 8628
rect 940 8440 992 8492
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2596 8440 2648 8492
rect 4436 8508 4488 8560
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 4068 8304 4120 8356
rect 3884 8236 3936 8288
rect 5264 8304 5316 8356
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 4068 8032 4120 8084
rect 1492 7896 1544 7948
rect 2688 7896 2740 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 1676 7760 1728 7812
rect 2596 7828 2648 7880
rect 3884 7828 3936 7880
rect 4068 7828 4120 7880
rect 2964 7803 3016 7812
rect 2964 7769 2973 7803
rect 2973 7769 3007 7803
rect 3007 7769 3016 7803
rect 2964 7760 3016 7769
rect 3792 7760 3844 7812
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4988 7760 5040 7812
rect 4712 7692 4764 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 4436 7488 4488 7540
rect 1584 7420 1636 7472
rect 1676 7352 1728 7404
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2504 7352 2556 7404
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3884 7463 3936 7472
rect 3884 7429 3893 7463
rect 3893 7429 3927 7463
rect 3927 7429 3936 7463
rect 3884 7420 3936 7429
rect 4528 7420 4580 7472
rect 3792 7352 3844 7404
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4436 7352 4488 7404
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 5448 7463 5500 7472
rect 5448 7429 5457 7463
rect 5457 7429 5491 7463
rect 5491 7429 5500 7463
rect 5448 7420 5500 7429
rect 5632 7463 5684 7472
rect 5632 7429 5641 7463
rect 5641 7429 5675 7463
rect 5675 7429 5684 7463
rect 5632 7420 5684 7429
rect 4988 7352 5040 7404
rect 6828 7352 6880 7404
rect 7380 7352 7432 7404
rect 6368 7284 6420 7336
rect 6920 7216 6972 7268
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4988 7148 5040 7200
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 2044 6944 2096 6996
rect 2872 6944 2924 6996
rect 6552 6944 6604 6996
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 7104 6808 7156 6860
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 6920 6740 6972 6792
rect 5080 6604 5132 6656
rect 7012 6604 7064 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 7104 6171 7156 6180
rect 7104 6137 7113 6171
rect 7113 6137 7147 6171
rect 7147 6137 7156 6171
rect 7104 6128 7156 6137
rect 940 6060 992 6112
rect 1860 6060 1912 6112
rect 5632 6060 5684 6112
rect 7564 6060 7616 6112
rect 8760 6060 8812 6112
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 4988 5856 5040 5908
rect 2688 5720 2740 5772
rect 940 5652 992 5704
rect 3056 5652 3108 5704
rect 5080 5584 5132 5636
rect 5264 5584 5316 5636
rect 2872 5516 2924 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 2504 5312 2556 5364
rect 1584 5176 1636 5228
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2872 5244 2924 5296
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 1492 5108 1544 5160
rect 3056 5108 3108 5160
rect 3792 4972 3844 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 4528 4743 4580 4752
rect 4528 4709 4537 4743
rect 4537 4709 4571 4743
rect 4571 4709 4580 4743
rect 4528 4700 4580 4709
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 5540 4632 5592 4684
rect 1492 4564 1544 4616
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 2780 4564 2832 4573
rect 3056 4564 3108 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 1676 4496 1728 4548
rect 4068 4496 4120 4548
rect 2044 4428 2096 4480
rect 2596 4428 2648 4480
rect 2780 4428 2832 4480
rect 5724 4428 5776 4480
rect 7196 4428 7248 4480
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1768 4224 1820 4276
rect 4252 4224 4304 4276
rect 5632 4267 5684 4276
rect 5632 4233 5641 4267
rect 5641 4233 5675 4267
rect 5675 4233 5684 4267
rect 5632 4224 5684 4233
rect 2504 4156 2556 4208
rect 2688 4156 2740 4208
rect 3332 4156 3384 4208
rect 4068 4156 4120 4208
rect 940 4088 992 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2780 4088 2832 4140
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 4160 4088 4212 4140
rect 3332 3995 3384 4004
rect 3332 3961 3341 3995
rect 3341 3961 3375 3995
rect 3375 3961 3384 3995
rect 3332 3952 3384 3961
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 4436 3952 4488 4004
rect 5632 4088 5684 4140
rect 7196 4156 7248 4208
rect 7564 4088 7616 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8852 4088 8904 4140
rect 7472 3952 7524 4004
rect 8668 4020 8720 4072
rect 8760 4020 8812 4072
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 4344 3884 4396 3936
rect 5080 3884 5132 3936
rect 7380 3884 7432 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 2688 3680 2740 3732
rect 4160 3723 4212 3732
rect 4160 3689 4169 3723
rect 4169 3689 4203 3723
rect 4203 3689 4212 3723
rect 4160 3680 4212 3689
rect 2504 3544 2556 3596
rect 2044 3476 2096 3528
rect 3332 3476 3384 3528
rect 4528 3476 4580 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 6736 3544 6788 3596
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 8300 3544 8352 3596
rect 9864 3544 9916 3596
rect 5080 3476 5132 3485
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 8668 3476 8720 3528
rect 3792 3408 3844 3460
rect 4436 3408 4488 3460
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 3976 3340 4028 3392
rect 5264 3340 5316 3392
rect 8116 3340 8168 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 1492 3068 1544 3120
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 8760 3000 8812 3052
rect 11060 2932 11112 2984
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 1676 2592 1728 2644
rect 2688 2592 2740 2644
rect 940 2388 992 2440
rect 1952 2388 2004 2440
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9864 2388 9916 2440
rect 2228 2320 2280 2372
rect 4252 2363 4304 2372
rect 4252 2329 4261 2363
rect 4261 2329 4295 2363
rect 4295 2329 4304 2363
rect 4252 2320 4304 2329
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 6920 2320 6972 2372
rect 8668 2320 8720 2372
rect 9588 2320 9640 2372
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 756 892 808 944
rect 1768 892 1820 944
rect 3700 892 3752 944
rect 4252 892 4304 944
rect 8116 892 8168 944
rect 8668 892 8720 944
<< metal2 >>
rect 938 16552 994 16561
rect 938 16487 994 16496
rect 952 15502 980 16487
rect 2169 15804 2477 15813
rect 2169 15802 2175 15804
rect 2231 15802 2255 15804
rect 2311 15802 2335 15804
rect 2391 15802 2415 15804
rect 2471 15802 2477 15804
rect 2231 15750 2233 15802
rect 2413 15750 2415 15802
rect 2169 15748 2175 15750
rect 2231 15748 2255 15750
rect 2311 15748 2335 15750
rect 2391 15748 2415 15750
rect 2471 15748 2477 15750
rect 2169 15739 2477 15748
rect 4607 15804 4915 15813
rect 4607 15802 4613 15804
rect 4669 15802 4693 15804
rect 4749 15802 4773 15804
rect 4829 15802 4853 15804
rect 4909 15802 4915 15804
rect 4669 15750 4671 15802
rect 4851 15750 4853 15802
rect 4607 15748 4613 15750
rect 4669 15748 4693 15750
rect 4749 15748 4773 15750
rect 4829 15748 4853 15750
rect 4909 15748 4915 15750
rect 4607 15739 4915 15748
rect 7045 15804 7353 15813
rect 7045 15802 7051 15804
rect 7107 15802 7131 15804
rect 7187 15802 7211 15804
rect 7267 15802 7291 15804
rect 7347 15802 7353 15804
rect 7107 15750 7109 15802
rect 7289 15750 7291 15802
rect 7045 15748 7051 15750
rect 7107 15748 7131 15750
rect 7187 15748 7211 15750
rect 7267 15748 7291 15750
rect 7347 15748 7353 15750
rect 7045 15739 7353 15748
rect 9483 15804 9791 15813
rect 9483 15802 9489 15804
rect 9545 15802 9569 15804
rect 9625 15802 9649 15804
rect 9705 15802 9729 15804
rect 9785 15802 9791 15804
rect 9545 15750 9547 15802
rect 9727 15750 9729 15802
rect 9483 15748 9489 15750
rect 9545 15748 9569 15750
rect 9625 15748 9649 15750
rect 9705 15748 9729 15750
rect 9785 15748 9791 15750
rect 9483 15739 9791 15748
rect 940 15496 992 15502
rect 940 15438 992 15444
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15162 1624 15438
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 3388 15260 3696 15269
rect 3388 15258 3394 15260
rect 3450 15258 3474 15260
rect 3530 15258 3554 15260
rect 3610 15258 3634 15260
rect 3690 15258 3696 15260
rect 3450 15206 3452 15258
rect 3632 15206 3634 15258
rect 3388 15204 3394 15206
rect 3450 15204 3474 15206
rect 3530 15204 3554 15206
rect 3610 15204 3634 15206
rect 3690 15204 3696 15206
rect 3388 15195 3696 15204
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 2169 14716 2477 14725
rect 2169 14714 2175 14716
rect 2231 14714 2255 14716
rect 2311 14714 2335 14716
rect 2391 14714 2415 14716
rect 2471 14714 2477 14716
rect 2231 14662 2233 14714
rect 2413 14662 2415 14714
rect 2169 14660 2175 14662
rect 2231 14660 2255 14662
rect 2311 14660 2335 14662
rect 2391 14660 2415 14662
rect 2471 14660 2477 14662
rect 2169 14651 2477 14660
rect 4607 14716 4915 14725
rect 4607 14714 4613 14716
rect 4669 14714 4693 14716
rect 4749 14714 4773 14716
rect 4829 14714 4853 14716
rect 4909 14714 4915 14716
rect 4669 14662 4671 14714
rect 4851 14662 4853 14714
rect 4607 14660 4613 14662
rect 4669 14660 4693 14662
rect 4749 14660 4773 14662
rect 4829 14660 4853 14662
rect 4909 14660 4915 14662
rect 4607 14651 4915 14660
rect 938 14376 994 14385
rect 938 14311 940 14320
rect 992 14311 994 14320
rect 2688 14340 2740 14346
rect 940 14282 992 14288
rect 2688 14282 2740 14288
rect 952 14074 980 14282
rect 940 14068 992 14074
rect 940 14010 992 14016
rect 2169 13628 2477 13637
rect 2169 13626 2175 13628
rect 2231 13626 2255 13628
rect 2311 13626 2335 13628
rect 2391 13626 2415 13628
rect 2471 13626 2477 13628
rect 2231 13574 2233 13626
rect 2413 13574 2415 13626
rect 2169 13572 2175 13574
rect 2231 13572 2255 13574
rect 2311 13572 2335 13574
rect 2391 13572 2415 13574
rect 2471 13572 2477 13574
rect 2169 13563 2477 13572
rect 2169 12540 2477 12549
rect 2169 12538 2175 12540
rect 2231 12538 2255 12540
rect 2311 12538 2335 12540
rect 2391 12538 2415 12540
rect 2471 12538 2477 12540
rect 2231 12486 2233 12538
rect 2413 12486 2415 12538
rect 2169 12484 2175 12486
rect 2231 12484 2255 12486
rect 2311 12484 2335 12486
rect 2391 12484 2415 12486
rect 2471 12484 2477 12486
rect 2169 12475 2477 12484
rect 938 12200 994 12209
rect 938 12135 940 12144
rect 992 12135 994 12144
rect 2044 12164 2096 12170
rect 940 12106 992 12112
rect 2044 12106 2096 12112
rect 952 11898 980 12106
rect 940 11892 992 11898
rect 940 11834 992 11840
rect 2056 11762 2084 12106
rect 2700 11830 2728 14282
rect 3388 14172 3696 14181
rect 3388 14170 3394 14172
rect 3450 14170 3474 14172
rect 3530 14170 3554 14172
rect 3610 14170 3634 14172
rect 3690 14170 3696 14172
rect 3450 14118 3452 14170
rect 3632 14118 3634 14170
rect 3388 14116 3394 14118
rect 3450 14116 3474 14118
rect 3530 14116 3554 14118
rect 3610 14116 3634 14118
rect 3690 14116 3696 14118
rect 3388 14107 3696 14116
rect 4607 13628 4915 13637
rect 4607 13626 4613 13628
rect 4669 13626 4693 13628
rect 4749 13626 4773 13628
rect 4829 13626 4853 13628
rect 4909 13626 4915 13628
rect 4669 13574 4671 13626
rect 4851 13574 4853 13626
rect 4607 13572 4613 13574
rect 4669 13572 4693 13574
rect 4749 13572 4773 13574
rect 4829 13572 4853 13574
rect 4909 13572 4915 13574
rect 4607 13563 4915 13572
rect 3388 13084 3696 13093
rect 3388 13082 3394 13084
rect 3450 13082 3474 13084
rect 3530 13082 3554 13084
rect 3610 13082 3634 13084
rect 3690 13082 3696 13084
rect 3450 13030 3452 13082
rect 3632 13030 3634 13082
rect 3388 13028 3394 13030
rect 3450 13028 3474 13030
rect 3530 13028 3554 13030
rect 3610 13028 3634 13030
rect 3690 13028 3696 13030
rect 3388 13019 3696 13028
rect 4607 12540 4915 12549
rect 4607 12538 4613 12540
rect 4669 12538 4693 12540
rect 4749 12538 4773 12540
rect 4829 12538 4853 12540
rect 4909 12538 4915 12540
rect 4669 12486 4671 12538
rect 4851 12486 4853 12538
rect 4607 12484 4613 12486
rect 4669 12484 4693 12486
rect 4749 12484 4773 12486
rect 4829 12484 4853 12486
rect 4909 12484 4915 12486
rect 4607 12475 4915 12484
rect 3388 11996 3696 12005
rect 3388 11994 3394 11996
rect 3450 11994 3474 11996
rect 3530 11994 3554 11996
rect 3610 11994 3634 11996
rect 3690 11994 3696 11996
rect 3450 11942 3452 11994
rect 3632 11942 3634 11994
rect 3388 11940 3394 11942
rect 3450 11940 3474 11942
rect 3530 11940 3554 11942
rect 3610 11940 3634 11942
rect 3690 11940 3696 11942
rect 3388 11931 3696 11940
rect 5460 11914 5488 15302
rect 5826 15260 6134 15269
rect 5826 15258 5832 15260
rect 5888 15258 5912 15260
rect 5968 15258 5992 15260
rect 6048 15258 6072 15260
rect 6128 15258 6134 15260
rect 5888 15206 5890 15258
rect 6070 15206 6072 15258
rect 5826 15204 5832 15206
rect 5888 15204 5912 15206
rect 5968 15204 5992 15206
rect 6048 15204 6072 15206
rect 6128 15204 6134 15206
rect 5826 15195 6134 15204
rect 8264 15260 8572 15269
rect 8264 15258 8270 15260
rect 8326 15258 8350 15260
rect 8406 15258 8430 15260
rect 8486 15258 8510 15260
rect 8566 15258 8572 15260
rect 8326 15206 8328 15258
rect 8508 15206 8510 15258
rect 8264 15204 8270 15206
rect 8326 15204 8350 15206
rect 8406 15204 8430 15206
rect 8486 15204 8510 15206
rect 8566 15204 8572 15206
rect 8264 15195 8572 15204
rect 10702 15260 11010 15269
rect 10702 15258 10708 15260
rect 10764 15258 10788 15260
rect 10844 15258 10868 15260
rect 10924 15258 10948 15260
rect 11004 15258 11010 15260
rect 10764 15206 10766 15258
rect 10946 15206 10948 15258
rect 10702 15204 10708 15206
rect 10764 15204 10788 15206
rect 10844 15204 10868 15206
rect 10924 15204 10948 15206
rect 11004 15204 11010 15206
rect 10702 15195 11010 15204
rect 7045 14716 7353 14725
rect 7045 14714 7051 14716
rect 7107 14714 7131 14716
rect 7187 14714 7211 14716
rect 7267 14714 7291 14716
rect 7347 14714 7353 14716
rect 7107 14662 7109 14714
rect 7289 14662 7291 14714
rect 7045 14660 7051 14662
rect 7107 14660 7131 14662
rect 7187 14660 7211 14662
rect 7267 14660 7291 14662
rect 7347 14660 7353 14662
rect 7045 14651 7353 14660
rect 9483 14716 9791 14725
rect 9483 14714 9489 14716
rect 9545 14714 9569 14716
rect 9625 14714 9649 14716
rect 9705 14714 9729 14716
rect 9785 14714 9791 14716
rect 9545 14662 9547 14714
rect 9727 14662 9729 14714
rect 9483 14660 9489 14662
rect 9545 14660 9569 14662
rect 9625 14660 9649 14662
rect 9705 14660 9729 14662
rect 9785 14660 9791 14662
rect 9483 14651 9791 14660
rect 5826 14172 6134 14181
rect 5826 14170 5832 14172
rect 5888 14170 5912 14172
rect 5968 14170 5992 14172
rect 6048 14170 6072 14172
rect 6128 14170 6134 14172
rect 5888 14118 5890 14170
rect 6070 14118 6072 14170
rect 5826 14116 5832 14118
rect 5888 14116 5912 14118
rect 5968 14116 5992 14118
rect 6048 14116 6072 14118
rect 6128 14116 6134 14118
rect 5826 14107 6134 14116
rect 8264 14172 8572 14181
rect 8264 14170 8270 14172
rect 8326 14170 8350 14172
rect 8406 14170 8430 14172
rect 8486 14170 8510 14172
rect 8566 14170 8572 14172
rect 8326 14118 8328 14170
rect 8508 14118 8510 14170
rect 8264 14116 8270 14118
rect 8326 14116 8350 14118
rect 8406 14116 8430 14118
rect 8486 14116 8510 14118
rect 8566 14116 8572 14118
rect 8264 14107 8572 14116
rect 10702 14172 11010 14181
rect 10702 14170 10708 14172
rect 10764 14170 10788 14172
rect 10844 14170 10868 14172
rect 10924 14170 10948 14172
rect 11004 14170 11010 14172
rect 10764 14118 10766 14170
rect 10946 14118 10948 14170
rect 10702 14116 10708 14118
rect 10764 14116 10788 14118
rect 10844 14116 10868 14118
rect 10924 14116 10948 14118
rect 11004 14116 11010 14118
rect 10702 14107 11010 14116
rect 7045 13628 7353 13637
rect 7045 13626 7051 13628
rect 7107 13626 7131 13628
rect 7187 13626 7211 13628
rect 7267 13626 7291 13628
rect 7347 13626 7353 13628
rect 7107 13574 7109 13626
rect 7289 13574 7291 13626
rect 7045 13572 7051 13574
rect 7107 13572 7131 13574
rect 7187 13572 7211 13574
rect 7267 13572 7291 13574
rect 7347 13572 7353 13574
rect 7045 13563 7353 13572
rect 9483 13628 9791 13637
rect 9483 13626 9489 13628
rect 9545 13626 9569 13628
rect 9625 13626 9649 13628
rect 9705 13626 9729 13628
rect 9785 13626 9791 13628
rect 9545 13574 9547 13626
rect 9727 13574 9729 13626
rect 9483 13572 9489 13574
rect 9545 13572 9569 13574
rect 9625 13572 9649 13574
rect 9705 13572 9729 13574
rect 9785 13572 9791 13574
rect 9483 13563 9791 13572
rect 5826 13084 6134 13093
rect 5826 13082 5832 13084
rect 5888 13082 5912 13084
rect 5968 13082 5992 13084
rect 6048 13082 6072 13084
rect 6128 13082 6134 13084
rect 5888 13030 5890 13082
rect 6070 13030 6072 13082
rect 5826 13028 5832 13030
rect 5888 13028 5912 13030
rect 5968 13028 5992 13030
rect 6048 13028 6072 13030
rect 6128 13028 6134 13030
rect 5826 13019 6134 13028
rect 8264 13084 8572 13093
rect 8264 13082 8270 13084
rect 8326 13082 8350 13084
rect 8406 13082 8430 13084
rect 8486 13082 8510 13084
rect 8566 13082 8572 13084
rect 8326 13030 8328 13082
rect 8508 13030 8510 13082
rect 8264 13028 8270 13030
rect 8326 13028 8350 13030
rect 8406 13028 8430 13030
rect 8486 13028 8510 13030
rect 8566 13028 8572 13030
rect 8264 13019 8572 13028
rect 10702 13084 11010 13093
rect 10702 13082 10708 13084
rect 10764 13082 10788 13084
rect 10844 13082 10868 13084
rect 10924 13082 10948 13084
rect 11004 13082 11010 13084
rect 10764 13030 10766 13082
rect 10946 13030 10948 13082
rect 10702 13028 10708 13030
rect 10764 13028 10788 13030
rect 10844 13028 10868 13030
rect 10924 13028 10948 13030
rect 11004 13028 11010 13030
rect 10702 13019 11010 13028
rect 7045 12540 7353 12549
rect 7045 12538 7051 12540
rect 7107 12538 7131 12540
rect 7187 12538 7211 12540
rect 7267 12538 7291 12540
rect 7347 12538 7353 12540
rect 7107 12486 7109 12538
rect 7289 12486 7291 12538
rect 7045 12484 7051 12486
rect 7107 12484 7131 12486
rect 7187 12484 7211 12486
rect 7267 12484 7291 12486
rect 7347 12484 7353 12486
rect 7045 12475 7353 12484
rect 9483 12540 9791 12549
rect 9483 12538 9489 12540
rect 9545 12538 9569 12540
rect 9625 12538 9649 12540
rect 9705 12538 9729 12540
rect 9785 12538 9791 12540
rect 9545 12486 9547 12538
rect 9727 12486 9729 12538
rect 9483 12484 9489 12486
rect 9545 12484 9569 12486
rect 9625 12484 9649 12486
rect 9705 12484 9729 12486
rect 9785 12484 9791 12486
rect 9483 12475 9791 12484
rect 5826 11996 6134 12005
rect 5826 11994 5832 11996
rect 5888 11994 5912 11996
rect 5968 11994 5992 11996
rect 6048 11994 6072 11996
rect 6128 11994 6134 11996
rect 5888 11942 5890 11994
rect 6070 11942 6072 11994
rect 5826 11940 5832 11942
rect 5888 11940 5912 11942
rect 5968 11940 5992 11942
rect 6048 11940 6072 11942
rect 6128 11940 6134 11942
rect 5826 11931 6134 11940
rect 8264 11996 8572 12005
rect 8264 11994 8270 11996
rect 8326 11994 8350 11996
rect 8406 11994 8430 11996
rect 8486 11994 8510 11996
rect 8566 11994 8572 11996
rect 8326 11942 8328 11994
rect 8508 11942 8510 11994
rect 8264 11940 8270 11942
rect 8326 11940 8350 11942
rect 8406 11940 8430 11942
rect 8486 11940 8510 11942
rect 8566 11940 8572 11942
rect 8264 11931 8572 11940
rect 10702 11996 11010 12005
rect 10702 11994 10708 11996
rect 10764 11994 10788 11996
rect 10844 11994 10868 11996
rect 10924 11994 10948 11996
rect 11004 11994 11010 11996
rect 10764 11942 10766 11994
rect 10946 11942 10948 11994
rect 10702 11940 10708 11942
rect 10764 11940 10788 11942
rect 10844 11940 10868 11942
rect 10924 11940 10948 11942
rect 11004 11940 11010 11942
rect 10702 11931 11010 11940
rect 5368 11898 5488 11914
rect 5368 11892 5500 11898
rect 5368 11886 5448 11892
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2056 11150 2084 11698
rect 2169 11452 2477 11461
rect 2169 11450 2175 11452
rect 2231 11450 2255 11452
rect 2311 11450 2335 11452
rect 2391 11450 2415 11452
rect 2471 11450 2477 11452
rect 2231 11398 2233 11450
rect 2413 11398 2415 11450
rect 2169 11396 2175 11398
rect 2231 11396 2255 11398
rect 2311 11396 2335 11398
rect 2391 11396 2415 11398
rect 2471 11396 2477 11398
rect 2169 11387 2477 11396
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1504 10674 1532 11086
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10674 1900 11018
rect 2056 10674 2084 11086
rect 2516 11082 2544 11698
rect 2700 11234 2728 11766
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 2608 11206 2728 11234
rect 2964 11212 3016 11218
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 940 10056 992 10062
rect 938 10024 940 10033
rect 992 10024 994 10033
rect 1504 9994 1532 10610
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 938 9959 994 9968
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 952 8498 980 8774
rect 940 8492 992 8498
rect 940 8434 992 8440
rect 952 7857 980 8434
rect 1504 7954 1532 9930
rect 1596 9722 1624 9998
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1872 8906 1900 10610
rect 2056 10010 2084 10610
rect 2169 10364 2477 10373
rect 2169 10362 2175 10364
rect 2231 10362 2255 10364
rect 2311 10362 2335 10364
rect 2391 10362 2415 10364
rect 2471 10362 2477 10364
rect 2231 10310 2233 10362
rect 2413 10310 2415 10362
rect 2169 10308 2175 10310
rect 2231 10308 2255 10310
rect 2311 10308 2335 10310
rect 2391 10308 2415 10310
rect 2471 10308 2477 10310
rect 2169 10299 2477 10308
rect 2608 10282 2636 11206
rect 2964 11154 3016 11160
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 10674 2728 11086
rect 2976 11082 3004 11154
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10538 2728 10610
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 1964 9982 2084 10010
rect 2516 10254 2636 10282
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8566 1900 8842
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 938 7848 994 7857
rect 938 7783 994 7792
rect 940 6112 992 6118
rect 940 6054 992 6060
rect 952 5710 980 6054
rect 940 5704 992 5710
rect 938 5672 940 5681
rect 992 5672 994 5681
rect 938 5607 994 5616
rect 1504 5166 1532 7890
rect 1964 7886 1992 9982
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2516 8498 2544 10254
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1596 7478 1624 7822
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1596 5234 1624 7414
rect 1688 7410 1716 7754
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1504 4622 1532 5102
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3505 980 4082
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 1504 3126 1532 4558
rect 1688 4554 1716 7346
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1780 4622 1808 5170
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1492 3120 1544 3126
rect 1492 3062 1544 3068
rect 1688 2650 1716 4490
rect 1780 4282 1808 4558
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1872 4146 1900 6054
rect 1964 5234 1992 7822
rect 2516 7410 2544 8434
rect 2608 7886 2636 8434
rect 2700 7954 2728 10474
rect 2976 10062 3004 11018
rect 3252 10674 3280 11494
rect 4607 11452 4915 11461
rect 4607 11450 4613 11452
rect 4669 11450 4693 11452
rect 4749 11450 4773 11452
rect 4829 11450 4853 11452
rect 4909 11450 4915 11452
rect 4669 11398 4671 11450
rect 4851 11398 4853 11450
rect 4607 11396 4613 11398
rect 4669 11396 4693 11398
rect 4749 11396 4773 11398
rect 4829 11396 4853 11398
rect 4909 11396 4915 11398
rect 4607 11387 4915 11396
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 3388 10908 3696 10917
rect 3388 10906 3394 10908
rect 3450 10906 3474 10908
rect 3530 10906 3554 10908
rect 3610 10906 3634 10908
rect 3690 10906 3696 10908
rect 3450 10854 3452 10906
rect 3632 10854 3634 10906
rect 3388 10852 3394 10854
rect 3450 10852 3474 10854
rect 3530 10852 3554 10854
rect 3610 10852 3634 10854
rect 3690 10852 3696 10854
rect 3388 10843 3696 10852
rect 4264 10674 4292 11154
rect 5368 11150 5396 11886
rect 5448 11834 5500 11840
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11150 5488 11698
rect 5644 11218 5672 11834
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5920 11150 5948 11766
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5448 11144 5500 11150
rect 5908 11144 5960 11150
rect 5448 11086 5500 11092
rect 5736 11092 5908 11098
rect 5736 11086 5960 11092
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10674 4936 11018
rect 5460 10962 5488 11086
rect 5736 11070 5948 11086
rect 5460 10934 5580 10962
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3068 10062 3096 10202
rect 3252 10198 3280 10610
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3988 10062 4016 10610
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2056 7002 2084 7346
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2700 5778 2728 7890
rect 2976 7818 3004 9862
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3896 8294 3924 9862
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7886 3924 8230
rect 3988 7970 4016 8366
rect 4080 8362 4108 10406
rect 4540 10266 4568 10610
rect 5552 10606 5580 10934
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 4607 10364 4915 10373
rect 4607 10362 4613 10364
rect 4669 10362 4693 10364
rect 4749 10362 4773 10364
rect 4829 10362 4853 10364
rect 4909 10362 4915 10364
rect 4669 10310 4671 10362
rect 4851 10310 4853 10362
rect 4607 10308 4613 10310
rect 4669 10308 4693 10310
rect 4749 10308 4773 10310
rect 4829 10308 4853 10310
rect 4909 10308 4915 10310
rect 4607 10299 4915 10308
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 8090 4108 8298
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3988 7942 4108 7970
rect 4080 7886 4108 7942
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 7002 2912 7346
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 5658 2728 5714
rect 2700 5630 2820 5658
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4622 1992 5170
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2056 3534 2084 4422
rect 2516 4214 2544 5306
rect 2792 4622 2820 5630
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5302 2912 5510
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2976 5234 3004 7754
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3804 7410 3832 7754
rect 3896 7478 3924 7822
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4080 7410 4108 7822
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3068 5166 3096 5646
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4622 3096 5102
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2516 3602 2544 4014
rect 2608 3942 2636 4422
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2700 3738 2728 4150
rect 2792 4146 2820 4422
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3344 4010 3372 4150
rect 3804 4078 3832 4966
rect 4264 4622 4292 7142
rect 4356 4622 4384 7890
rect 4448 7546 4476 8502
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7478 4568 7822
rect 5000 7818 5028 8570
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4724 7410 4752 7686
rect 5000 7410 5028 7754
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4214 4108 4490
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 952 1329 980 2382
rect 938 1320 994 1329
rect 938 1255 994 1264
rect 1780 950 1808 2926
rect 1964 2446 1992 3334
rect 2516 3194 2544 3538
rect 3344 3534 3372 3946
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3804 3466 3832 4014
rect 4172 3738 4200 4082
rect 4356 3942 4384 4558
rect 4448 4010 4476 7346
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5000 6322 5028 7142
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6458 5120 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5000 5914 5028 6258
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5642 5120 6394
rect 5276 6322 5304 8298
rect 5460 7478 5488 10474
rect 5552 8974 5580 10542
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5644 7478 5672 10066
rect 5736 8974 5764 11070
rect 5826 10908 6134 10917
rect 5826 10906 5832 10908
rect 5888 10906 5912 10908
rect 5968 10906 5992 10908
rect 6048 10906 6072 10908
rect 6128 10906 6134 10908
rect 5888 10854 5890 10906
rect 6070 10854 6072 10906
rect 5826 10852 5832 10854
rect 5888 10852 5912 10854
rect 5968 10852 5992 10854
rect 6048 10852 6072 10854
rect 6128 10852 6134 10854
rect 5826 10843 6134 10852
rect 6472 10674 6500 11698
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 11218 6592 11494
rect 6748 11354 6776 11698
rect 7045 11452 7353 11461
rect 7045 11450 7051 11452
rect 7107 11450 7131 11452
rect 7187 11450 7211 11452
rect 7267 11450 7291 11452
rect 7347 11450 7353 11452
rect 7107 11398 7109 11450
rect 7289 11398 7291 11450
rect 7045 11396 7051 11398
rect 7107 11396 7131 11398
rect 7187 11396 7211 11398
rect 7267 11396 7291 11398
rect 7347 11396 7353 11398
rect 7045 11387 7353 11396
rect 9483 11452 9791 11461
rect 9483 11450 9489 11452
rect 9545 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9791 11452
rect 9545 11398 9547 11450
rect 9727 11398 9729 11450
rect 9483 11396 9489 11398
rect 9545 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9791 11398
rect 9483 11387 9791 11396
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6564 8974 6592 11018
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10674 6684 10950
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6748 10470 6776 11290
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 8974 6960 10406
rect 7045 10364 7353 10373
rect 7045 10362 7051 10364
rect 7107 10362 7131 10364
rect 7187 10362 7211 10364
rect 7267 10362 7291 10364
rect 7347 10362 7353 10364
rect 7107 10310 7109 10362
rect 7289 10310 7291 10362
rect 7045 10308 7051 10310
rect 7107 10308 7131 10310
rect 7187 10308 7211 10310
rect 7267 10308 7291 10310
rect 7347 10308 7353 10310
rect 7045 10299 7353 10308
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7392 8974 7420 9046
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5460 6914 5488 7414
rect 5460 6886 5580 6914
rect 5552 6798 5580 6886
rect 5644 6798 5672 7414
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 6798 6408 7278
rect 6564 7002 6592 8910
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7392 7410 7420 8910
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6840 6798 6868 7346
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6932 6798 6960 7210
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 7024 6322 7052 6598
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 5276 5642 5304 6258
rect 7116 6186 7144 6802
rect 7944 6322 7972 11222
rect 8264 10908 8572 10917
rect 8264 10906 8270 10908
rect 8326 10906 8350 10908
rect 8406 10906 8430 10908
rect 8486 10906 8510 10908
rect 8566 10906 8572 10908
rect 8326 10854 8328 10906
rect 8508 10854 8510 10906
rect 8264 10852 8270 10854
rect 8326 10852 8350 10854
rect 8406 10852 8430 10854
rect 8486 10852 8510 10854
rect 8566 10852 8572 10854
rect 8264 10843 8572 10852
rect 10702 10908 11010 10917
rect 10702 10906 10708 10908
rect 10764 10906 10788 10908
rect 10844 10906 10868 10908
rect 10924 10906 10948 10908
rect 11004 10906 11010 10908
rect 10764 10854 10766 10906
rect 10946 10854 10948 10906
rect 10702 10852 10708 10854
rect 10764 10852 10788 10854
rect 10844 10852 10868 10854
rect 10924 10852 10948 10854
rect 11004 10852 11010 10854
rect 10702 10843 11010 10852
rect 9483 10364 9791 10373
rect 9483 10362 9489 10364
rect 9545 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9791 10364
rect 9545 10310 9547 10362
rect 9727 10310 9729 10362
rect 9483 10308 9489 10310
rect 9545 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9791 10310
rect 9483 10299 9791 10308
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4448 3466 4476 3946
rect 4540 3534 4568 4694
rect 5552 4690 5580 5510
rect 5644 4758 5672 6054
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4162 5580 4626
rect 5644 4282 5672 4694
rect 7576 4622 7604 6054
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5552 4146 5672 4162
rect 5552 4140 5684 4146
rect 5552 4134 5632 4140
rect 5632 4082 5684 4088
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 5092 3534 5120 3878
rect 5736 3534 5764 4422
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 7208 4214 7236 4422
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7576 4146 7604 4558
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2700 2650 2728 2994
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 3988 2446 4016 3334
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 5276 2446 5304 3334
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 6748 2446 6776 3538
rect 7392 3534 7420 3878
rect 7484 3602 7512 3946
rect 8312 3602 8340 4082
rect 8680 4078 8708 8774
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 4078 8800 6054
rect 8864 4146 8892 8910
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8680 3534 8708 4014
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 8128 2446 8156 3334
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8772 3058 8800 3878
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9876 2446 9904 3538
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 756 944 808 950
rect 756 886 808 892
rect 1768 944 1820 950
rect 1768 886 1820 892
rect 768 800 796 886
rect 2240 800 2268 2314
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 4264 950 4292 2314
rect 3700 944 3752 950
rect 3700 886 3752 892
rect 4252 944 4304 950
rect 5552 898 5580 2314
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6932 898 6960 2314
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8680 950 8708 2314
rect 4252 886 4304 892
rect 3712 800 3740 886
rect 5184 870 5580 898
rect 6656 870 6960 898
rect 8116 944 8168 950
rect 8116 886 8168 892
rect 8668 944 8720 950
rect 8668 886 8720 892
rect 5184 800 5212 870
rect 6656 800 6684 870
rect 8128 800 8156 886
rect 9600 800 9628 2314
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 11072 800 11100 2926
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
<< via2 >>
rect 938 16496 994 16552
rect 2175 15802 2231 15804
rect 2255 15802 2311 15804
rect 2335 15802 2391 15804
rect 2415 15802 2471 15804
rect 2175 15750 2221 15802
rect 2221 15750 2231 15802
rect 2255 15750 2285 15802
rect 2285 15750 2297 15802
rect 2297 15750 2311 15802
rect 2335 15750 2349 15802
rect 2349 15750 2361 15802
rect 2361 15750 2391 15802
rect 2415 15750 2425 15802
rect 2425 15750 2471 15802
rect 2175 15748 2231 15750
rect 2255 15748 2311 15750
rect 2335 15748 2391 15750
rect 2415 15748 2471 15750
rect 4613 15802 4669 15804
rect 4693 15802 4749 15804
rect 4773 15802 4829 15804
rect 4853 15802 4909 15804
rect 4613 15750 4659 15802
rect 4659 15750 4669 15802
rect 4693 15750 4723 15802
rect 4723 15750 4735 15802
rect 4735 15750 4749 15802
rect 4773 15750 4787 15802
rect 4787 15750 4799 15802
rect 4799 15750 4829 15802
rect 4853 15750 4863 15802
rect 4863 15750 4909 15802
rect 4613 15748 4669 15750
rect 4693 15748 4749 15750
rect 4773 15748 4829 15750
rect 4853 15748 4909 15750
rect 7051 15802 7107 15804
rect 7131 15802 7187 15804
rect 7211 15802 7267 15804
rect 7291 15802 7347 15804
rect 7051 15750 7097 15802
rect 7097 15750 7107 15802
rect 7131 15750 7161 15802
rect 7161 15750 7173 15802
rect 7173 15750 7187 15802
rect 7211 15750 7225 15802
rect 7225 15750 7237 15802
rect 7237 15750 7267 15802
rect 7291 15750 7301 15802
rect 7301 15750 7347 15802
rect 7051 15748 7107 15750
rect 7131 15748 7187 15750
rect 7211 15748 7267 15750
rect 7291 15748 7347 15750
rect 9489 15802 9545 15804
rect 9569 15802 9625 15804
rect 9649 15802 9705 15804
rect 9729 15802 9785 15804
rect 9489 15750 9535 15802
rect 9535 15750 9545 15802
rect 9569 15750 9599 15802
rect 9599 15750 9611 15802
rect 9611 15750 9625 15802
rect 9649 15750 9663 15802
rect 9663 15750 9675 15802
rect 9675 15750 9705 15802
rect 9729 15750 9739 15802
rect 9739 15750 9785 15802
rect 9489 15748 9545 15750
rect 9569 15748 9625 15750
rect 9649 15748 9705 15750
rect 9729 15748 9785 15750
rect 3394 15258 3450 15260
rect 3474 15258 3530 15260
rect 3554 15258 3610 15260
rect 3634 15258 3690 15260
rect 3394 15206 3440 15258
rect 3440 15206 3450 15258
rect 3474 15206 3504 15258
rect 3504 15206 3516 15258
rect 3516 15206 3530 15258
rect 3554 15206 3568 15258
rect 3568 15206 3580 15258
rect 3580 15206 3610 15258
rect 3634 15206 3644 15258
rect 3644 15206 3690 15258
rect 3394 15204 3450 15206
rect 3474 15204 3530 15206
rect 3554 15204 3610 15206
rect 3634 15204 3690 15206
rect 2175 14714 2231 14716
rect 2255 14714 2311 14716
rect 2335 14714 2391 14716
rect 2415 14714 2471 14716
rect 2175 14662 2221 14714
rect 2221 14662 2231 14714
rect 2255 14662 2285 14714
rect 2285 14662 2297 14714
rect 2297 14662 2311 14714
rect 2335 14662 2349 14714
rect 2349 14662 2361 14714
rect 2361 14662 2391 14714
rect 2415 14662 2425 14714
rect 2425 14662 2471 14714
rect 2175 14660 2231 14662
rect 2255 14660 2311 14662
rect 2335 14660 2391 14662
rect 2415 14660 2471 14662
rect 4613 14714 4669 14716
rect 4693 14714 4749 14716
rect 4773 14714 4829 14716
rect 4853 14714 4909 14716
rect 4613 14662 4659 14714
rect 4659 14662 4669 14714
rect 4693 14662 4723 14714
rect 4723 14662 4735 14714
rect 4735 14662 4749 14714
rect 4773 14662 4787 14714
rect 4787 14662 4799 14714
rect 4799 14662 4829 14714
rect 4853 14662 4863 14714
rect 4863 14662 4909 14714
rect 4613 14660 4669 14662
rect 4693 14660 4749 14662
rect 4773 14660 4829 14662
rect 4853 14660 4909 14662
rect 938 14340 994 14376
rect 938 14320 940 14340
rect 940 14320 992 14340
rect 992 14320 994 14340
rect 2175 13626 2231 13628
rect 2255 13626 2311 13628
rect 2335 13626 2391 13628
rect 2415 13626 2471 13628
rect 2175 13574 2221 13626
rect 2221 13574 2231 13626
rect 2255 13574 2285 13626
rect 2285 13574 2297 13626
rect 2297 13574 2311 13626
rect 2335 13574 2349 13626
rect 2349 13574 2361 13626
rect 2361 13574 2391 13626
rect 2415 13574 2425 13626
rect 2425 13574 2471 13626
rect 2175 13572 2231 13574
rect 2255 13572 2311 13574
rect 2335 13572 2391 13574
rect 2415 13572 2471 13574
rect 2175 12538 2231 12540
rect 2255 12538 2311 12540
rect 2335 12538 2391 12540
rect 2415 12538 2471 12540
rect 2175 12486 2221 12538
rect 2221 12486 2231 12538
rect 2255 12486 2285 12538
rect 2285 12486 2297 12538
rect 2297 12486 2311 12538
rect 2335 12486 2349 12538
rect 2349 12486 2361 12538
rect 2361 12486 2391 12538
rect 2415 12486 2425 12538
rect 2425 12486 2471 12538
rect 2175 12484 2231 12486
rect 2255 12484 2311 12486
rect 2335 12484 2391 12486
rect 2415 12484 2471 12486
rect 938 12164 994 12200
rect 938 12144 940 12164
rect 940 12144 992 12164
rect 992 12144 994 12164
rect 3394 14170 3450 14172
rect 3474 14170 3530 14172
rect 3554 14170 3610 14172
rect 3634 14170 3690 14172
rect 3394 14118 3440 14170
rect 3440 14118 3450 14170
rect 3474 14118 3504 14170
rect 3504 14118 3516 14170
rect 3516 14118 3530 14170
rect 3554 14118 3568 14170
rect 3568 14118 3580 14170
rect 3580 14118 3610 14170
rect 3634 14118 3644 14170
rect 3644 14118 3690 14170
rect 3394 14116 3450 14118
rect 3474 14116 3530 14118
rect 3554 14116 3610 14118
rect 3634 14116 3690 14118
rect 4613 13626 4669 13628
rect 4693 13626 4749 13628
rect 4773 13626 4829 13628
rect 4853 13626 4909 13628
rect 4613 13574 4659 13626
rect 4659 13574 4669 13626
rect 4693 13574 4723 13626
rect 4723 13574 4735 13626
rect 4735 13574 4749 13626
rect 4773 13574 4787 13626
rect 4787 13574 4799 13626
rect 4799 13574 4829 13626
rect 4853 13574 4863 13626
rect 4863 13574 4909 13626
rect 4613 13572 4669 13574
rect 4693 13572 4749 13574
rect 4773 13572 4829 13574
rect 4853 13572 4909 13574
rect 3394 13082 3450 13084
rect 3474 13082 3530 13084
rect 3554 13082 3610 13084
rect 3634 13082 3690 13084
rect 3394 13030 3440 13082
rect 3440 13030 3450 13082
rect 3474 13030 3504 13082
rect 3504 13030 3516 13082
rect 3516 13030 3530 13082
rect 3554 13030 3568 13082
rect 3568 13030 3580 13082
rect 3580 13030 3610 13082
rect 3634 13030 3644 13082
rect 3644 13030 3690 13082
rect 3394 13028 3450 13030
rect 3474 13028 3530 13030
rect 3554 13028 3610 13030
rect 3634 13028 3690 13030
rect 4613 12538 4669 12540
rect 4693 12538 4749 12540
rect 4773 12538 4829 12540
rect 4853 12538 4909 12540
rect 4613 12486 4659 12538
rect 4659 12486 4669 12538
rect 4693 12486 4723 12538
rect 4723 12486 4735 12538
rect 4735 12486 4749 12538
rect 4773 12486 4787 12538
rect 4787 12486 4799 12538
rect 4799 12486 4829 12538
rect 4853 12486 4863 12538
rect 4863 12486 4909 12538
rect 4613 12484 4669 12486
rect 4693 12484 4749 12486
rect 4773 12484 4829 12486
rect 4853 12484 4909 12486
rect 3394 11994 3450 11996
rect 3474 11994 3530 11996
rect 3554 11994 3610 11996
rect 3634 11994 3690 11996
rect 3394 11942 3440 11994
rect 3440 11942 3450 11994
rect 3474 11942 3504 11994
rect 3504 11942 3516 11994
rect 3516 11942 3530 11994
rect 3554 11942 3568 11994
rect 3568 11942 3580 11994
rect 3580 11942 3610 11994
rect 3634 11942 3644 11994
rect 3644 11942 3690 11994
rect 3394 11940 3450 11942
rect 3474 11940 3530 11942
rect 3554 11940 3610 11942
rect 3634 11940 3690 11942
rect 5832 15258 5888 15260
rect 5912 15258 5968 15260
rect 5992 15258 6048 15260
rect 6072 15258 6128 15260
rect 5832 15206 5878 15258
rect 5878 15206 5888 15258
rect 5912 15206 5942 15258
rect 5942 15206 5954 15258
rect 5954 15206 5968 15258
rect 5992 15206 6006 15258
rect 6006 15206 6018 15258
rect 6018 15206 6048 15258
rect 6072 15206 6082 15258
rect 6082 15206 6128 15258
rect 5832 15204 5888 15206
rect 5912 15204 5968 15206
rect 5992 15204 6048 15206
rect 6072 15204 6128 15206
rect 8270 15258 8326 15260
rect 8350 15258 8406 15260
rect 8430 15258 8486 15260
rect 8510 15258 8566 15260
rect 8270 15206 8316 15258
rect 8316 15206 8326 15258
rect 8350 15206 8380 15258
rect 8380 15206 8392 15258
rect 8392 15206 8406 15258
rect 8430 15206 8444 15258
rect 8444 15206 8456 15258
rect 8456 15206 8486 15258
rect 8510 15206 8520 15258
rect 8520 15206 8566 15258
rect 8270 15204 8326 15206
rect 8350 15204 8406 15206
rect 8430 15204 8486 15206
rect 8510 15204 8566 15206
rect 10708 15258 10764 15260
rect 10788 15258 10844 15260
rect 10868 15258 10924 15260
rect 10948 15258 11004 15260
rect 10708 15206 10754 15258
rect 10754 15206 10764 15258
rect 10788 15206 10818 15258
rect 10818 15206 10830 15258
rect 10830 15206 10844 15258
rect 10868 15206 10882 15258
rect 10882 15206 10894 15258
rect 10894 15206 10924 15258
rect 10948 15206 10958 15258
rect 10958 15206 11004 15258
rect 10708 15204 10764 15206
rect 10788 15204 10844 15206
rect 10868 15204 10924 15206
rect 10948 15204 11004 15206
rect 7051 14714 7107 14716
rect 7131 14714 7187 14716
rect 7211 14714 7267 14716
rect 7291 14714 7347 14716
rect 7051 14662 7097 14714
rect 7097 14662 7107 14714
rect 7131 14662 7161 14714
rect 7161 14662 7173 14714
rect 7173 14662 7187 14714
rect 7211 14662 7225 14714
rect 7225 14662 7237 14714
rect 7237 14662 7267 14714
rect 7291 14662 7301 14714
rect 7301 14662 7347 14714
rect 7051 14660 7107 14662
rect 7131 14660 7187 14662
rect 7211 14660 7267 14662
rect 7291 14660 7347 14662
rect 9489 14714 9545 14716
rect 9569 14714 9625 14716
rect 9649 14714 9705 14716
rect 9729 14714 9785 14716
rect 9489 14662 9535 14714
rect 9535 14662 9545 14714
rect 9569 14662 9599 14714
rect 9599 14662 9611 14714
rect 9611 14662 9625 14714
rect 9649 14662 9663 14714
rect 9663 14662 9675 14714
rect 9675 14662 9705 14714
rect 9729 14662 9739 14714
rect 9739 14662 9785 14714
rect 9489 14660 9545 14662
rect 9569 14660 9625 14662
rect 9649 14660 9705 14662
rect 9729 14660 9785 14662
rect 5832 14170 5888 14172
rect 5912 14170 5968 14172
rect 5992 14170 6048 14172
rect 6072 14170 6128 14172
rect 5832 14118 5878 14170
rect 5878 14118 5888 14170
rect 5912 14118 5942 14170
rect 5942 14118 5954 14170
rect 5954 14118 5968 14170
rect 5992 14118 6006 14170
rect 6006 14118 6018 14170
rect 6018 14118 6048 14170
rect 6072 14118 6082 14170
rect 6082 14118 6128 14170
rect 5832 14116 5888 14118
rect 5912 14116 5968 14118
rect 5992 14116 6048 14118
rect 6072 14116 6128 14118
rect 8270 14170 8326 14172
rect 8350 14170 8406 14172
rect 8430 14170 8486 14172
rect 8510 14170 8566 14172
rect 8270 14118 8316 14170
rect 8316 14118 8326 14170
rect 8350 14118 8380 14170
rect 8380 14118 8392 14170
rect 8392 14118 8406 14170
rect 8430 14118 8444 14170
rect 8444 14118 8456 14170
rect 8456 14118 8486 14170
rect 8510 14118 8520 14170
rect 8520 14118 8566 14170
rect 8270 14116 8326 14118
rect 8350 14116 8406 14118
rect 8430 14116 8486 14118
rect 8510 14116 8566 14118
rect 10708 14170 10764 14172
rect 10788 14170 10844 14172
rect 10868 14170 10924 14172
rect 10948 14170 11004 14172
rect 10708 14118 10754 14170
rect 10754 14118 10764 14170
rect 10788 14118 10818 14170
rect 10818 14118 10830 14170
rect 10830 14118 10844 14170
rect 10868 14118 10882 14170
rect 10882 14118 10894 14170
rect 10894 14118 10924 14170
rect 10948 14118 10958 14170
rect 10958 14118 11004 14170
rect 10708 14116 10764 14118
rect 10788 14116 10844 14118
rect 10868 14116 10924 14118
rect 10948 14116 11004 14118
rect 7051 13626 7107 13628
rect 7131 13626 7187 13628
rect 7211 13626 7267 13628
rect 7291 13626 7347 13628
rect 7051 13574 7097 13626
rect 7097 13574 7107 13626
rect 7131 13574 7161 13626
rect 7161 13574 7173 13626
rect 7173 13574 7187 13626
rect 7211 13574 7225 13626
rect 7225 13574 7237 13626
rect 7237 13574 7267 13626
rect 7291 13574 7301 13626
rect 7301 13574 7347 13626
rect 7051 13572 7107 13574
rect 7131 13572 7187 13574
rect 7211 13572 7267 13574
rect 7291 13572 7347 13574
rect 9489 13626 9545 13628
rect 9569 13626 9625 13628
rect 9649 13626 9705 13628
rect 9729 13626 9785 13628
rect 9489 13574 9535 13626
rect 9535 13574 9545 13626
rect 9569 13574 9599 13626
rect 9599 13574 9611 13626
rect 9611 13574 9625 13626
rect 9649 13574 9663 13626
rect 9663 13574 9675 13626
rect 9675 13574 9705 13626
rect 9729 13574 9739 13626
rect 9739 13574 9785 13626
rect 9489 13572 9545 13574
rect 9569 13572 9625 13574
rect 9649 13572 9705 13574
rect 9729 13572 9785 13574
rect 5832 13082 5888 13084
rect 5912 13082 5968 13084
rect 5992 13082 6048 13084
rect 6072 13082 6128 13084
rect 5832 13030 5878 13082
rect 5878 13030 5888 13082
rect 5912 13030 5942 13082
rect 5942 13030 5954 13082
rect 5954 13030 5968 13082
rect 5992 13030 6006 13082
rect 6006 13030 6018 13082
rect 6018 13030 6048 13082
rect 6072 13030 6082 13082
rect 6082 13030 6128 13082
rect 5832 13028 5888 13030
rect 5912 13028 5968 13030
rect 5992 13028 6048 13030
rect 6072 13028 6128 13030
rect 8270 13082 8326 13084
rect 8350 13082 8406 13084
rect 8430 13082 8486 13084
rect 8510 13082 8566 13084
rect 8270 13030 8316 13082
rect 8316 13030 8326 13082
rect 8350 13030 8380 13082
rect 8380 13030 8392 13082
rect 8392 13030 8406 13082
rect 8430 13030 8444 13082
rect 8444 13030 8456 13082
rect 8456 13030 8486 13082
rect 8510 13030 8520 13082
rect 8520 13030 8566 13082
rect 8270 13028 8326 13030
rect 8350 13028 8406 13030
rect 8430 13028 8486 13030
rect 8510 13028 8566 13030
rect 10708 13082 10764 13084
rect 10788 13082 10844 13084
rect 10868 13082 10924 13084
rect 10948 13082 11004 13084
rect 10708 13030 10754 13082
rect 10754 13030 10764 13082
rect 10788 13030 10818 13082
rect 10818 13030 10830 13082
rect 10830 13030 10844 13082
rect 10868 13030 10882 13082
rect 10882 13030 10894 13082
rect 10894 13030 10924 13082
rect 10948 13030 10958 13082
rect 10958 13030 11004 13082
rect 10708 13028 10764 13030
rect 10788 13028 10844 13030
rect 10868 13028 10924 13030
rect 10948 13028 11004 13030
rect 7051 12538 7107 12540
rect 7131 12538 7187 12540
rect 7211 12538 7267 12540
rect 7291 12538 7347 12540
rect 7051 12486 7097 12538
rect 7097 12486 7107 12538
rect 7131 12486 7161 12538
rect 7161 12486 7173 12538
rect 7173 12486 7187 12538
rect 7211 12486 7225 12538
rect 7225 12486 7237 12538
rect 7237 12486 7267 12538
rect 7291 12486 7301 12538
rect 7301 12486 7347 12538
rect 7051 12484 7107 12486
rect 7131 12484 7187 12486
rect 7211 12484 7267 12486
rect 7291 12484 7347 12486
rect 9489 12538 9545 12540
rect 9569 12538 9625 12540
rect 9649 12538 9705 12540
rect 9729 12538 9785 12540
rect 9489 12486 9535 12538
rect 9535 12486 9545 12538
rect 9569 12486 9599 12538
rect 9599 12486 9611 12538
rect 9611 12486 9625 12538
rect 9649 12486 9663 12538
rect 9663 12486 9675 12538
rect 9675 12486 9705 12538
rect 9729 12486 9739 12538
rect 9739 12486 9785 12538
rect 9489 12484 9545 12486
rect 9569 12484 9625 12486
rect 9649 12484 9705 12486
rect 9729 12484 9785 12486
rect 5832 11994 5888 11996
rect 5912 11994 5968 11996
rect 5992 11994 6048 11996
rect 6072 11994 6128 11996
rect 5832 11942 5878 11994
rect 5878 11942 5888 11994
rect 5912 11942 5942 11994
rect 5942 11942 5954 11994
rect 5954 11942 5968 11994
rect 5992 11942 6006 11994
rect 6006 11942 6018 11994
rect 6018 11942 6048 11994
rect 6072 11942 6082 11994
rect 6082 11942 6128 11994
rect 5832 11940 5888 11942
rect 5912 11940 5968 11942
rect 5992 11940 6048 11942
rect 6072 11940 6128 11942
rect 8270 11994 8326 11996
rect 8350 11994 8406 11996
rect 8430 11994 8486 11996
rect 8510 11994 8566 11996
rect 8270 11942 8316 11994
rect 8316 11942 8326 11994
rect 8350 11942 8380 11994
rect 8380 11942 8392 11994
rect 8392 11942 8406 11994
rect 8430 11942 8444 11994
rect 8444 11942 8456 11994
rect 8456 11942 8486 11994
rect 8510 11942 8520 11994
rect 8520 11942 8566 11994
rect 8270 11940 8326 11942
rect 8350 11940 8406 11942
rect 8430 11940 8486 11942
rect 8510 11940 8566 11942
rect 10708 11994 10764 11996
rect 10788 11994 10844 11996
rect 10868 11994 10924 11996
rect 10948 11994 11004 11996
rect 10708 11942 10754 11994
rect 10754 11942 10764 11994
rect 10788 11942 10818 11994
rect 10818 11942 10830 11994
rect 10830 11942 10844 11994
rect 10868 11942 10882 11994
rect 10882 11942 10894 11994
rect 10894 11942 10924 11994
rect 10948 11942 10958 11994
rect 10958 11942 11004 11994
rect 10708 11940 10764 11942
rect 10788 11940 10844 11942
rect 10868 11940 10924 11942
rect 10948 11940 11004 11942
rect 2175 11450 2231 11452
rect 2255 11450 2311 11452
rect 2335 11450 2391 11452
rect 2415 11450 2471 11452
rect 2175 11398 2221 11450
rect 2221 11398 2231 11450
rect 2255 11398 2285 11450
rect 2285 11398 2297 11450
rect 2297 11398 2311 11450
rect 2335 11398 2349 11450
rect 2349 11398 2361 11450
rect 2361 11398 2391 11450
rect 2415 11398 2425 11450
rect 2425 11398 2471 11450
rect 2175 11396 2231 11398
rect 2255 11396 2311 11398
rect 2335 11396 2391 11398
rect 2415 11396 2471 11398
rect 938 10004 940 10024
rect 940 10004 992 10024
rect 992 10004 994 10024
rect 938 9968 994 10004
rect 2175 10362 2231 10364
rect 2255 10362 2311 10364
rect 2335 10362 2391 10364
rect 2415 10362 2471 10364
rect 2175 10310 2221 10362
rect 2221 10310 2231 10362
rect 2255 10310 2285 10362
rect 2285 10310 2297 10362
rect 2297 10310 2311 10362
rect 2335 10310 2349 10362
rect 2349 10310 2361 10362
rect 2361 10310 2391 10362
rect 2415 10310 2425 10362
rect 2425 10310 2471 10362
rect 2175 10308 2231 10310
rect 2255 10308 2311 10310
rect 2335 10308 2391 10310
rect 2415 10308 2471 10310
rect 938 7792 994 7848
rect 938 5652 940 5672
rect 940 5652 992 5672
rect 992 5652 994 5672
rect 938 5616 994 5652
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 938 3440 994 3496
rect 4613 11450 4669 11452
rect 4693 11450 4749 11452
rect 4773 11450 4829 11452
rect 4853 11450 4909 11452
rect 4613 11398 4659 11450
rect 4659 11398 4669 11450
rect 4693 11398 4723 11450
rect 4723 11398 4735 11450
rect 4735 11398 4749 11450
rect 4773 11398 4787 11450
rect 4787 11398 4799 11450
rect 4799 11398 4829 11450
rect 4853 11398 4863 11450
rect 4863 11398 4909 11450
rect 4613 11396 4669 11398
rect 4693 11396 4749 11398
rect 4773 11396 4829 11398
rect 4853 11396 4909 11398
rect 3394 10906 3450 10908
rect 3474 10906 3530 10908
rect 3554 10906 3610 10908
rect 3634 10906 3690 10908
rect 3394 10854 3440 10906
rect 3440 10854 3450 10906
rect 3474 10854 3504 10906
rect 3504 10854 3516 10906
rect 3516 10854 3530 10906
rect 3554 10854 3568 10906
rect 3568 10854 3580 10906
rect 3580 10854 3610 10906
rect 3634 10854 3644 10906
rect 3644 10854 3690 10906
rect 3394 10852 3450 10854
rect 3474 10852 3530 10854
rect 3554 10852 3610 10854
rect 3634 10852 3690 10854
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 4613 10362 4669 10364
rect 4693 10362 4749 10364
rect 4773 10362 4829 10364
rect 4853 10362 4909 10364
rect 4613 10310 4659 10362
rect 4659 10310 4669 10362
rect 4693 10310 4723 10362
rect 4723 10310 4735 10362
rect 4735 10310 4749 10362
rect 4773 10310 4787 10362
rect 4787 10310 4799 10362
rect 4799 10310 4829 10362
rect 4853 10310 4863 10362
rect 4863 10310 4909 10362
rect 4613 10308 4669 10310
rect 4693 10308 4749 10310
rect 4773 10308 4829 10310
rect 4853 10308 4909 10310
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 938 1264 994 1320
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 5832 10906 5888 10908
rect 5912 10906 5968 10908
rect 5992 10906 6048 10908
rect 6072 10906 6128 10908
rect 5832 10854 5878 10906
rect 5878 10854 5888 10906
rect 5912 10854 5942 10906
rect 5942 10854 5954 10906
rect 5954 10854 5968 10906
rect 5992 10854 6006 10906
rect 6006 10854 6018 10906
rect 6018 10854 6048 10906
rect 6072 10854 6082 10906
rect 6082 10854 6128 10906
rect 5832 10852 5888 10854
rect 5912 10852 5968 10854
rect 5992 10852 6048 10854
rect 6072 10852 6128 10854
rect 7051 11450 7107 11452
rect 7131 11450 7187 11452
rect 7211 11450 7267 11452
rect 7291 11450 7347 11452
rect 7051 11398 7097 11450
rect 7097 11398 7107 11450
rect 7131 11398 7161 11450
rect 7161 11398 7173 11450
rect 7173 11398 7187 11450
rect 7211 11398 7225 11450
rect 7225 11398 7237 11450
rect 7237 11398 7267 11450
rect 7291 11398 7301 11450
rect 7301 11398 7347 11450
rect 7051 11396 7107 11398
rect 7131 11396 7187 11398
rect 7211 11396 7267 11398
rect 7291 11396 7347 11398
rect 9489 11450 9545 11452
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9489 11398 9535 11450
rect 9535 11398 9545 11450
rect 9569 11398 9599 11450
rect 9599 11398 9611 11450
rect 9611 11398 9625 11450
rect 9649 11398 9663 11450
rect 9663 11398 9675 11450
rect 9675 11398 9705 11450
rect 9729 11398 9739 11450
rect 9739 11398 9785 11450
rect 9489 11396 9545 11398
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 7051 10362 7107 10364
rect 7131 10362 7187 10364
rect 7211 10362 7267 10364
rect 7291 10362 7347 10364
rect 7051 10310 7097 10362
rect 7097 10310 7107 10362
rect 7131 10310 7161 10362
rect 7161 10310 7173 10362
rect 7173 10310 7187 10362
rect 7211 10310 7225 10362
rect 7225 10310 7237 10362
rect 7237 10310 7267 10362
rect 7291 10310 7301 10362
rect 7301 10310 7347 10362
rect 7051 10308 7107 10310
rect 7131 10308 7187 10310
rect 7211 10308 7267 10310
rect 7291 10308 7347 10310
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 8270 10906 8326 10908
rect 8350 10906 8406 10908
rect 8430 10906 8486 10908
rect 8510 10906 8566 10908
rect 8270 10854 8316 10906
rect 8316 10854 8326 10906
rect 8350 10854 8380 10906
rect 8380 10854 8392 10906
rect 8392 10854 8406 10906
rect 8430 10854 8444 10906
rect 8444 10854 8456 10906
rect 8456 10854 8486 10906
rect 8510 10854 8520 10906
rect 8520 10854 8566 10906
rect 8270 10852 8326 10854
rect 8350 10852 8406 10854
rect 8430 10852 8486 10854
rect 8510 10852 8566 10854
rect 10708 10906 10764 10908
rect 10788 10906 10844 10908
rect 10868 10906 10924 10908
rect 10948 10906 11004 10908
rect 10708 10854 10754 10906
rect 10754 10854 10764 10906
rect 10788 10854 10818 10906
rect 10818 10854 10830 10906
rect 10830 10854 10844 10906
rect 10868 10854 10882 10906
rect 10882 10854 10894 10906
rect 10894 10854 10924 10906
rect 10948 10854 10958 10906
rect 10958 10854 11004 10906
rect 10708 10852 10764 10854
rect 10788 10852 10844 10854
rect 10868 10852 10924 10854
rect 10948 10852 11004 10854
rect 9489 10362 9545 10364
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9489 10310 9535 10362
rect 9535 10310 9545 10362
rect 9569 10310 9599 10362
rect 9599 10310 9611 10362
rect 9611 10310 9625 10362
rect 9649 10310 9663 10362
rect 9663 10310 9675 10362
rect 9675 10310 9705 10362
rect 9729 10310 9739 10362
rect 9739 10310 9785 10362
rect 9489 10308 9545 10310
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
<< metal3 >>
rect 0 16554 800 16584
rect 933 16554 999 16557
rect 0 16552 999 16554
rect 0 16496 938 16552
rect 994 16496 999 16552
rect 0 16494 999 16496
rect 0 16464 800 16494
rect 933 16491 999 16494
rect 2165 15808 2481 15809
rect 2165 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2481 15808
rect 2165 15743 2481 15744
rect 4603 15808 4919 15809
rect 4603 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4919 15808
rect 4603 15743 4919 15744
rect 7041 15808 7357 15809
rect 7041 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7357 15808
rect 7041 15743 7357 15744
rect 9479 15808 9795 15809
rect 9479 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9795 15808
rect 9479 15743 9795 15744
rect 3384 15264 3700 15265
rect 3384 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3700 15264
rect 3384 15199 3700 15200
rect 5822 15264 6138 15265
rect 5822 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6138 15264
rect 5822 15199 6138 15200
rect 8260 15264 8576 15265
rect 8260 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8576 15264
rect 8260 15199 8576 15200
rect 10698 15264 11014 15265
rect 10698 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11014 15264
rect 10698 15199 11014 15200
rect 2165 14720 2481 14721
rect 2165 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2481 14720
rect 2165 14655 2481 14656
rect 4603 14720 4919 14721
rect 4603 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4919 14720
rect 4603 14655 4919 14656
rect 7041 14720 7357 14721
rect 7041 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7357 14720
rect 7041 14655 7357 14656
rect 9479 14720 9795 14721
rect 9479 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9795 14720
rect 9479 14655 9795 14656
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 3384 14176 3700 14177
rect 3384 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3700 14176
rect 3384 14111 3700 14112
rect 5822 14176 6138 14177
rect 5822 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6138 14176
rect 5822 14111 6138 14112
rect 8260 14176 8576 14177
rect 8260 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8576 14176
rect 8260 14111 8576 14112
rect 10698 14176 11014 14177
rect 10698 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11014 14176
rect 10698 14111 11014 14112
rect 2165 13632 2481 13633
rect 2165 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2481 13632
rect 2165 13567 2481 13568
rect 4603 13632 4919 13633
rect 4603 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4919 13632
rect 4603 13567 4919 13568
rect 7041 13632 7357 13633
rect 7041 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7357 13632
rect 7041 13567 7357 13568
rect 9479 13632 9795 13633
rect 9479 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9795 13632
rect 9479 13567 9795 13568
rect 3384 13088 3700 13089
rect 3384 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3700 13088
rect 3384 13023 3700 13024
rect 5822 13088 6138 13089
rect 5822 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6138 13088
rect 5822 13023 6138 13024
rect 8260 13088 8576 13089
rect 8260 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8576 13088
rect 8260 13023 8576 13024
rect 10698 13088 11014 13089
rect 10698 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11014 13088
rect 10698 13023 11014 13024
rect 2165 12544 2481 12545
rect 2165 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2481 12544
rect 2165 12479 2481 12480
rect 4603 12544 4919 12545
rect 4603 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4919 12544
rect 4603 12479 4919 12480
rect 7041 12544 7357 12545
rect 7041 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7357 12544
rect 7041 12479 7357 12480
rect 9479 12544 9795 12545
rect 9479 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9795 12544
rect 9479 12479 9795 12480
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 3384 12000 3700 12001
rect 3384 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3700 12000
rect 3384 11935 3700 11936
rect 5822 12000 6138 12001
rect 5822 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6138 12000
rect 5822 11935 6138 11936
rect 8260 12000 8576 12001
rect 8260 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8576 12000
rect 8260 11935 8576 11936
rect 10698 12000 11014 12001
rect 10698 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11014 12000
rect 10698 11935 11014 11936
rect 2165 11456 2481 11457
rect 2165 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2481 11456
rect 2165 11391 2481 11392
rect 4603 11456 4919 11457
rect 4603 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4919 11456
rect 4603 11391 4919 11392
rect 7041 11456 7357 11457
rect 7041 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7357 11456
rect 7041 11391 7357 11392
rect 9479 11456 9795 11457
rect 9479 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9795 11456
rect 9479 11391 9795 11392
rect 3384 10912 3700 10913
rect 3384 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3700 10912
rect 3384 10847 3700 10848
rect 5822 10912 6138 10913
rect 5822 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6138 10912
rect 5822 10847 6138 10848
rect 8260 10912 8576 10913
rect 8260 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8576 10912
rect 8260 10847 8576 10848
rect 10698 10912 11014 10913
rect 10698 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11014 10912
rect 10698 10847 11014 10848
rect 2165 10368 2481 10369
rect 2165 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2481 10368
rect 2165 10303 2481 10304
rect 4603 10368 4919 10369
rect 4603 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4919 10368
rect 4603 10303 4919 10304
rect 7041 10368 7357 10369
rect 7041 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7357 10368
rect 7041 10303 7357 10304
rect 9479 10368 9795 10369
rect 9479 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9795 10368
rect 9479 10303 9795 10304
rect 0 10026 800 10056
rect 933 10026 999 10029
rect 0 10024 999 10026
rect 0 9968 938 10024
rect 994 9968 999 10024
rect 0 9966 999 9968
rect 0 9936 800 9966
rect 933 9963 999 9966
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7850 800 7880
rect 933 7850 999 7853
rect 0 7848 999 7850
rect 0 7792 938 7848
rect 994 7792 999 7848
rect 0 7790 999 7792
rect 0 7760 800 7790
rect 933 7787 999 7790
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 0 5674 800 5704
rect 933 5674 999 5677
rect 0 5672 999 5674
rect 0 5616 938 5672
rect 994 5616 999 5672
rect 0 5614 999 5616
rect 0 5584 800 5614
rect 933 5611 999 5614
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 0 1322 800 1352
rect 933 1322 999 1325
rect 0 1320 999 1322
rect 0 1264 938 1320
rect 994 1264 999 1320
rect 0 1262 999 1264
rect 0 1232 800 1262
rect 933 1259 999 1262
<< via3 >>
rect 2171 15804 2235 15808
rect 2171 15748 2175 15804
rect 2175 15748 2231 15804
rect 2231 15748 2235 15804
rect 2171 15744 2235 15748
rect 2251 15804 2315 15808
rect 2251 15748 2255 15804
rect 2255 15748 2311 15804
rect 2311 15748 2315 15804
rect 2251 15744 2315 15748
rect 2331 15804 2395 15808
rect 2331 15748 2335 15804
rect 2335 15748 2391 15804
rect 2391 15748 2395 15804
rect 2331 15744 2395 15748
rect 2411 15804 2475 15808
rect 2411 15748 2415 15804
rect 2415 15748 2471 15804
rect 2471 15748 2475 15804
rect 2411 15744 2475 15748
rect 4609 15804 4673 15808
rect 4609 15748 4613 15804
rect 4613 15748 4669 15804
rect 4669 15748 4673 15804
rect 4609 15744 4673 15748
rect 4689 15804 4753 15808
rect 4689 15748 4693 15804
rect 4693 15748 4749 15804
rect 4749 15748 4753 15804
rect 4689 15744 4753 15748
rect 4769 15804 4833 15808
rect 4769 15748 4773 15804
rect 4773 15748 4829 15804
rect 4829 15748 4833 15804
rect 4769 15744 4833 15748
rect 4849 15804 4913 15808
rect 4849 15748 4853 15804
rect 4853 15748 4909 15804
rect 4909 15748 4913 15804
rect 4849 15744 4913 15748
rect 7047 15804 7111 15808
rect 7047 15748 7051 15804
rect 7051 15748 7107 15804
rect 7107 15748 7111 15804
rect 7047 15744 7111 15748
rect 7127 15804 7191 15808
rect 7127 15748 7131 15804
rect 7131 15748 7187 15804
rect 7187 15748 7191 15804
rect 7127 15744 7191 15748
rect 7207 15804 7271 15808
rect 7207 15748 7211 15804
rect 7211 15748 7267 15804
rect 7267 15748 7271 15804
rect 7207 15744 7271 15748
rect 7287 15804 7351 15808
rect 7287 15748 7291 15804
rect 7291 15748 7347 15804
rect 7347 15748 7351 15804
rect 7287 15744 7351 15748
rect 9485 15804 9549 15808
rect 9485 15748 9489 15804
rect 9489 15748 9545 15804
rect 9545 15748 9549 15804
rect 9485 15744 9549 15748
rect 9565 15804 9629 15808
rect 9565 15748 9569 15804
rect 9569 15748 9625 15804
rect 9625 15748 9629 15804
rect 9565 15744 9629 15748
rect 9645 15804 9709 15808
rect 9645 15748 9649 15804
rect 9649 15748 9705 15804
rect 9705 15748 9709 15804
rect 9645 15744 9709 15748
rect 9725 15804 9789 15808
rect 9725 15748 9729 15804
rect 9729 15748 9785 15804
rect 9785 15748 9789 15804
rect 9725 15744 9789 15748
rect 3390 15260 3454 15264
rect 3390 15204 3394 15260
rect 3394 15204 3450 15260
rect 3450 15204 3454 15260
rect 3390 15200 3454 15204
rect 3470 15260 3534 15264
rect 3470 15204 3474 15260
rect 3474 15204 3530 15260
rect 3530 15204 3534 15260
rect 3470 15200 3534 15204
rect 3550 15260 3614 15264
rect 3550 15204 3554 15260
rect 3554 15204 3610 15260
rect 3610 15204 3614 15260
rect 3550 15200 3614 15204
rect 3630 15260 3694 15264
rect 3630 15204 3634 15260
rect 3634 15204 3690 15260
rect 3690 15204 3694 15260
rect 3630 15200 3694 15204
rect 5828 15260 5892 15264
rect 5828 15204 5832 15260
rect 5832 15204 5888 15260
rect 5888 15204 5892 15260
rect 5828 15200 5892 15204
rect 5908 15260 5972 15264
rect 5908 15204 5912 15260
rect 5912 15204 5968 15260
rect 5968 15204 5972 15260
rect 5908 15200 5972 15204
rect 5988 15260 6052 15264
rect 5988 15204 5992 15260
rect 5992 15204 6048 15260
rect 6048 15204 6052 15260
rect 5988 15200 6052 15204
rect 6068 15260 6132 15264
rect 6068 15204 6072 15260
rect 6072 15204 6128 15260
rect 6128 15204 6132 15260
rect 6068 15200 6132 15204
rect 8266 15260 8330 15264
rect 8266 15204 8270 15260
rect 8270 15204 8326 15260
rect 8326 15204 8330 15260
rect 8266 15200 8330 15204
rect 8346 15260 8410 15264
rect 8346 15204 8350 15260
rect 8350 15204 8406 15260
rect 8406 15204 8410 15260
rect 8346 15200 8410 15204
rect 8426 15260 8490 15264
rect 8426 15204 8430 15260
rect 8430 15204 8486 15260
rect 8486 15204 8490 15260
rect 8426 15200 8490 15204
rect 8506 15260 8570 15264
rect 8506 15204 8510 15260
rect 8510 15204 8566 15260
rect 8566 15204 8570 15260
rect 8506 15200 8570 15204
rect 10704 15260 10768 15264
rect 10704 15204 10708 15260
rect 10708 15204 10764 15260
rect 10764 15204 10768 15260
rect 10704 15200 10768 15204
rect 10784 15260 10848 15264
rect 10784 15204 10788 15260
rect 10788 15204 10844 15260
rect 10844 15204 10848 15260
rect 10784 15200 10848 15204
rect 10864 15260 10928 15264
rect 10864 15204 10868 15260
rect 10868 15204 10924 15260
rect 10924 15204 10928 15260
rect 10864 15200 10928 15204
rect 10944 15260 11008 15264
rect 10944 15204 10948 15260
rect 10948 15204 11004 15260
rect 11004 15204 11008 15260
rect 10944 15200 11008 15204
rect 2171 14716 2235 14720
rect 2171 14660 2175 14716
rect 2175 14660 2231 14716
rect 2231 14660 2235 14716
rect 2171 14656 2235 14660
rect 2251 14716 2315 14720
rect 2251 14660 2255 14716
rect 2255 14660 2311 14716
rect 2311 14660 2315 14716
rect 2251 14656 2315 14660
rect 2331 14716 2395 14720
rect 2331 14660 2335 14716
rect 2335 14660 2391 14716
rect 2391 14660 2395 14716
rect 2331 14656 2395 14660
rect 2411 14716 2475 14720
rect 2411 14660 2415 14716
rect 2415 14660 2471 14716
rect 2471 14660 2475 14716
rect 2411 14656 2475 14660
rect 4609 14716 4673 14720
rect 4609 14660 4613 14716
rect 4613 14660 4669 14716
rect 4669 14660 4673 14716
rect 4609 14656 4673 14660
rect 4689 14716 4753 14720
rect 4689 14660 4693 14716
rect 4693 14660 4749 14716
rect 4749 14660 4753 14716
rect 4689 14656 4753 14660
rect 4769 14716 4833 14720
rect 4769 14660 4773 14716
rect 4773 14660 4829 14716
rect 4829 14660 4833 14716
rect 4769 14656 4833 14660
rect 4849 14716 4913 14720
rect 4849 14660 4853 14716
rect 4853 14660 4909 14716
rect 4909 14660 4913 14716
rect 4849 14656 4913 14660
rect 7047 14716 7111 14720
rect 7047 14660 7051 14716
rect 7051 14660 7107 14716
rect 7107 14660 7111 14716
rect 7047 14656 7111 14660
rect 7127 14716 7191 14720
rect 7127 14660 7131 14716
rect 7131 14660 7187 14716
rect 7187 14660 7191 14716
rect 7127 14656 7191 14660
rect 7207 14716 7271 14720
rect 7207 14660 7211 14716
rect 7211 14660 7267 14716
rect 7267 14660 7271 14716
rect 7207 14656 7271 14660
rect 7287 14716 7351 14720
rect 7287 14660 7291 14716
rect 7291 14660 7347 14716
rect 7347 14660 7351 14716
rect 7287 14656 7351 14660
rect 9485 14716 9549 14720
rect 9485 14660 9489 14716
rect 9489 14660 9545 14716
rect 9545 14660 9549 14716
rect 9485 14656 9549 14660
rect 9565 14716 9629 14720
rect 9565 14660 9569 14716
rect 9569 14660 9625 14716
rect 9625 14660 9629 14716
rect 9565 14656 9629 14660
rect 9645 14716 9709 14720
rect 9645 14660 9649 14716
rect 9649 14660 9705 14716
rect 9705 14660 9709 14716
rect 9645 14656 9709 14660
rect 9725 14716 9789 14720
rect 9725 14660 9729 14716
rect 9729 14660 9785 14716
rect 9785 14660 9789 14716
rect 9725 14656 9789 14660
rect 3390 14172 3454 14176
rect 3390 14116 3394 14172
rect 3394 14116 3450 14172
rect 3450 14116 3454 14172
rect 3390 14112 3454 14116
rect 3470 14172 3534 14176
rect 3470 14116 3474 14172
rect 3474 14116 3530 14172
rect 3530 14116 3534 14172
rect 3470 14112 3534 14116
rect 3550 14172 3614 14176
rect 3550 14116 3554 14172
rect 3554 14116 3610 14172
rect 3610 14116 3614 14172
rect 3550 14112 3614 14116
rect 3630 14172 3694 14176
rect 3630 14116 3634 14172
rect 3634 14116 3690 14172
rect 3690 14116 3694 14172
rect 3630 14112 3694 14116
rect 5828 14172 5892 14176
rect 5828 14116 5832 14172
rect 5832 14116 5888 14172
rect 5888 14116 5892 14172
rect 5828 14112 5892 14116
rect 5908 14172 5972 14176
rect 5908 14116 5912 14172
rect 5912 14116 5968 14172
rect 5968 14116 5972 14172
rect 5908 14112 5972 14116
rect 5988 14172 6052 14176
rect 5988 14116 5992 14172
rect 5992 14116 6048 14172
rect 6048 14116 6052 14172
rect 5988 14112 6052 14116
rect 6068 14172 6132 14176
rect 6068 14116 6072 14172
rect 6072 14116 6128 14172
rect 6128 14116 6132 14172
rect 6068 14112 6132 14116
rect 8266 14172 8330 14176
rect 8266 14116 8270 14172
rect 8270 14116 8326 14172
rect 8326 14116 8330 14172
rect 8266 14112 8330 14116
rect 8346 14172 8410 14176
rect 8346 14116 8350 14172
rect 8350 14116 8406 14172
rect 8406 14116 8410 14172
rect 8346 14112 8410 14116
rect 8426 14172 8490 14176
rect 8426 14116 8430 14172
rect 8430 14116 8486 14172
rect 8486 14116 8490 14172
rect 8426 14112 8490 14116
rect 8506 14172 8570 14176
rect 8506 14116 8510 14172
rect 8510 14116 8566 14172
rect 8566 14116 8570 14172
rect 8506 14112 8570 14116
rect 10704 14172 10768 14176
rect 10704 14116 10708 14172
rect 10708 14116 10764 14172
rect 10764 14116 10768 14172
rect 10704 14112 10768 14116
rect 10784 14172 10848 14176
rect 10784 14116 10788 14172
rect 10788 14116 10844 14172
rect 10844 14116 10848 14172
rect 10784 14112 10848 14116
rect 10864 14172 10928 14176
rect 10864 14116 10868 14172
rect 10868 14116 10924 14172
rect 10924 14116 10928 14172
rect 10864 14112 10928 14116
rect 10944 14172 11008 14176
rect 10944 14116 10948 14172
rect 10948 14116 11004 14172
rect 11004 14116 11008 14172
rect 10944 14112 11008 14116
rect 2171 13628 2235 13632
rect 2171 13572 2175 13628
rect 2175 13572 2231 13628
rect 2231 13572 2235 13628
rect 2171 13568 2235 13572
rect 2251 13628 2315 13632
rect 2251 13572 2255 13628
rect 2255 13572 2311 13628
rect 2311 13572 2315 13628
rect 2251 13568 2315 13572
rect 2331 13628 2395 13632
rect 2331 13572 2335 13628
rect 2335 13572 2391 13628
rect 2391 13572 2395 13628
rect 2331 13568 2395 13572
rect 2411 13628 2475 13632
rect 2411 13572 2415 13628
rect 2415 13572 2471 13628
rect 2471 13572 2475 13628
rect 2411 13568 2475 13572
rect 4609 13628 4673 13632
rect 4609 13572 4613 13628
rect 4613 13572 4669 13628
rect 4669 13572 4673 13628
rect 4609 13568 4673 13572
rect 4689 13628 4753 13632
rect 4689 13572 4693 13628
rect 4693 13572 4749 13628
rect 4749 13572 4753 13628
rect 4689 13568 4753 13572
rect 4769 13628 4833 13632
rect 4769 13572 4773 13628
rect 4773 13572 4829 13628
rect 4829 13572 4833 13628
rect 4769 13568 4833 13572
rect 4849 13628 4913 13632
rect 4849 13572 4853 13628
rect 4853 13572 4909 13628
rect 4909 13572 4913 13628
rect 4849 13568 4913 13572
rect 7047 13628 7111 13632
rect 7047 13572 7051 13628
rect 7051 13572 7107 13628
rect 7107 13572 7111 13628
rect 7047 13568 7111 13572
rect 7127 13628 7191 13632
rect 7127 13572 7131 13628
rect 7131 13572 7187 13628
rect 7187 13572 7191 13628
rect 7127 13568 7191 13572
rect 7207 13628 7271 13632
rect 7207 13572 7211 13628
rect 7211 13572 7267 13628
rect 7267 13572 7271 13628
rect 7207 13568 7271 13572
rect 7287 13628 7351 13632
rect 7287 13572 7291 13628
rect 7291 13572 7347 13628
rect 7347 13572 7351 13628
rect 7287 13568 7351 13572
rect 9485 13628 9549 13632
rect 9485 13572 9489 13628
rect 9489 13572 9545 13628
rect 9545 13572 9549 13628
rect 9485 13568 9549 13572
rect 9565 13628 9629 13632
rect 9565 13572 9569 13628
rect 9569 13572 9625 13628
rect 9625 13572 9629 13628
rect 9565 13568 9629 13572
rect 9645 13628 9709 13632
rect 9645 13572 9649 13628
rect 9649 13572 9705 13628
rect 9705 13572 9709 13628
rect 9645 13568 9709 13572
rect 9725 13628 9789 13632
rect 9725 13572 9729 13628
rect 9729 13572 9785 13628
rect 9785 13572 9789 13628
rect 9725 13568 9789 13572
rect 3390 13084 3454 13088
rect 3390 13028 3394 13084
rect 3394 13028 3450 13084
rect 3450 13028 3454 13084
rect 3390 13024 3454 13028
rect 3470 13084 3534 13088
rect 3470 13028 3474 13084
rect 3474 13028 3530 13084
rect 3530 13028 3534 13084
rect 3470 13024 3534 13028
rect 3550 13084 3614 13088
rect 3550 13028 3554 13084
rect 3554 13028 3610 13084
rect 3610 13028 3614 13084
rect 3550 13024 3614 13028
rect 3630 13084 3694 13088
rect 3630 13028 3634 13084
rect 3634 13028 3690 13084
rect 3690 13028 3694 13084
rect 3630 13024 3694 13028
rect 5828 13084 5892 13088
rect 5828 13028 5832 13084
rect 5832 13028 5888 13084
rect 5888 13028 5892 13084
rect 5828 13024 5892 13028
rect 5908 13084 5972 13088
rect 5908 13028 5912 13084
rect 5912 13028 5968 13084
rect 5968 13028 5972 13084
rect 5908 13024 5972 13028
rect 5988 13084 6052 13088
rect 5988 13028 5992 13084
rect 5992 13028 6048 13084
rect 6048 13028 6052 13084
rect 5988 13024 6052 13028
rect 6068 13084 6132 13088
rect 6068 13028 6072 13084
rect 6072 13028 6128 13084
rect 6128 13028 6132 13084
rect 6068 13024 6132 13028
rect 8266 13084 8330 13088
rect 8266 13028 8270 13084
rect 8270 13028 8326 13084
rect 8326 13028 8330 13084
rect 8266 13024 8330 13028
rect 8346 13084 8410 13088
rect 8346 13028 8350 13084
rect 8350 13028 8406 13084
rect 8406 13028 8410 13084
rect 8346 13024 8410 13028
rect 8426 13084 8490 13088
rect 8426 13028 8430 13084
rect 8430 13028 8486 13084
rect 8486 13028 8490 13084
rect 8426 13024 8490 13028
rect 8506 13084 8570 13088
rect 8506 13028 8510 13084
rect 8510 13028 8566 13084
rect 8566 13028 8570 13084
rect 8506 13024 8570 13028
rect 10704 13084 10768 13088
rect 10704 13028 10708 13084
rect 10708 13028 10764 13084
rect 10764 13028 10768 13084
rect 10704 13024 10768 13028
rect 10784 13084 10848 13088
rect 10784 13028 10788 13084
rect 10788 13028 10844 13084
rect 10844 13028 10848 13084
rect 10784 13024 10848 13028
rect 10864 13084 10928 13088
rect 10864 13028 10868 13084
rect 10868 13028 10924 13084
rect 10924 13028 10928 13084
rect 10864 13024 10928 13028
rect 10944 13084 11008 13088
rect 10944 13028 10948 13084
rect 10948 13028 11004 13084
rect 11004 13028 11008 13084
rect 10944 13024 11008 13028
rect 2171 12540 2235 12544
rect 2171 12484 2175 12540
rect 2175 12484 2231 12540
rect 2231 12484 2235 12540
rect 2171 12480 2235 12484
rect 2251 12540 2315 12544
rect 2251 12484 2255 12540
rect 2255 12484 2311 12540
rect 2311 12484 2315 12540
rect 2251 12480 2315 12484
rect 2331 12540 2395 12544
rect 2331 12484 2335 12540
rect 2335 12484 2391 12540
rect 2391 12484 2395 12540
rect 2331 12480 2395 12484
rect 2411 12540 2475 12544
rect 2411 12484 2415 12540
rect 2415 12484 2471 12540
rect 2471 12484 2475 12540
rect 2411 12480 2475 12484
rect 4609 12540 4673 12544
rect 4609 12484 4613 12540
rect 4613 12484 4669 12540
rect 4669 12484 4673 12540
rect 4609 12480 4673 12484
rect 4689 12540 4753 12544
rect 4689 12484 4693 12540
rect 4693 12484 4749 12540
rect 4749 12484 4753 12540
rect 4689 12480 4753 12484
rect 4769 12540 4833 12544
rect 4769 12484 4773 12540
rect 4773 12484 4829 12540
rect 4829 12484 4833 12540
rect 4769 12480 4833 12484
rect 4849 12540 4913 12544
rect 4849 12484 4853 12540
rect 4853 12484 4909 12540
rect 4909 12484 4913 12540
rect 4849 12480 4913 12484
rect 7047 12540 7111 12544
rect 7047 12484 7051 12540
rect 7051 12484 7107 12540
rect 7107 12484 7111 12540
rect 7047 12480 7111 12484
rect 7127 12540 7191 12544
rect 7127 12484 7131 12540
rect 7131 12484 7187 12540
rect 7187 12484 7191 12540
rect 7127 12480 7191 12484
rect 7207 12540 7271 12544
rect 7207 12484 7211 12540
rect 7211 12484 7267 12540
rect 7267 12484 7271 12540
rect 7207 12480 7271 12484
rect 7287 12540 7351 12544
rect 7287 12484 7291 12540
rect 7291 12484 7347 12540
rect 7347 12484 7351 12540
rect 7287 12480 7351 12484
rect 9485 12540 9549 12544
rect 9485 12484 9489 12540
rect 9489 12484 9545 12540
rect 9545 12484 9549 12540
rect 9485 12480 9549 12484
rect 9565 12540 9629 12544
rect 9565 12484 9569 12540
rect 9569 12484 9625 12540
rect 9625 12484 9629 12540
rect 9565 12480 9629 12484
rect 9645 12540 9709 12544
rect 9645 12484 9649 12540
rect 9649 12484 9705 12540
rect 9705 12484 9709 12540
rect 9645 12480 9709 12484
rect 9725 12540 9789 12544
rect 9725 12484 9729 12540
rect 9729 12484 9785 12540
rect 9785 12484 9789 12540
rect 9725 12480 9789 12484
rect 3390 11996 3454 12000
rect 3390 11940 3394 11996
rect 3394 11940 3450 11996
rect 3450 11940 3454 11996
rect 3390 11936 3454 11940
rect 3470 11996 3534 12000
rect 3470 11940 3474 11996
rect 3474 11940 3530 11996
rect 3530 11940 3534 11996
rect 3470 11936 3534 11940
rect 3550 11996 3614 12000
rect 3550 11940 3554 11996
rect 3554 11940 3610 11996
rect 3610 11940 3614 11996
rect 3550 11936 3614 11940
rect 3630 11996 3694 12000
rect 3630 11940 3634 11996
rect 3634 11940 3690 11996
rect 3690 11940 3694 11996
rect 3630 11936 3694 11940
rect 5828 11996 5892 12000
rect 5828 11940 5832 11996
rect 5832 11940 5888 11996
rect 5888 11940 5892 11996
rect 5828 11936 5892 11940
rect 5908 11996 5972 12000
rect 5908 11940 5912 11996
rect 5912 11940 5968 11996
rect 5968 11940 5972 11996
rect 5908 11936 5972 11940
rect 5988 11996 6052 12000
rect 5988 11940 5992 11996
rect 5992 11940 6048 11996
rect 6048 11940 6052 11996
rect 5988 11936 6052 11940
rect 6068 11996 6132 12000
rect 6068 11940 6072 11996
rect 6072 11940 6128 11996
rect 6128 11940 6132 11996
rect 6068 11936 6132 11940
rect 8266 11996 8330 12000
rect 8266 11940 8270 11996
rect 8270 11940 8326 11996
rect 8326 11940 8330 11996
rect 8266 11936 8330 11940
rect 8346 11996 8410 12000
rect 8346 11940 8350 11996
rect 8350 11940 8406 11996
rect 8406 11940 8410 11996
rect 8346 11936 8410 11940
rect 8426 11996 8490 12000
rect 8426 11940 8430 11996
rect 8430 11940 8486 11996
rect 8486 11940 8490 11996
rect 8426 11936 8490 11940
rect 8506 11996 8570 12000
rect 8506 11940 8510 11996
rect 8510 11940 8566 11996
rect 8566 11940 8570 11996
rect 8506 11936 8570 11940
rect 10704 11996 10768 12000
rect 10704 11940 10708 11996
rect 10708 11940 10764 11996
rect 10764 11940 10768 11996
rect 10704 11936 10768 11940
rect 10784 11996 10848 12000
rect 10784 11940 10788 11996
rect 10788 11940 10844 11996
rect 10844 11940 10848 11996
rect 10784 11936 10848 11940
rect 10864 11996 10928 12000
rect 10864 11940 10868 11996
rect 10868 11940 10924 11996
rect 10924 11940 10928 11996
rect 10864 11936 10928 11940
rect 10944 11996 11008 12000
rect 10944 11940 10948 11996
rect 10948 11940 11004 11996
rect 11004 11940 11008 11996
rect 10944 11936 11008 11940
rect 2171 11452 2235 11456
rect 2171 11396 2175 11452
rect 2175 11396 2231 11452
rect 2231 11396 2235 11452
rect 2171 11392 2235 11396
rect 2251 11452 2315 11456
rect 2251 11396 2255 11452
rect 2255 11396 2311 11452
rect 2311 11396 2315 11452
rect 2251 11392 2315 11396
rect 2331 11452 2395 11456
rect 2331 11396 2335 11452
rect 2335 11396 2391 11452
rect 2391 11396 2395 11452
rect 2331 11392 2395 11396
rect 2411 11452 2475 11456
rect 2411 11396 2415 11452
rect 2415 11396 2471 11452
rect 2471 11396 2475 11452
rect 2411 11392 2475 11396
rect 4609 11452 4673 11456
rect 4609 11396 4613 11452
rect 4613 11396 4669 11452
rect 4669 11396 4673 11452
rect 4609 11392 4673 11396
rect 4689 11452 4753 11456
rect 4689 11396 4693 11452
rect 4693 11396 4749 11452
rect 4749 11396 4753 11452
rect 4689 11392 4753 11396
rect 4769 11452 4833 11456
rect 4769 11396 4773 11452
rect 4773 11396 4829 11452
rect 4829 11396 4833 11452
rect 4769 11392 4833 11396
rect 4849 11452 4913 11456
rect 4849 11396 4853 11452
rect 4853 11396 4909 11452
rect 4909 11396 4913 11452
rect 4849 11392 4913 11396
rect 7047 11452 7111 11456
rect 7047 11396 7051 11452
rect 7051 11396 7107 11452
rect 7107 11396 7111 11452
rect 7047 11392 7111 11396
rect 7127 11452 7191 11456
rect 7127 11396 7131 11452
rect 7131 11396 7187 11452
rect 7187 11396 7191 11452
rect 7127 11392 7191 11396
rect 7207 11452 7271 11456
rect 7207 11396 7211 11452
rect 7211 11396 7267 11452
rect 7267 11396 7271 11452
rect 7207 11392 7271 11396
rect 7287 11452 7351 11456
rect 7287 11396 7291 11452
rect 7291 11396 7347 11452
rect 7347 11396 7351 11452
rect 7287 11392 7351 11396
rect 9485 11452 9549 11456
rect 9485 11396 9489 11452
rect 9489 11396 9545 11452
rect 9545 11396 9549 11452
rect 9485 11392 9549 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 3390 10908 3454 10912
rect 3390 10852 3394 10908
rect 3394 10852 3450 10908
rect 3450 10852 3454 10908
rect 3390 10848 3454 10852
rect 3470 10908 3534 10912
rect 3470 10852 3474 10908
rect 3474 10852 3530 10908
rect 3530 10852 3534 10908
rect 3470 10848 3534 10852
rect 3550 10908 3614 10912
rect 3550 10852 3554 10908
rect 3554 10852 3610 10908
rect 3610 10852 3614 10908
rect 3550 10848 3614 10852
rect 3630 10908 3694 10912
rect 3630 10852 3634 10908
rect 3634 10852 3690 10908
rect 3690 10852 3694 10908
rect 3630 10848 3694 10852
rect 5828 10908 5892 10912
rect 5828 10852 5832 10908
rect 5832 10852 5888 10908
rect 5888 10852 5892 10908
rect 5828 10848 5892 10852
rect 5908 10908 5972 10912
rect 5908 10852 5912 10908
rect 5912 10852 5968 10908
rect 5968 10852 5972 10908
rect 5908 10848 5972 10852
rect 5988 10908 6052 10912
rect 5988 10852 5992 10908
rect 5992 10852 6048 10908
rect 6048 10852 6052 10908
rect 5988 10848 6052 10852
rect 6068 10908 6132 10912
rect 6068 10852 6072 10908
rect 6072 10852 6128 10908
rect 6128 10852 6132 10908
rect 6068 10848 6132 10852
rect 8266 10908 8330 10912
rect 8266 10852 8270 10908
rect 8270 10852 8326 10908
rect 8326 10852 8330 10908
rect 8266 10848 8330 10852
rect 8346 10908 8410 10912
rect 8346 10852 8350 10908
rect 8350 10852 8406 10908
rect 8406 10852 8410 10908
rect 8346 10848 8410 10852
rect 8426 10908 8490 10912
rect 8426 10852 8430 10908
rect 8430 10852 8486 10908
rect 8486 10852 8490 10908
rect 8426 10848 8490 10852
rect 8506 10908 8570 10912
rect 8506 10852 8510 10908
rect 8510 10852 8566 10908
rect 8566 10852 8570 10908
rect 8506 10848 8570 10852
rect 10704 10908 10768 10912
rect 10704 10852 10708 10908
rect 10708 10852 10764 10908
rect 10764 10852 10768 10908
rect 10704 10848 10768 10852
rect 10784 10908 10848 10912
rect 10784 10852 10788 10908
rect 10788 10852 10844 10908
rect 10844 10852 10848 10908
rect 10784 10848 10848 10852
rect 10864 10908 10928 10912
rect 10864 10852 10868 10908
rect 10868 10852 10924 10908
rect 10924 10852 10928 10908
rect 10864 10848 10928 10852
rect 10944 10908 11008 10912
rect 10944 10852 10948 10908
rect 10948 10852 11004 10908
rect 11004 10852 11008 10908
rect 10944 10848 11008 10852
rect 2171 10364 2235 10368
rect 2171 10308 2175 10364
rect 2175 10308 2231 10364
rect 2231 10308 2235 10364
rect 2171 10304 2235 10308
rect 2251 10364 2315 10368
rect 2251 10308 2255 10364
rect 2255 10308 2311 10364
rect 2311 10308 2315 10364
rect 2251 10304 2315 10308
rect 2331 10364 2395 10368
rect 2331 10308 2335 10364
rect 2335 10308 2391 10364
rect 2391 10308 2395 10364
rect 2331 10304 2395 10308
rect 2411 10364 2475 10368
rect 2411 10308 2415 10364
rect 2415 10308 2471 10364
rect 2471 10308 2475 10364
rect 2411 10304 2475 10308
rect 4609 10364 4673 10368
rect 4609 10308 4613 10364
rect 4613 10308 4669 10364
rect 4669 10308 4673 10364
rect 4609 10304 4673 10308
rect 4689 10364 4753 10368
rect 4689 10308 4693 10364
rect 4693 10308 4749 10364
rect 4749 10308 4753 10364
rect 4689 10304 4753 10308
rect 4769 10364 4833 10368
rect 4769 10308 4773 10364
rect 4773 10308 4829 10364
rect 4829 10308 4833 10364
rect 4769 10304 4833 10308
rect 4849 10364 4913 10368
rect 4849 10308 4853 10364
rect 4853 10308 4909 10364
rect 4909 10308 4913 10364
rect 4849 10304 4913 10308
rect 7047 10364 7111 10368
rect 7047 10308 7051 10364
rect 7051 10308 7107 10364
rect 7107 10308 7111 10364
rect 7047 10304 7111 10308
rect 7127 10364 7191 10368
rect 7127 10308 7131 10364
rect 7131 10308 7187 10364
rect 7187 10308 7191 10364
rect 7127 10304 7191 10308
rect 7207 10364 7271 10368
rect 7207 10308 7211 10364
rect 7211 10308 7267 10364
rect 7267 10308 7271 10364
rect 7207 10304 7271 10308
rect 7287 10364 7351 10368
rect 7287 10308 7291 10364
rect 7291 10308 7347 10364
rect 7347 10308 7351 10364
rect 7287 10304 7351 10308
rect 9485 10364 9549 10368
rect 9485 10308 9489 10364
rect 9489 10308 9545 10364
rect 9545 10308 9549 10364
rect 9485 10304 9549 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 15808 2483 15824
rect 2163 15744 2171 15808
rect 2235 15744 2251 15808
rect 2315 15744 2331 15808
rect 2395 15744 2411 15808
rect 2475 15744 2483 15808
rect 2163 14720 2483 15744
rect 2163 14656 2171 14720
rect 2235 14656 2251 14720
rect 2315 14656 2331 14720
rect 2395 14656 2411 14720
rect 2475 14656 2483 14720
rect 2163 13632 2483 14656
rect 2163 13568 2171 13632
rect 2235 13568 2251 13632
rect 2315 13568 2331 13632
rect 2395 13568 2411 13632
rect 2475 13568 2483 13632
rect 2163 12544 2483 13568
rect 2163 12480 2171 12544
rect 2235 12480 2251 12544
rect 2315 12480 2331 12544
rect 2395 12480 2411 12544
rect 2475 12480 2483 12544
rect 2163 11456 2483 12480
rect 2163 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2483 11456
rect 2163 10368 2483 11392
rect 2163 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2483 10368
rect 2163 9280 2483 10304
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 15264 3702 15824
rect 3382 15200 3390 15264
rect 3454 15200 3470 15264
rect 3534 15200 3550 15264
rect 3614 15200 3630 15264
rect 3694 15200 3702 15264
rect 3382 14176 3702 15200
rect 3382 14112 3390 14176
rect 3454 14112 3470 14176
rect 3534 14112 3550 14176
rect 3614 14112 3630 14176
rect 3694 14112 3702 14176
rect 3382 13088 3702 14112
rect 3382 13024 3390 13088
rect 3454 13024 3470 13088
rect 3534 13024 3550 13088
rect 3614 13024 3630 13088
rect 3694 13024 3702 13088
rect 3382 12000 3702 13024
rect 3382 11936 3390 12000
rect 3454 11936 3470 12000
rect 3534 11936 3550 12000
rect 3614 11936 3630 12000
rect 3694 11936 3702 12000
rect 3382 10912 3702 11936
rect 3382 10848 3390 10912
rect 3454 10848 3470 10912
rect 3534 10848 3550 10912
rect 3614 10848 3630 10912
rect 3694 10848 3702 10912
rect 3382 9824 3702 10848
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 15808 4921 15824
rect 4601 15744 4609 15808
rect 4673 15744 4689 15808
rect 4753 15744 4769 15808
rect 4833 15744 4849 15808
rect 4913 15744 4921 15808
rect 4601 14720 4921 15744
rect 4601 14656 4609 14720
rect 4673 14656 4689 14720
rect 4753 14656 4769 14720
rect 4833 14656 4849 14720
rect 4913 14656 4921 14720
rect 4601 13632 4921 14656
rect 4601 13568 4609 13632
rect 4673 13568 4689 13632
rect 4753 13568 4769 13632
rect 4833 13568 4849 13632
rect 4913 13568 4921 13632
rect 4601 12544 4921 13568
rect 4601 12480 4609 12544
rect 4673 12480 4689 12544
rect 4753 12480 4769 12544
rect 4833 12480 4849 12544
rect 4913 12480 4921 12544
rect 4601 11456 4921 12480
rect 4601 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4921 11456
rect 4601 10368 4921 11392
rect 4601 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4921 10368
rect 4601 9280 4921 10304
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 15264 6140 15824
rect 5820 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6140 15264
rect 5820 14176 6140 15200
rect 5820 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6140 14176
rect 5820 13088 6140 14112
rect 5820 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6140 13088
rect 5820 12000 6140 13024
rect 5820 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6140 12000
rect 5820 10912 6140 11936
rect 5820 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6140 10912
rect 5820 9824 6140 10848
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 15808 7359 15824
rect 7039 15744 7047 15808
rect 7111 15744 7127 15808
rect 7191 15744 7207 15808
rect 7271 15744 7287 15808
rect 7351 15744 7359 15808
rect 7039 14720 7359 15744
rect 7039 14656 7047 14720
rect 7111 14656 7127 14720
rect 7191 14656 7207 14720
rect 7271 14656 7287 14720
rect 7351 14656 7359 14720
rect 7039 13632 7359 14656
rect 7039 13568 7047 13632
rect 7111 13568 7127 13632
rect 7191 13568 7207 13632
rect 7271 13568 7287 13632
rect 7351 13568 7359 13632
rect 7039 12544 7359 13568
rect 7039 12480 7047 12544
rect 7111 12480 7127 12544
rect 7191 12480 7207 12544
rect 7271 12480 7287 12544
rect 7351 12480 7359 12544
rect 7039 11456 7359 12480
rect 7039 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7359 11456
rect 7039 10368 7359 11392
rect 7039 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7359 10368
rect 7039 9280 7359 10304
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 15264 8578 15824
rect 8258 15200 8266 15264
rect 8330 15200 8346 15264
rect 8410 15200 8426 15264
rect 8490 15200 8506 15264
rect 8570 15200 8578 15264
rect 8258 14176 8578 15200
rect 8258 14112 8266 14176
rect 8330 14112 8346 14176
rect 8410 14112 8426 14176
rect 8490 14112 8506 14176
rect 8570 14112 8578 14176
rect 8258 13088 8578 14112
rect 8258 13024 8266 13088
rect 8330 13024 8346 13088
rect 8410 13024 8426 13088
rect 8490 13024 8506 13088
rect 8570 13024 8578 13088
rect 8258 12000 8578 13024
rect 8258 11936 8266 12000
rect 8330 11936 8346 12000
rect 8410 11936 8426 12000
rect 8490 11936 8506 12000
rect 8570 11936 8578 12000
rect 8258 10912 8578 11936
rect 8258 10848 8266 10912
rect 8330 10848 8346 10912
rect 8410 10848 8426 10912
rect 8490 10848 8506 10912
rect 8570 10848 8578 10912
rect 8258 9824 8578 10848
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 15808 9797 15824
rect 9477 15744 9485 15808
rect 9549 15744 9565 15808
rect 9629 15744 9645 15808
rect 9709 15744 9725 15808
rect 9789 15744 9797 15808
rect 9477 14720 9797 15744
rect 9477 14656 9485 14720
rect 9549 14656 9565 14720
rect 9629 14656 9645 14720
rect 9709 14656 9725 14720
rect 9789 14656 9797 14720
rect 9477 13632 9797 14656
rect 9477 13568 9485 13632
rect 9549 13568 9565 13632
rect 9629 13568 9645 13632
rect 9709 13568 9725 13632
rect 9789 13568 9797 13632
rect 9477 12544 9797 13568
rect 9477 12480 9485 12544
rect 9549 12480 9565 12544
rect 9629 12480 9645 12544
rect 9709 12480 9725 12544
rect 9789 12480 9797 12544
rect 9477 11456 9797 12480
rect 9477 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9797 11456
rect 9477 10368 9797 11392
rect 9477 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9797 10368
rect 9477 9280 9797 10304
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 15264 11016 15824
rect 10696 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11016 15264
rect 10696 14176 11016 15200
rect 10696 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11016 14176
rect 10696 13088 11016 14112
rect 10696 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11016 13088
rect 10696 12000 11016 13024
rect 10696 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11016 12000
rect 10696 10912 11016 11936
rect 10696 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11016 10912
rect 10696 9824 11016 10848
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1676037725
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67
timestamp 1676037725
transform 1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1676037725
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_18
timestamp 1676037725
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_37
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_36
timestamp 1676037725
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1676037725
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_63
timestamp 1676037725
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1676037725
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_94
timestamp 1676037725
transform 1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1676037725
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_30
timestamp 1676037725
transform 1 0 3864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_41
timestamp 1676037725
transform 1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1676037725
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1676037725
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_84
timestamp 1676037725
transform 1 0 8832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_96
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1676037725
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_19
timestamp 1676037725
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1676037725
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_38
timestamp 1676037725
transform 1 0 4600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1676037725
transform 1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_54
timestamp 1676037725
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_71
timestamp 1676037725
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 1676037725
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_16
timestamp 1676037725
transform 1 0 2576 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1676037725
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_14
timestamp 1676037725
transform 1 0 2392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_49
timestamp 1676037725
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_61
timestamp 1676037725
transform 1 0 6716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1676037725
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1676037725
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_13
timestamp 1676037725
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_25
timestamp 1676037725
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp 1676037725
transform 1 0 4876 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1676037725
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1676037725
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1676037725
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_79
timestamp 1676037725
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1676037725
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1676037725
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1676037725
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1676037725
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1676037725
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1676037725
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1676037725
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_72
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_84
timestamp 1676037725
transform 1 0 8832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_96
timestamp 1676037725
transform 1 0 9936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1676037725
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_50
timestamp 1676037725
transform 1 0 5704 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_62
timestamp 1676037725
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_20
timestamp 1676037725
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1676037725
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_7
timestamp 1676037725
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1676037725
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_71
timestamp 1676037725
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1676037725
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_39
timestamp 1676037725
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_51
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_63
timestamp 1676037725
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1676037725
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1676037725
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_77
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_89
timestamp 1676037725
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1676037725
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1676037725
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1676037725
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_62
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_74
timestamp 1676037725
transform 1 0 7912 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_86
timestamp 1676037725
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1676037725
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_102
timestamp 1676037725
transform 1 0 10488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1676037725
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1676037725
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1676037725
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1676037725
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_7
timestamp 1676037725
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_19
timestamp 1676037725
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1676037725
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1676037725
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp 1676037725
transform -1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _057_
timestamp 1676037725
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _060_
timestamp 1676037725
transform -1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_4  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__a21o_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3864 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _067_
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _068_
timestamp 1676037725
transform 1 0 2852 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _069_
timestamp 1676037725
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7728 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _071_
timestamp 1676037725
transform -1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3128 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__nand3_2  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _076_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _078_
timestamp 1676037725
transform 1 0 5152 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _080_
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5704 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _082_
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _083_
timestamp 1676037725
transform -1 0 3496 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _086_
timestamp 1676037725
transform 1 0 5152 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _087_
timestamp 1676037725
transform -1 0 5520 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _089_
timestamp 1676037725
transform 1 0 3680 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _090_
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4784 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_2  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6072 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _095_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _099_
timestamp 1676037725
transform -1 0 7544 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1676037725
transform -1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _101_
timestamp 1676037725
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _102_
timestamp 1676037725
transform -1 0 6072 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _103_
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _104_
timestamp 1676037725
transform 1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _105_
timestamp 1676037725
transform 1 0 6992 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _106_
timestamp 1676037725
transform 1 0 8004 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 1676037725
transform -1 0 7912 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _108_
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _109_
timestamp 1676037725
transform -1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _111_
timestamp 1676037725
transform -1 0 8832 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1676037725
transform -1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform -1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 9844 0 -1 3264
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_in[3]
port 3 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 io_in[6]
port 6 nsew signal input
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 io_in[7]
port 7 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 2163 2128 2483 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 4601 2128 4921 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7039 2128 7359 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 9477 2128 9797 15824 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 3382 2128 3702 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 15824 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 18000
<< end >>
