magic
tech sky130B
magscale 1 2
timestamp 1676307443
<< obsli1 >>
rect 1104 2159 54832 53329
<< obsm1 >>
rect 1104 1980 54832 53360
<< metal2 >>
rect 1674 55200 1730 56000
rect 2870 55200 2926 56000
rect 4066 55200 4122 56000
rect 5262 55200 5318 56000
rect 6458 55200 6514 56000
rect 7654 55200 7710 56000
rect 8850 55200 8906 56000
rect 10046 55200 10102 56000
rect 11242 55200 11298 56000
rect 12438 55200 12494 56000
rect 13634 55200 13690 56000
rect 14830 55200 14886 56000
rect 16026 55200 16082 56000
rect 17222 55200 17278 56000
rect 18418 55200 18474 56000
rect 19614 55200 19670 56000
rect 20810 55200 20866 56000
rect 22006 55200 22062 56000
rect 23202 55200 23258 56000
rect 24398 55200 24454 56000
rect 25594 55200 25650 56000
rect 26790 55200 26846 56000
rect 27986 55200 28042 56000
rect 29182 55200 29238 56000
rect 30378 55200 30434 56000
rect 31574 55200 31630 56000
rect 32770 55200 32826 56000
rect 33966 55200 34022 56000
rect 35162 55200 35218 56000
rect 36358 55200 36414 56000
rect 37554 55200 37610 56000
rect 38750 55200 38806 56000
rect 39946 55200 40002 56000
rect 41142 55200 41198 56000
rect 42338 55200 42394 56000
rect 43534 55200 43590 56000
rect 44730 55200 44786 56000
rect 45926 55200 45982 56000
rect 47122 55200 47178 56000
rect 48318 55200 48374 56000
rect 49514 55200 49570 56000
rect 50710 55200 50766 56000
rect 51906 55200 51962 56000
rect 53102 55200 53158 56000
rect 54298 55200 54354 56000
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50986 0 51042 800
<< obsm2 >>
rect 1490 55144 1618 55298
rect 1786 55144 2814 55298
rect 2982 55144 4010 55298
rect 4178 55144 5206 55298
rect 5374 55144 6402 55298
rect 6570 55144 7598 55298
rect 7766 55144 8794 55298
rect 8962 55144 9990 55298
rect 10158 55144 11186 55298
rect 11354 55144 12382 55298
rect 12550 55144 13578 55298
rect 13746 55144 14774 55298
rect 14942 55144 15970 55298
rect 16138 55144 17166 55298
rect 17334 55144 18362 55298
rect 18530 55144 19558 55298
rect 19726 55144 20754 55298
rect 20922 55144 21950 55298
rect 22118 55144 23146 55298
rect 23314 55144 24342 55298
rect 24510 55144 25538 55298
rect 25706 55144 26734 55298
rect 26902 55144 27930 55298
rect 28098 55144 29126 55298
rect 29294 55144 30322 55298
rect 30490 55144 31518 55298
rect 31686 55144 32714 55298
rect 32882 55144 33910 55298
rect 34078 55144 35106 55298
rect 35274 55144 36302 55298
rect 36470 55144 37498 55298
rect 37666 55144 38694 55298
rect 38862 55144 39890 55298
rect 40058 55144 41086 55298
rect 41254 55144 42282 55298
rect 42450 55144 43478 55298
rect 43646 55144 44674 55298
rect 44842 55144 45870 55298
rect 46038 55144 47066 55298
rect 47234 55144 48262 55298
rect 48430 55144 49458 55298
rect 49626 55144 50654 55298
rect 50822 55144 51850 55298
rect 52018 55144 53046 55298
rect 53214 55144 54242 55298
rect 54410 55144 54538 55298
rect 1490 856 54538 55144
rect 1490 734 4930 856
rect 5098 734 5298 856
rect 5466 734 5666 856
rect 5834 734 6034 856
rect 6202 734 6402 856
rect 6570 734 6770 856
rect 6938 734 7138 856
rect 7306 734 7506 856
rect 7674 734 7874 856
rect 8042 734 8242 856
rect 8410 734 8610 856
rect 8778 734 8978 856
rect 9146 734 9346 856
rect 9514 734 9714 856
rect 9882 734 10082 856
rect 10250 734 10450 856
rect 10618 734 10818 856
rect 10986 734 11186 856
rect 11354 734 11554 856
rect 11722 734 11922 856
rect 12090 734 12290 856
rect 12458 734 12658 856
rect 12826 734 13026 856
rect 13194 734 13394 856
rect 13562 734 13762 856
rect 13930 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14866 856
rect 15034 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15970 856
rect 16138 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17810 856
rect 17978 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18914 856
rect 19082 734 19282 856
rect 19450 734 19650 856
rect 19818 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20754 856
rect 20922 734 21122 856
rect 21290 734 21490 856
rect 21658 734 21858 856
rect 22026 734 22226 856
rect 22394 734 22594 856
rect 22762 734 22962 856
rect 23130 734 23330 856
rect 23498 734 23698 856
rect 23866 734 24066 856
rect 24234 734 24434 856
rect 24602 734 24802 856
rect 24970 734 25170 856
rect 25338 734 25538 856
rect 25706 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 27010 856
rect 27178 734 27378 856
rect 27546 734 27746 856
rect 27914 734 28114 856
rect 28282 734 28482 856
rect 28650 734 28850 856
rect 29018 734 29218 856
rect 29386 734 29586 856
rect 29754 734 29954 856
rect 30122 734 30322 856
rect 30490 734 30690 856
rect 30858 734 31058 856
rect 31226 734 31426 856
rect 31594 734 31794 856
rect 31962 734 32162 856
rect 32330 734 32530 856
rect 32698 734 32898 856
rect 33066 734 33266 856
rect 33434 734 33634 856
rect 33802 734 34002 856
rect 34170 734 34370 856
rect 34538 734 34738 856
rect 34906 734 35106 856
rect 35274 734 35474 856
rect 35642 734 35842 856
rect 36010 734 36210 856
rect 36378 734 36578 856
rect 36746 734 36946 856
rect 37114 734 37314 856
rect 37482 734 37682 856
rect 37850 734 38050 856
rect 38218 734 38418 856
rect 38586 734 38786 856
rect 38954 734 39154 856
rect 39322 734 39522 856
rect 39690 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40626 856
rect 40794 734 40994 856
rect 41162 734 41362 856
rect 41530 734 41730 856
rect 41898 734 42098 856
rect 42266 734 42466 856
rect 42634 734 42834 856
rect 43002 734 43202 856
rect 43370 734 43570 856
rect 43738 734 43938 856
rect 44106 734 44306 856
rect 44474 734 44674 856
rect 44842 734 45042 856
rect 45210 734 45410 856
rect 45578 734 45778 856
rect 45946 734 46146 856
rect 46314 734 46514 856
rect 46682 734 46882 856
rect 47050 734 47250 856
rect 47418 734 47618 856
rect 47786 734 47986 856
rect 48154 734 48354 856
rect 48522 734 48722 856
rect 48890 734 49090 856
rect 49258 734 49458 856
rect 49626 734 49826 856
rect 49994 734 50194 856
rect 50362 734 50562 856
rect 50730 734 50930 856
rect 51098 734 54538 856
<< metal3 >>
rect 0 52640 800 52760
rect 0 52096 800 52216
rect 0 51552 800 51672
rect 0 51008 800 51128
rect 0 50464 800 50584
rect 0 49920 800 50040
rect 0 49376 800 49496
rect 55200 49240 56000 49360
rect 0 48832 800 48952
rect 55200 48968 56000 49088
rect 55200 48696 56000 48816
rect 0 48288 800 48408
rect 55200 48424 56000 48544
rect 55200 48152 56000 48272
rect 0 47744 800 47864
rect 55200 47880 56000 48000
rect 55200 47608 56000 47728
rect 0 47200 800 47320
rect 55200 47336 56000 47456
rect 55200 47064 56000 47184
rect 0 46656 800 46776
rect 55200 46792 56000 46912
rect 55200 46520 56000 46640
rect 0 46112 800 46232
rect 55200 46248 56000 46368
rect 55200 45976 56000 46096
rect 0 45568 800 45688
rect 55200 45704 56000 45824
rect 55200 45432 56000 45552
rect 0 45024 800 45144
rect 55200 45160 56000 45280
rect 55200 44888 56000 45008
rect 0 44480 800 44600
rect 55200 44616 56000 44736
rect 55200 44344 56000 44464
rect 0 43936 800 44056
rect 55200 44072 56000 44192
rect 55200 43800 56000 43920
rect 0 43392 800 43512
rect 55200 43528 56000 43648
rect 55200 43256 56000 43376
rect 0 42848 800 42968
rect 55200 42984 56000 43104
rect 55200 42712 56000 42832
rect 0 42304 800 42424
rect 55200 42440 56000 42560
rect 55200 42168 56000 42288
rect 0 41760 800 41880
rect 55200 41896 56000 42016
rect 55200 41624 56000 41744
rect 0 41216 800 41336
rect 55200 41352 56000 41472
rect 55200 41080 56000 41200
rect 0 40672 800 40792
rect 55200 40808 56000 40928
rect 55200 40536 56000 40656
rect 0 40128 800 40248
rect 55200 40264 56000 40384
rect 55200 39992 56000 40112
rect 0 39584 800 39704
rect 55200 39720 56000 39840
rect 55200 39448 56000 39568
rect 0 39040 800 39160
rect 55200 39176 56000 39296
rect 55200 38904 56000 39024
rect 0 38496 800 38616
rect 55200 38632 56000 38752
rect 55200 38360 56000 38480
rect 0 37952 800 38072
rect 55200 38088 56000 38208
rect 55200 37816 56000 37936
rect 0 37408 800 37528
rect 55200 37544 56000 37664
rect 55200 37272 56000 37392
rect 0 36864 800 36984
rect 55200 37000 56000 37120
rect 55200 36728 56000 36848
rect 0 36320 800 36440
rect 55200 36456 56000 36576
rect 55200 36184 56000 36304
rect 0 35776 800 35896
rect 55200 35912 56000 36032
rect 55200 35640 56000 35760
rect 0 35232 800 35352
rect 55200 35368 56000 35488
rect 55200 35096 56000 35216
rect 0 34688 800 34808
rect 55200 34824 56000 34944
rect 55200 34552 56000 34672
rect 0 34144 800 34264
rect 55200 34280 56000 34400
rect 55200 34008 56000 34128
rect 0 33600 800 33720
rect 55200 33736 56000 33856
rect 55200 33464 56000 33584
rect 0 33056 800 33176
rect 55200 33192 56000 33312
rect 55200 32920 56000 33040
rect 0 32512 800 32632
rect 55200 32648 56000 32768
rect 55200 32376 56000 32496
rect 0 31968 800 32088
rect 55200 32104 56000 32224
rect 55200 31832 56000 31952
rect 0 31424 800 31544
rect 55200 31560 56000 31680
rect 55200 31288 56000 31408
rect 0 30880 800 31000
rect 55200 31016 56000 31136
rect 55200 30744 56000 30864
rect 0 30336 800 30456
rect 55200 30472 56000 30592
rect 55200 30200 56000 30320
rect 0 29792 800 29912
rect 55200 29928 56000 30048
rect 55200 29656 56000 29776
rect 0 29248 800 29368
rect 55200 29384 56000 29504
rect 55200 29112 56000 29232
rect 0 28704 800 28824
rect 55200 28840 56000 28960
rect 55200 28568 56000 28688
rect 0 28160 800 28280
rect 55200 28296 56000 28416
rect 55200 28024 56000 28144
rect 0 27616 800 27736
rect 55200 27752 56000 27872
rect 55200 27480 56000 27600
rect 0 27072 800 27192
rect 55200 27208 56000 27328
rect 55200 26936 56000 27056
rect 0 26528 800 26648
rect 55200 26664 56000 26784
rect 55200 26392 56000 26512
rect 0 25984 800 26104
rect 55200 26120 56000 26240
rect 55200 25848 56000 25968
rect 0 25440 800 25560
rect 55200 25576 56000 25696
rect 55200 25304 56000 25424
rect 0 24896 800 25016
rect 55200 25032 56000 25152
rect 55200 24760 56000 24880
rect 0 24352 800 24472
rect 55200 24488 56000 24608
rect 55200 24216 56000 24336
rect 0 23808 800 23928
rect 55200 23944 56000 24064
rect 55200 23672 56000 23792
rect 0 23264 800 23384
rect 55200 23400 56000 23520
rect 55200 23128 56000 23248
rect 0 22720 800 22840
rect 55200 22856 56000 22976
rect 55200 22584 56000 22704
rect 0 22176 800 22296
rect 55200 22312 56000 22432
rect 55200 22040 56000 22160
rect 0 21632 800 21752
rect 55200 21768 56000 21888
rect 55200 21496 56000 21616
rect 0 21088 800 21208
rect 55200 21224 56000 21344
rect 55200 20952 56000 21072
rect 0 20544 800 20664
rect 55200 20680 56000 20800
rect 55200 20408 56000 20528
rect 0 20000 800 20120
rect 55200 20136 56000 20256
rect 55200 19864 56000 19984
rect 0 19456 800 19576
rect 55200 19592 56000 19712
rect 55200 19320 56000 19440
rect 0 18912 800 19032
rect 55200 19048 56000 19168
rect 55200 18776 56000 18896
rect 0 18368 800 18488
rect 55200 18504 56000 18624
rect 55200 18232 56000 18352
rect 0 17824 800 17944
rect 55200 17960 56000 18080
rect 55200 17688 56000 17808
rect 0 17280 800 17400
rect 55200 17416 56000 17536
rect 55200 17144 56000 17264
rect 0 16736 800 16856
rect 55200 16872 56000 16992
rect 55200 16600 56000 16720
rect 0 16192 800 16312
rect 55200 16328 56000 16448
rect 55200 16056 56000 16176
rect 0 15648 800 15768
rect 55200 15784 56000 15904
rect 55200 15512 56000 15632
rect 0 15104 800 15224
rect 55200 15240 56000 15360
rect 55200 14968 56000 15088
rect 0 14560 800 14680
rect 55200 14696 56000 14816
rect 55200 14424 56000 14544
rect 0 14016 800 14136
rect 55200 14152 56000 14272
rect 55200 13880 56000 14000
rect 0 13472 800 13592
rect 55200 13608 56000 13728
rect 55200 13336 56000 13456
rect 0 12928 800 13048
rect 55200 13064 56000 13184
rect 55200 12792 56000 12912
rect 0 12384 800 12504
rect 55200 12520 56000 12640
rect 55200 12248 56000 12368
rect 0 11840 800 11960
rect 55200 11976 56000 12096
rect 55200 11704 56000 11824
rect 0 11296 800 11416
rect 55200 11432 56000 11552
rect 55200 11160 56000 11280
rect 0 10752 800 10872
rect 55200 10888 56000 11008
rect 55200 10616 56000 10736
rect 0 10208 800 10328
rect 55200 10344 56000 10464
rect 55200 10072 56000 10192
rect 0 9664 800 9784
rect 55200 9800 56000 9920
rect 55200 9528 56000 9648
rect 0 9120 800 9240
rect 55200 9256 56000 9376
rect 55200 8984 56000 9104
rect 0 8576 800 8696
rect 55200 8712 56000 8832
rect 55200 8440 56000 8560
rect 0 8032 800 8152
rect 55200 8168 56000 8288
rect 55200 7896 56000 8016
rect 0 7488 800 7608
rect 55200 7624 56000 7744
rect 55200 7352 56000 7472
rect 0 6944 800 7064
rect 55200 7080 56000 7200
rect 55200 6808 56000 6928
rect 0 6400 800 6520
rect 55200 6536 56000 6656
rect 0 5856 800 5976
rect 0 5312 800 5432
rect 0 4768 800 4888
rect 0 4224 800 4344
rect 0 3680 800 3800
rect 0 3136 800 3256
<< obsm3 >>
rect 800 52840 55200 53345
rect 880 52560 55200 52840
rect 800 52296 55200 52560
rect 880 52016 55200 52296
rect 800 51752 55200 52016
rect 880 51472 55200 51752
rect 800 51208 55200 51472
rect 880 50928 55200 51208
rect 800 50664 55200 50928
rect 880 50384 55200 50664
rect 800 50120 55200 50384
rect 880 49840 55200 50120
rect 800 49576 55200 49840
rect 880 49440 55200 49576
rect 880 49296 55120 49440
rect 800 49032 55120 49296
rect 880 48752 55120 49032
rect 800 48488 55120 48752
rect 880 48208 55120 48488
rect 800 47944 55120 48208
rect 880 47664 55120 47944
rect 800 47400 55120 47664
rect 880 47120 55120 47400
rect 800 46856 55120 47120
rect 880 46576 55120 46856
rect 800 46312 55120 46576
rect 880 46032 55120 46312
rect 800 45768 55120 46032
rect 880 45488 55120 45768
rect 800 45224 55120 45488
rect 880 44944 55120 45224
rect 800 44680 55120 44944
rect 880 44400 55120 44680
rect 800 44136 55120 44400
rect 880 43856 55120 44136
rect 800 43592 55120 43856
rect 880 43312 55120 43592
rect 800 43048 55120 43312
rect 880 42768 55120 43048
rect 800 42504 55120 42768
rect 880 42224 55120 42504
rect 800 41960 55120 42224
rect 880 41680 55120 41960
rect 800 41416 55120 41680
rect 880 41136 55120 41416
rect 800 40872 55120 41136
rect 880 40592 55120 40872
rect 800 40328 55120 40592
rect 880 40048 55120 40328
rect 800 39784 55120 40048
rect 880 39504 55120 39784
rect 800 39240 55120 39504
rect 880 38960 55120 39240
rect 800 38696 55120 38960
rect 880 38416 55120 38696
rect 800 38152 55120 38416
rect 880 37872 55120 38152
rect 800 37608 55120 37872
rect 880 37328 55120 37608
rect 800 37064 55120 37328
rect 880 36784 55120 37064
rect 800 36520 55120 36784
rect 880 36240 55120 36520
rect 800 35976 55120 36240
rect 880 35696 55120 35976
rect 800 35432 55120 35696
rect 880 35152 55120 35432
rect 800 34888 55120 35152
rect 880 34608 55120 34888
rect 800 34344 55120 34608
rect 880 34064 55120 34344
rect 800 33800 55120 34064
rect 880 33520 55120 33800
rect 800 33256 55120 33520
rect 880 32976 55120 33256
rect 800 32712 55120 32976
rect 880 32432 55120 32712
rect 800 32168 55120 32432
rect 880 31888 55120 32168
rect 800 31624 55120 31888
rect 880 31344 55120 31624
rect 800 31080 55120 31344
rect 880 30800 55120 31080
rect 800 30536 55120 30800
rect 880 30256 55120 30536
rect 800 29992 55120 30256
rect 880 29712 55120 29992
rect 800 29448 55120 29712
rect 880 29168 55120 29448
rect 800 28904 55120 29168
rect 880 28624 55120 28904
rect 800 28360 55120 28624
rect 880 28080 55120 28360
rect 800 27816 55120 28080
rect 880 27536 55120 27816
rect 800 27272 55120 27536
rect 880 26992 55120 27272
rect 800 26728 55120 26992
rect 880 26448 55120 26728
rect 800 26184 55120 26448
rect 880 25904 55120 26184
rect 800 25640 55120 25904
rect 880 25360 55120 25640
rect 800 25096 55120 25360
rect 880 24816 55120 25096
rect 800 24552 55120 24816
rect 880 24272 55120 24552
rect 800 24008 55120 24272
rect 880 23728 55120 24008
rect 800 23464 55120 23728
rect 880 23184 55120 23464
rect 800 22920 55120 23184
rect 880 22640 55120 22920
rect 800 22376 55120 22640
rect 880 22096 55120 22376
rect 800 21832 55120 22096
rect 880 21552 55120 21832
rect 800 21288 55120 21552
rect 880 21008 55120 21288
rect 800 20744 55120 21008
rect 880 20464 55120 20744
rect 800 20200 55120 20464
rect 880 19920 55120 20200
rect 800 19656 55120 19920
rect 880 19376 55120 19656
rect 800 19112 55120 19376
rect 880 18832 55120 19112
rect 800 18568 55120 18832
rect 880 18288 55120 18568
rect 800 18024 55120 18288
rect 880 17744 55120 18024
rect 800 17480 55120 17744
rect 880 17200 55120 17480
rect 800 16936 55120 17200
rect 880 16656 55120 16936
rect 800 16392 55120 16656
rect 880 16112 55120 16392
rect 800 15848 55120 16112
rect 880 15568 55120 15848
rect 800 15304 55120 15568
rect 880 15024 55120 15304
rect 800 14760 55120 15024
rect 880 14480 55120 14760
rect 800 14216 55120 14480
rect 880 13936 55120 14216
rect 800 13672 55120 13936
rect 880 13392 55120 13672
rect 800 13128 55120 13392
rect 880 12848 55120 13128
rect 800 12584 55120 12848
rect 880 12304 55120 12584
rect 800 12040 55120 12304
rect 880 11760 55120 12040
rect 800 11496 55120 11760
rect 880 11216 55120 11496
rect 800 10952 55120 11216
rect 880 10672 55120 10952
rect 800 10408 55120 10672
rect 880 10128 55120 10408
rect 800 9864 55120 10128
rect 880 9584 55120 9864
rect 800 9320 55120 9584
rect 880 9040 55120 9320
rect 800 8776 55120 9040
rect 880 8496 55120 8776
rect 800 8232 55120 8496
rect 880 7952 55120 8232
rect 800 7688 55120 7952
rect 880 7408 55120 7688
rect 800 7144 55120 7408
rect 880 6864 55120 7144
rect 800 6600 55120 6864
rect 880 6456 55120 6600
rect 880 6320 55200 6456
rect 800 6056 55200 6320
rect 880 5776 55200 6056
rect 800 5512 55200 5776
rect 880 5232 55200 5512
rect 800 4968 55200 5232
rect 880 4688 55200 4968
rect 800 4424 55200 4688
rect 880 4144 55200 4424
rect 800 3880 55200 4144
rect 880 3600 55200 3880
rect 800 3336 55200 3600
rect 880 3056 55200 3336
rect 800 2143 55200 3056
<< metal4 >>
rect 4208 2128 4528 53360
rect 19568 2128 19888 53360
rect 34928 2128 35248 53360
rect 50288 2128 50608 53360
<< obsm4 >>
rect 25819 2347 34848 52597
rect 35328 2347 38397 52597
<< labels >>
rlabel metal3 s 0 17824 800 17944 6 design_clk_o
port 1 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 dsi_all[0]
port 2 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 dsi_all[10]
port 3 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 dsi_all[11]
port 4 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 dsi_all[12]
port 5 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 dsi_all[13]
port 6 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 dsi_all[14]
port 7 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 dsi_all[15]
port 8 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 dsi_all[16]
port 9 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 dsi_all[17]
port 10 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 dsi_all[18]
port 11 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 dsi_all[19]
port 12 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 dsi_all[1]
port 13 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 dsi_all[20]
port 14 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 dsi_all[21]
port 15 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 dsi_all[22]
port 16 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 dsi_all[23]
port 17 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 dsi_all[24]
port 18 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 dsi_all[25]
port 19 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 dsi_all[26]
port 20 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 dsi_all[2]
port 21 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 dsi_all[3]
port 22 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 dsi_all[4]
port 23 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 dsi_all[5]
port 24 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 dsi_all[6]
port 25 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 dsi_all[7]
port 26 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 dsi_all[8]
port 27 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 dsi_all[9]
port 28 nsew signal output
rlabel metal3 s 55200 34552 56000 34672 6 dso_6502[0]
port 29 nsew signal input
rlabel metal3 s 55200 37272 56000 37392 6 dso_6502[10]
port 30 nsew signal input
rlabel metal3 s 55200 37544 56000 37664 6 dso_6502[11]
port 31 nsew signal input
rlabel metal3 s 55200 37816 56000 37936 6 dso_6502[12]
port 32 nsew signal input
rlabel metal3 s 55200 38088 56000 38208 6 dso_6502[13]
port 33 nsew signal input
rlabel metal3 s 55200 38360 56000 38480 6 dso_6502[14]
port 34 nsew signal input
rlabel metal3 s 55200 38632 56000 38752 6 dso_6502[15]
port 35 nsew signal input
rlabel metal3 s 55200 38904 56000 39024 6 dso_6502[16]
port 36 nsew signal input
rlabel metal3 s 55200 39176 56000 39296 6 dso_6502[17]
port 37 nsew signal input
rlabel metal3 s 55200 39448 56000 39568 6 dso_6502[18]
port 38 nsew signal input
rlabel metal3 s 55200 39720 56000 39840 6 dso_6502[19]
port 39 nsew signal input
rlabel metal3 s 55200 34824 56000 34944 6 dso_6502[1]
port 40 nsew signal input
rlabel metal3 s 55200 39992 56000 40112 6 dso_6502[20]
port 41 nsew signal input
rlabel metal3 s 55200 40264 56000 40384 6 dso_6502[21]
port 42 nsew signal input
rlabel metal3 s 55200 40536 56000 40656 6 dso_6502[22]
port 43 nsew signal input
rlabel metal3 s 55200 40808 56000 40928 6 dso_6502[23]
port 44 nsew signal input
rlabel metal3 s 55200 41080 56000 41200 6 dso_6502[24]
port 45 nsew signal input
rlabel metal3 s 55200 41352 56000 41472 6 dso_6502[25]
port 46 nsew signal input
rlabel metal3 s 55200 41624 56000 41744 6 dso_6502[26]
port 47 nsew signal input
rlabel metal3 s 55200 35096 56000 35216 6 dso_6502[2]
port 48 nsew signal input
rlabel metal3 s 55200 35368 56000 35488 6 dso_6502[3]
port 49 nsew signal input
rlabel metal3 s 55200 35640 56000 35760 6 dso_6502[4]
port 50 nsew signal input
rlabel metal3 s 55200 35912 56000 36032 6 dso_6502[5]
port 51 nsew signal input
rlabel metal3 s 55200 36184 56000 36304 6 dso_6502[6]
port 52 nsew signal input
rlabel metal3 s 55200 36456 56000 36576 6 dso_6502[7]
port 53 nsew signal input
rlabel metal3 s 55200 36728 56000 36848 6 dso_6502[8]
port 54 nsew signal input
rlabel metal3 s 55200 37000 56000 37120 6 dso_6502[9]
port 55 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 dso_LCD[0]
port 56 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 dso_LCD[1]
port 57 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 dso_LCD[2]
port 58 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 dso_LCD[3]
port 59 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 dso_LCD[4]
port 60 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 dso_LCD[5]
port 61 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 dso_LCD[6]
port 62 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 dso_LCD[7]
port 63 nsew signal input
rlabel metal3 s 55200 41896 56000 42016 6 dso_as1802[0]
port 64 nsew signal input
rlabel metal3 s 55200 44616 56000 44736 6 dso_as1802[10]
port 65 nsew signal input
rlabel metal3 s 55200 44888 56000 45008 6 dso_as1802[11]
port 66 nsew signal input
rlabel metal3 s 55200 45160 56000 45280 6 dso_as1802[12]
port 67 nsew signal input
rlabel metal3 s 55200 45432 56000 45552 6 dso_as1802[13]
port 68 nsew signal input
rlabel metal3 s 55200 45704 56000 45824 6 dso_as1802[14]
port 69 nsew signal input
rlabel metal3 s 55200 45976 56000 46096 6 dso_as1802[15]
port 70 nsew signal input
rlabel metal3 s 55200 46248 56000 46368 6 dso_as1802[16]
port 71 nsew signal input
rlabel metal3 s 55200 46520 56000 46640 6 dso_as1802[17]
port 72 nsew signal input
rlabel metal3 s 55200 46792 56000 46912 6 dso_as1802[18]
port 73 nsew signal input
rlabel metal3 s 55200 47064 56000 47184 6 dso_as1802[19]
port 74 nsew signal input
rlabel metal3 s 55200 42168 56000 42288 6 dso_as1802[1]
port 75 nsew signal input
rlabel metal3 s 55200 47336 56000 47456 6 dso_as1802[20]
port 76 nsew signal input
rlabel metal3 s 55200 47608 56000 47728 6 dso_as1802[21]
port 77 nsew signal input
rlabel metal3 s 55200 47880 56000 48000 6 dso_as1802[22]
port 78 nsew signal input
rlabel metal3 s 55200 48152 56000 48272 6 dso_as1802[23]
port 79 nsew signal input
rlabel metal3 s 55200 48424 56000 48544 6 dso_as1802[24]
port 80 nsew signal input
rlabel metal3 s 55200 48696 56000 48816 6 dso_as1802[25]
port 81 nsew signal input
rlabel metal3 s 55200 48968 56000 49088 6 dso_as1802[26]
port 82 nsew signal input
rlabel metal3 s 55200 42440 56000 42560 6 dso_as1802[2]
port 83 nsew signal input
rlabel metal3 s 55200 42712 56000 42832 6 dso_as1802[3]
port 84 nsew signal input
rlabel metal3 s 55200 42984 56000 43104 6 dso_as1802[4]
port 85 nsew signal input
rlabel metal3 s 55200 43256 56000 43376 6 dso_as1802[5]
port 86 nsew signal input
rlabel metal3 s 55200 43528 56000 43648 6 dso_as1802[6]
port 87 nsew signal input
rlabel metal3 s 55200 43800 56000 43920 6 dso_as1802[7]
port 88 nsew signal input
rlabel metal3 s 55200 44072 56000 44192 6 dso_as1802[8]
port 89 nsew signal input
rlabel metal3 s 55200 44344 56000 44464 6 dso_as1802[9]
port 90 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 dso_as2650[0]
port 91 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 dso_as2650[10]
port 92 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 dso_as2650[11]
port 93 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 dso_as2650[12]
port 94 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 dso_as2650[13]
port 95 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 dso_as2650[14]
port 96 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 dso_as2650[15]
port 97 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 dso_as2650[16]
port 98 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 dso_as2650[17]
port 99 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 dso_as2650[18]
port 100 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 dso_as2650[19]
port 101 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 dso_as2650[1]
port 102 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 dso_as2650[20]
port 103 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 dso_as2650[21]
port 104 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 dso_as2650[22]
port 105 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 dso_as2650[23]
port 106 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 dso_as2650[24]
port 107 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 dso_as2650[25]
port 108 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 dso_as2650[26]
port 109 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 dso_as2650[2]
port 110 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 dso_as2650[3]
port 111 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 dso_as2650[4]
port 112 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 dso_as2650[5]
port 113 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 dso_as2650[6]
port 114 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 dso_as2650[7]
port 115 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 dso_as2650[8]
port 116 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 dso_as2650[9]
port 117 nsew signal input
rlabel metal2 s 11242 55200 11298 56000 6 dso_as5401[0]
port 118 nsew signal input
rlabel metal2 s 23202 55200 23258 56000 6 dso_as5401[10]
port 119 nsew signal input
rlabel metal2 s 24398 55200 24454 56000 6 dso_as5401[11]
port 120 nsew signal input
rlabel metal2 s 25594 55200 25650 56000 6 dso_as5401[12]
port 121 nsew signal input
rlabel metal2 s 26790 55200 26846 56000 6 dso_as5401[13]
port 122 nsew signal input
rlabel metal2 s 27986 55200 28042 56000 6 dso_as5401[14]
port 123 nsew signal input
rlabel metal2 s 29182 55200 29238 56000 6 dso_as5401[15]
port 124 nsew signal input
rlabel metal2 s 30378 55200 30434 56000 6 dso_as5401[16]
port 125 nsew signal input
rlabel metal2 s 31574 55200 31630 56000 6 dso_as5401[17]
port 126 nsew signal input
rlabel metal2 s 32770 55200 32826 56000 6 dso_as5401[18]
port 127 nsew signal input
rlabel metal2 s 33966 55200 34022 56000 6 dso_as5401[19]
port 128 nsew signal input
rlabel metal2 s 12438 55200 12494 56000 6 dso_as5401[1]
port 129 nsew signal input
rlabel metal2 s 35162 55200 35218 56000 6 dso_as5401[20]
port 130 nsew signal input
rlabel metal2 s 36358 55200 36414 56000 6 dso_as5401[21]
port 131 nsew signal input
rlabel metal2 s 37554 55200 37610 56000 6 dso_as5401[22]
port 132 nsew signal input
rlabel metal2 s 38750 55200 38806 56000 6 dso_as5401[23]
port 133 nsew signal input
rlabel metal2 s 39946 55200 40002 56000 6 dso_as5401[24]
port 134 nsew signal input
rlabel metal2 s 41142 55200 41198 56000 6 dso_as5401[25]
port 135 nsew signal input
rlabel metal2 s 42338 55200 42394 56000 6 dso_as5401[26]
port 136 nsew signal input
rlabel metal2 s 13634 55200 13690 56000 6 dso_as5401[2]
port 137 nsew signal input
rlabel metal2 s 14830 55200 14886 56000 6 dso_as5401[3]
port 138 nsew signal input
rlabel metal2 s 16026 55200 16082 56000 6 dso_as5401[4]
port 139 nsew signal input
rlabel metal2 s 17222 55200 17278 56000 6 dso_as5401[5]
port 140 nsew signal input
rlabel metal2 s 18418 55200 18474 56000 6 dso_as5401[6]
port 141 nsew signal input
rlabel metal2 s 19614 55200 19670 56000 6 dso_as5401[7]
port 142 nsew signal input
rlabel metal2 s 20810 55200 20866 56000 6 dso_as5401[8]
port 143 nsew signal input
rlabel metal2 s 22006 55200 22062 56000 6 dso_as5401[9]
port 144 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 dso_counter[0]
port 145 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dso_counter[10]
port 146 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 dso_counter[11]
port 147 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 dso_counter[1]
port 148 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 dso_counter[2]
port 149 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 dso_counter[3]
port 150 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 dso_counter[4]
port 151 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 dso_counter[5]
port 152 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 dso_counter[6]
port 153 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 dso_counter[7]
port 154 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 dso_counter[8]
port 155 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 dso_counter[9]
port 156 nsew signal input
rlabel metal2 s 44730 55200 44786 56000 6 dso_diceroll[0]
port 157 nsew signal input
rlabel metal2 s 45926 55200 45982 56000 6 dso_diceroll[1]
port 158 nsew signal input
rlabel metal2 s 47122 55200 47178 56000 6 dso_diceroll[2]
port 159 nsew signal input
rlabel metal2 s 48318 55200 48374 56000 6 dso_diceroll[3]
port 160 nsew signal input
rlabel metal2 s 49514 55200 49570 56000 6 dso_diceroll[4]
port 161 nsew signal input
rlabel metal2 s 50710 55200 50766 56000 6 dso_diceroll[5]
port 162 nsew signal input
rlabel metal2 s 51906 55200 51962 56000 6 dso_diceroll[6]
port 163 nsew signal input
rlabel metal2 s 53102 55200 53158 56000 6 dso_diceroll[7]
port 164 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 dso_mc14500[0]
port 165 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 dso_mc14500[1]
port 166 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 dso_mc14500[2]
port 167 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 dso_mc14500[3]
port 168 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 dso_mc14500[4]
port 169 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 dso_mc14500[5]
port 170 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 dso_mc14500[6]
port 171 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 dso_mc14500[7]
port 172 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 dso_mc14500[8]
port 173 nsew signal input
rlabel metal2 s 1674 55200 1730 56000 6 dso_multiplier[0]
port 174 nsew signal input
rlabel metal2 s 2870 55200 2926 56000 6 dso_multiplier[1]
port 175 nsew signal input
rlabel metal2 s 4066 55200 4122 56000 6 dso_multiplier[2]
port 176 nsew signal input
rlabel metal2 s 5262 55200 5318 56000 6 dso_multiplier[3]
port 177 nsew signal input
rlabel metal2 s 6458 55200 6514 56000 6 dso_multiplier[4]
port 178 nsew signal input
rlabel metal2 s 7654 55200 7710 56000 6 dso_multiplier[5]
port 179 nsew signal input
rlabel metal2 s 8850 55200 8906 56000 6 dso_multiplier[6]
port 180 nsew signal input
rlabel metal2 s 10046 55200 10102 56000 6 dso_multiplier[7]
port 181 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 dso_tbb1143[0]
port 182 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 dso_tbb1143[1]
port 183 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 dso_tbb1143[2]
port 184 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 dso_tbb1143[3]
port 185 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 dso_tbb1143[4]
port 186 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 dso_tbb1143[5]
port 187 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 dso_tbb1143[6]
port 188 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 dso_tbb1143[7]
port 189 nsew signal input
rlabel metal2 s 54298 55200 54354 56000 6 dso_tune
port 190 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 io_in[0]
port 191 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 io_in[10]
port 192 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_in[11]
port 193 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 io_in[12]
port 194 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 io_in[13]
port 195 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 io_in[14]
port 196 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 io_in[15]
port 197 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_in[16]
port 198 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 io_in[17]
port 199 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_in[18]
port 200 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 io_in[19]
port 201 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 io_in[1]
port 202 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 io_in[20]
port 203 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 io_in[21]
port 204 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 io_in[22]
port 205 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 io_in[23]
port 206 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 io_in[24]
port 207 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[25]
port 208 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 io_in[26]
port 209 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 io_in[27]
port 210 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 io_in[28]
port 211 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 io_in[29]
port 212 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 io_in[2]
port 213 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 io_in[30]
port 214 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 io_in[31]
port 215 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 216 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 io_in[33]
port 217 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 io_in[34]
port 218 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 io_in[35]
port 219 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 io_in[36]
port 220 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 io_in[37]
port 221 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 io_in[3]
port 222 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_in[4]
port 223 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 io_in[5]
port 224 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 io_in[6]
port 225 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 io_in[7]
port 226 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 io_in[8]
port 227 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 io_in[9]
port 228 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 io_oeb[0]
port 229 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 io_oeb[10]
port 230 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 io_oeb[11]
port 231 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[12]
port 232 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 io_oeb[13]
port 233 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 io_oeb[14]
port 234 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 io_oeb[15]
port 235 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 io_oeb[16]
port 236 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 io_oeb[17]
port 237 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 io_oeb[18]
port 238 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 io_oeb[19]
port 239 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 io_oeb[1]
port 240 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 io_oeb[20]
port 241 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 io_oeb[21]
port 242 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 io_oeb[22]
port 243 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 io_oeb[23]
port 244 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 io_oeb[24]
port 245 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 io_oeb[25]
port 246 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 io_oeb[26]
port 247 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 io_oeb[27]
port 248 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 io_oeb[28]
port 249 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 io_oeb[29]
port 250 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 io_oeb[2]
port 251 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 io_oeb[30]
port 252 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 io_oeb[31]
port 253 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 io_oeb[32]
port 254 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 io_oeb[33]
port 255 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 io_oeb[34]
port 256 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 io_oeb[35]
port 257 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 io_oeb[36]
port 258 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 io_oeb[37]
port 259 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[3]
port 260 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 io_oeb[4]
port 261 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_oeb[5]
port 262 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 io_oeb[6]
port 263 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 io_oeb[7]
port 264 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 io_oeb[8]
port 265 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 io_oeb[9]
port 266 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 io_out[0]
port 267 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 io_out[10]
port 268 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 io_out[11]
port 269 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 io_out[12]
port 270 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 io_out[13]
port 271 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_out[14]
port 272 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_out[15]
port 273 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 io_out[16]
port 274 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 io_out[17]
port 275 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 io_out[18]
port 276 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 io_out[19]
port 277 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_out[1]
port 278 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 io_out[20]
port 279 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 io_out[21]
port 280 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 io_out[22]
port 281 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_out[23]
port 282 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 io_out[24]
port 283 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 io_out[25]
port 284 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 io_out[26]
port 285 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 io_out[27]
port 286 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 io_out[28]
port 287 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_out[29]
port 288 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 io_out[2]
port 289 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 io_out[30]
port 290 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 io_out[31]
port 291 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_out[32]
port 292 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 io_out[33]
port 293 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 io_out[34]
port 294 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 io_out[35]
port 295 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 io_out[36]
port 296 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 io_out[37]
port 297 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 io_out[3]
port 298 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 io_out[4]
port 299 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_out[5]
port 300 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 io_out[6]
port 301 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 io_out[7]
port 302 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_out[8]
port 303 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 io_out[9]
port 304 nsew signal output
rlabel metal3 s 55200 34280 56000 34400 6 oeb_6502
port 305 nsew signal input
rlabel metal3 s 55200 49240 56000 49360 6 oeb_as1802
port 306 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 oeb_as2650
port 307 nsew signal input
rlabel metal2 s 43534 55200 43590 56000 6 oeb_as5401
port 308 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 oeb_mc14500
port 309 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 rst_6502
port 310 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 rst_LCD
port 311 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 rst_as1802
port 312 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 rst_as2650
port 313 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 rst_as5401
port 314 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 rst_counter
port 315 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 rst_diceroll
port 316 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 rst_mc14500
port 317 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 rst_tbb1143
port 318 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 rst_tune
port 319 nsew signal output
rlabel metal4 s 4208 2128 4528 53360 6 vccd1
port 320 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 53360 6 vccd1
port 320 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 53360 6 vssd1
port 321 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 53360 6 vssd1
port 321 nsew ground bidirectional
rlabel metal3 s 55200 6536 56000 6656 6 wb_clk_i
port 322 nsew signal input
rlabel metal3 s 55200 6808 56000 6928 6 wb_rst_i
port 323 nsew signal input
rlabel metal3 s 55200 7080 56000 7200 6 wbs_ack_o
port 324 nsew signal output
rlabel metal3 s 55200 8168 56000 8288 6 wbs_adr_i[0]
port 325 nsew signal input
rlabel metal3 s 55200 16328 56000 16448 6 wbs_adr_i[10]
port 326 nsew signal input
rlabel metal3 s 55200 17144 56000 17264 6 wbs_adr_i[11]
port 327 nsew signal input
rlabel metal3 s 55200 17960 56000 18080 6 wbs_adr_i[12]
port 328 nsew signal input
rlabel metal3 s 55200 18776 56000 18896 6 wbs_adr_i[13]
port 329 nsew signal input
rlabel metal3 s 55200 19592 56000 19712 6 wbs_adr_i[14]
port 330 nsew signal input
rlabel metal3 s 55200 20408 56000 20528 6 wbs_adr_i[15]
port 331 nsew signal input
rlabel metal3 s 55200 21224 56000 21344 6 wbs_adr_i[16]
port 332 nsew signal input
rlabel metal3 s 55200 22040 56000 22160 6 wbs_adr_i[17]
port 333 nsew signal input
rlabel metal3 s 55200 22856 56000 22976 6 wbs_adr_i[18]
port 334 nsew signal input
rlabel metal3 s 55200 23672 56000 23792 6 wbs_adr_i[19]
port 335 nsew signal input
rlabel metal3 s 55200 8984 56000 9104 6 wbs_adr_i[1]
port 336 nsew signal input
rlabel metal3 s 55200 24488 56000 24608 6 wbs_adr_i[20]
port 337 nsew signal input
rlabel metal3 s 55200 25304 56000 25424 6 wbs_adr_i[21]
port 338 nsew signal input
rlabel metal3 s 55200 26120 56000 26240 6 wbs_adr_i[22]
port 339 nsew signal input
rlabel metal3 s 55200 26936 56000 27056 6 wbs_adr_i[23]
port 340 nsew signal input
rlabel metal3 s 55200 27752 56000 27872 6 wbs_adr_i[24]
port 341 nsew signal input
rlabel metal3 s 55200 28568 56000 28688 6 wbs_adr_i[25]
port 342 nsew signal input
rlabel metal3 s 55200 29384 56000 29504 6 wbs_adr_i[26]
port 343 nsew signal input
rlabel metal3 s 55200 30200 56000 30320 6 wbs_adr_i[27]
port 344 nsew signal input
rlabel metal3 s 55200 31016 56000 31136 6 wbs_adr_i[28]
port 345 nsew signal input
rlabel metal3 s 55200 31832 56000 31952 6 wbs_adr_i[29]
port 346 nsew signal input
rlabel metal3 s 55200 9800 56000 9920 6 wbs_adr_i[2]
port 347 nsew signal input
rlabel metal3 s 55200 32648 56000 32768 6 wbs_adr_i[30]
port 348 nsew signal input
rlabel metal3 s 55200 33464 56000 33584 6 wbs_adr_i[31]
port 349 nsew signal input
rlabel metal3 s 55200 10616 56000 10736 6 wbs_adr_i[3]
port 350 nsew signal input
rlabel metal3 s 55200 11432 56000 11552 6 wbs_adr_i[4]
port 351 nsew signal input
rlabel metal3 s 55200 12248 56000 12368 6 wbs_adr_i[5]
port 352 nsew signal input
rlabel metal3 s 55200 13064 56000 13184 6 wbs_adr_i[6]
port 353 nsew signal input
rlabel metal3 s 55200 13880 56000 14000 6 wbs_adr_i[7]
port 354 nsew signal input
rlabel metal3 s 55200 14696 56000 14816 6 wbs_adr_i[8]
port 355 nsew signal input
rlabel metal3 s 55200 15512 56000 15632 6 wbs_adr_i[9]
port 356 nsew signal input
rlabel metal3 s 55200 7352 56000 7472 6 wbs_cyc_i
port 357 nsew signal input
rlabel metal3 s 55200 8440 56000 8560 6 wbs_dat_i[0]
port 358 nsew signal input
rlabel metal3 s 55200 16600 56000 16720 6 wbs_dat_i[10]
port 359 nsew signal input
rlabel metal3 s 55200 17416 56000 17536 6 wbs_dat_i[11]
port 360 nsew signal input
rlabel metal3 s 55200 18232 56000 18352 6 wbs_dat_i[12]
port 361 nsew signal input
rlabel metal3 s 55200 19048 56000 19168 6 wbs_dat_i[13]
port 362 nsew signal input
rlabel metal3 s 55200 19864 56000 19984 6 wbs_dat_i[14]
port 363 nsew signal input
rlabel metal3 s 55200 20680 56000 20800 6 wbs_dat_i[15]
port 364 nsew signal input
rlabel metal3 s 55200 21496 56000 21616 6 wbs_dat_i[16]
port 365 nsew signal input
rlabel metal3 s 55200 22312 56000 22432 6 wbs_dat_i[17]
port 366 nsew signal input
rlabel metal3 s 55200 23128 56000 23248 6 wbs_dat_i[18]
port 367 nsew signal input
rlabel metal3 s 55200 23944 56000 24064 6 wbs_dat_i[19]
port 368 nsew signal input
rlabel metal3 s 55200 9256 56000 9376 6 wbs_dat_i[1]
port 369 nsew signal input
rlabel metal3 s 55200 24760 56000 24880 6 wbs_dat_i[20]
port 370 nsew signal input
rlabel metal3 s 55200 25576 56000 25696 6 wbs_dat_i[21]
port 371 nsew signal input
rlabel metal3 s 55200 26392 56000 26512 6 wbs_dat_i[22]
port 372 nsew signal input
rlabel metal3 s 55200 27208 56000 27328 6 wbs_dat_i[23]
port 373 nsew signal input
rlabel metal3 s 55200 28024 56000 28144 6 wbs_dat_i[24]
port 374 nsew signal input
rlabel metal3 s 55200 28840 56000 28960 6 wbs_dat_i[25]
port 375 nsew signal input
rlabel metal3 s 55200 29656 56000 29776 6 wbs_dat_i[26]
port 376 nsew signal input
rlabel metal3 s 55200 30472 56000 30592 6 wbs_dat_i[27]
port 377 nsew signal input
rlabel metal3 s 55200 31288 56000 31408 6 wbs_dat_i[28]
port 378 nsew signal input
rlabel metal3 s 55200 32104 56000 32224 6 wbs_dat_i[29]
port 379 nsew signal input
rlabel metal3 s 55200 10072 56000 10192 6 wbs_dat_i[2]
port 380 nsew signal input
rlabel metal3 s 55200 32920 56000 33040 6 wbs_dat_i[30]
port 381 nsew signal input
rlabel metal3 s 55200 33736 56000 33856 6 wbs_dat_i[31]
port 382 nsew signal input
rlabel metal3 s 55200 10888 56000 11008 6 wbs_dat_i[3]
port 383 nsew signal input
rlabel metal3 s 55200 11704 56000 11824 6 wbs_dat_i[4]
port 384 nsew signal input
rlabel metal3 s 55200 12520 56000 12640 6 wbs_dat_i[5]
port 385 nsew signal input
rlabel metal3 s 55200 13336 56000 13456 6 wbs_dat_i[6]
port 386 nsew signal input
rlabel metal3 s 55200 14152 56000 14272 6 wbs_dat_i[7]
port 387 nsew signal input
rlabel metal3 s 55200 14968 56000 15088 6 wbs_dat_i[8]
port 388 nsew signal input
rlabel metal3 s 55200 15784 56000 15904 6 wbs_dat_i[9]
port 389 nsew signal input
rlabel metal3 s 55200 8712 56000 8832 6 wbs_dat_o[0]
port 390 nsew signal output
rlabel metal3 s 55200 16872 56000 16992 6 wbs_dat_o[10]
port 391 nsew signal output
rlabel metal3 s 55200 17688 56000 17808 6 wbs_dat_o[11]
port 392 nsew signal output
rlabel metal3 s 55200 18504 56000 18624 6 wbs_dat_o[12]
port 393 nsew signal output
rlabel metal3 s 55200 19320 56000 19440 6 wbs_dat_o[13]
port 394 nsew signal output
rlabel metal3 s 55200 20136 56000 20256 6 wbs_dat_o[14]
port 395 nsew signal output
rlabel metal3 s 55200 20952 56000 21072 6 wbs_dat_o[15]
port 396 nsew signal output
rlabel metal3 s 55200 21768 56000 21888 6 wbs_dat_o[16]
port 397 nsew signal output
rlabel metal3 s 55200 22584 56000 22704 6 wbs_dat_o[17]
port 398 nsew signal output
rlabel metal3 s 55200 23400 56000 23520 6 wbs_dat_o[18]
port 399 nsew signal output
rlabel metal3 s 55200 24216 56000 24336 6 wbs_dat_o[19]
port 400 nsew signal output
rlabel metal3 s 55200 9528 56000 9648 6 wbs_dat_o[1]
port 401 nsew signal output
rlabel metal3 s 55200 25032 56000 25152 6 wbs_dat_o[20]
port 402 nsew signal output
rlabel metal3 s 55200 25848 56000 25968 6 wbs_dat_o[21]
port 403 nsew signal output
rlabel metal3 s 55200 26664 56000 26784 6 wbs_dat_o[22]
port 404 nsew signal output
rlabel metal3 s 55200 27480 56000 27600 6 wbs_dat_o[23]
port 405 nsew signal output
rlabel metal3 s 55200 28296 56000 28416 6 wbs_dat_o[24]
port 406 nsew signal output
rlabel metal3 s 55200 29112 56000 29232 6 wbs_dat_o[25]
port 407 nsew signal output
rlabel metal3 s 55200 29928 56000 30048 6 wbs_dat_o[26]
port 408 nsew signal output
rlabel metal3 s 55200 30744 56000 30864 6 wbs_dat_o[27]
port 409 nsew signal output
rlabel metal3 s 55200 31560 56000 31680 6 wbs_dat_o[28]
port 410 nsew signal output
rlabel metal3 s 55200 32376 56000 32496 6 wbs_dat_o[29]
port 411 nsew signal output
rlabel metal3 s 55200 10344 56000 10464 6 wbs_dat_o[2]
port 412 nsew signal output
rlabel metal3 s 55200 33192 56000 33312 6 wbs_dat_o[30]
port 413 nsew signal output
rlabel metal3 s 55200 34008 56000 34128 6 wbs_dat_o[31]
port 414 nsew signal output
rlabel metal3 s 55200 11160 56000 11280 6 wbs_dat_o[3]
port 415 nsew signal output
rlabel metal3 s 55200 11976 56000 12096 6 wbs_dat_o[4]
port 416 nsew signal output
rlabel metal3 s 55200 12792 56000 12912 6 wbs_dat_o[5]
port 417 nsew signal output
rlabel metal3 s 55200 13608 56000 13728 6 wbs_dat_o[6]
port 418 nsew signal output
rlabel metal3 s 55200 14424 56000 14544 6 wbs_dat_o[7]
port 419 nsew signal output
rlabel metal3 s 55200 15240 56000 15360 6 wbs_dat_o[8]
port 420 nsew signal output
rlabel metal3 s 55200 16056 56000 16176 6 wbs_dat_o[9]
port 421 nsew signal output
rlabel metal3 s 55200 7624 56000 7744 6 wbs_stb_i
port 422 nsew signal input
rlabel metal3 s 55200 7896 56000 8016 6 wbs_we_i
port 423 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 56000 56000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4654602
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Multiplexer/runs/23_02_13_17_50/results/signoff/multiplexer.magic.gds
string GDS_START 417362
<< end >>

