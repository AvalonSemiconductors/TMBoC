VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tune_player
  CLASS BLOCK ;
  FOREIGN tune_player ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN OP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END OP
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.080 10.640 18.680 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.805 10.640 43.405 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.530 10.640 68.130 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.255 10.640 92.855 98.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.440 10.640 31.040 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.165 10.640 55.765 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.890 10.640 80.490 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.615 10.640 105.215 98.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 4.670 10.640 105.215 98.160 ;
      LAYER met2 ;
        RECT 4.690 10.695 105.185 98.105 ;
      LAYER met3 ;
        RECT 4.000 92.160 105.205 98.085 ;
        RECT 4.400 90.760 105.205 92.160 ;
        RECT 4.000 55.440 105.205 90.760 ;
        RECT 4.400 54.040 105.205 55.440 ;
        RECT 4.000 18.720 105.205 54.040 ;
        RECT 4.400 17.320 105.205 18.720 ;
        RECT 4.000 10.715 105.205 17.320 ;
  END
END tune_player
END LIBRARY

