magic
tech sky130B
magscale 1 2
timestamp 1680008814
<< nwell >>
rect 1066 28549 30858 29115
rect 1066 27461 30858 28027
rect 1066 26373 30858 26939
rect 1066 25285 30858 25851
rect 1066 24197 30858 24763
rect 1066 23109 30858 23675
rect 1066 22021 30858 22587
rect 1066 20933 30858 21499
rect 1066 19845 30858 20411
rect 1066 18757 30858 19323
rect 1066 17669 30858 18235
rect 1066 16581 30858 17147
rect 1066 15493 30858 16059
rect 1066 14405 30858 14971
rect 1066 13317 30858 13883
rect 1066 12229 30858 12795
rect 1066 11141 30858 11707
rect 1066 10053 30858 10619
rect 1066 8965 30858 9531
rect 1066 7877 30858 8443
rect 1066 6789 30858 7355
rect 1066 5701 30858 6267
rect 1066 4613 30858 5179
rect 1066 3525 30858 4091
rect 1066 2437 30858 3003
<< obsli1 >>
rect 1104 2159 30820 29393
<< obsm1 >>
rect 1104 2128 31082 29424
<< metal2 >>
rect 2134 31200 2190 32000
rect 6090 31200 6146 32000
rect 10046 31200 10102 32000
rect 14002 31200 14058 32000
rect 17958 31200 18014 32000
rect 21914 31200 21970 32000
rect 25870 31200 25926 32000
rect 29826 31200 29882 32000
<< obsm2 >>
rect 1860 31144 2078 31362
rect 2246 31144 6034 31362
rect 6202 31144 9990 31362
rect 10158 31144 13946 31362
rect 14114 31144 17902 31362
rect 18070 31144 21858 31362
rect 22026 31144 25814 31362
rect 25982 31144 29770 31362
rect 29938 31144 31078 31362
rect 1860 1935 31078 31144
<< metal3 >>
rect 31200 29656 32000 29776
rect 31200 25712 32000 25832
rect 31200 21768 32000 21888
rect 31200 17824 32000 17944
rect 31200 13880 32000 14000
rect 31200 9936 32000 10056
rect 31200 5992 32000 6112
rect 31200 2048 32000 2168
<< obsm3 >>
rect 4660 29576 31120 29749
rect 4660 25912 31218 29576
rect 4660 25632 31120 25912
rect 4660 21968 31218 25632
rect 4660 21688 31120 21968
rect 4660 18024 31218 21688
rect 4660 17744 31120 18024
rect 4660 14080 31218 17744
rect 4660 13800 31120 14080
rect 4660 10136 31218 13800
rect 4660 9856 31120 10136
rect 4660 6192 31218 9856
rect 4660 5912 31120 6192
rect 4660 2248 31218 5912
rect 4660 1968 31120 2248
rect 4660 1939 31218 1968
<< metal4 >>
rect 4658 2128 4978 29424
rect 8372 2128 8692 29424
rect 12086 2128 12406 29424
rect 15800 2128 16120 29424
rect 19514 2128 19834 29424
rect 23228 2128 23548 29424
rect 26942 2128 27262 29424
rect 30656 2128 30976 29424
<< labels >>
rlabel metal2 s 2134 31200 2190 32000 6 clk
port 1 nsew signal input
rlabel metal2 s 10046 31200 10102 32000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 14002 31200 14058 32000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 17958 31200 18014 32000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 21914 31200 21970 32000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 25870 31200 25926 32000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 29826 31200 29882 32000 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 31200 2048 32000 2168 6 io_out[0]
port 8 nsew signal output
rlabel metal3 s 31200 5992 32000 6112 6 io_out[1]
port 9 nsew signal output
rlabel metal3 s 31200 9936 32000 10056 6 io_out[2]
port 10 nsew signal output
rlabel metal3 s 31200 13880 32000 14000 6 io_out[3]
port 11 nsew signal output
rlabel metal3 s 31200 17824 32000 17944 6 io_out[4]
port 12 nsew signal output
rlabel metal3 s 31200 21768 32000 21888 6 io_out[5]
port 13 nsew signal output
rlabel metal3 s 31200 25712 32000 25832 6 io_out[6]
port 14 nsew signal output
rlabel metal3 s 31200 29656 32000 29776 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 6090 31200 6146 32000 6 rst
port 16 nsew signal input
rlabel metal4 s 4658 2128 4978 29424 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 12086 2128 12406 29424 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 19514 2128 19834 29424 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 26942 2128 27262 29424 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 8372 2128 8692 29424 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 15800 2128 16120 29424 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 23228 2128 23548 29424 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 30656 2128 30976 29424 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32000 32000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1829308
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/TBB1143/runs/23_03_28_15_05/results/signoff/tholin_avalonsemi_tbb1143.magic.gds
string GDS_START 460618
<< end >>

