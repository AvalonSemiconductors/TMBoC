VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt2_tholin_namebadge
  CLASS BLOCK ;
  FOREIGN tt2_tholin_namebadge ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 125.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 121.000 12.790 125.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 121.000 62.470 125.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 121.000 87.310 125.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 121.000 112.150 125.000 ;
    END
  END io_in[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END io_out[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 121.000 37.630 125.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.920 10.640 20.520 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.325 10.640 48.925 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.730 10.640 77.330 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.135 10.640 105.735 111.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 33.120 10.640 34.720 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.525 10.640 63.125 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.930 10.640 91.530 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.335 10.640 119.935 111.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 110.105 119.330 111.710 ;
        RECT 5.330 104.665 119.330 107.495 ;
        RECT 5.330 99.225 119.330 102.055 ;
        RECT 5.330 93.785 119.330 96.615 ;
        RECT 5.330 88.345 119.330 91.175 ;
        RECT 5.330 82.905 119.330 85.735 ;
        RECT 5.330 77.465 119.330 80.295 ;
        RECT 5.330 72.025 119.330 74.855 ;
        RECT 5.330 66.585 119.330 69.415 ;
        RECT 5.330 61.145 119.330 63.975 ;
        RECT 5.330 55.705 119.330 58.535 ;
        RECT 5.330 50.265 119.330 53.095 ;
        RECT 5.330 44.825 119.330 47.655 ;
        RECT 5.330 39.385 119.330 42.215 ;
        RECT 5.330 33.945 119.330 36.775 ;
        RECT 5.330 28.505 119.330 31.335 ;
        RECT 5.330 23.065 119.330 25.895 ;
        RECT 5.330 17.625 119.330 20.455 ;
        RECT 5.330 12.185 119.330 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 119.140 111.605 ;
      LAYER met1 ;
        RECT 5.520 4.460 119.935 111.760 ;
      LAYER met2 ;
        RECT 7.450 120.720 12.230 121.000 ;
        RECT 13.070 120.720 37.070 121.000 ;
        RECT 37.910 120.720 61.910 121.000 ;
        RECT 62.750 120.720 86.750 121.000 ;
        RECT 87.590 120.720 111.590 121.000 ;
        RECT 112.430 120.720 119.905 121.000 ;
        RECT 7.450 4.280 119.905 120.720 ;
        RECT 8.010 3.670 10.390 4.280 ;
        RECT 11.230 3.670 13.610 4.280 ;
        RECT 14.450 3.670 16.830 4.280 ;
        RECT 17.670 3.670 20.050 4.280 ;
        RECT 20.890 3.670 23.270 4.280 ;
        RECT 24.110 3.670 26.490 4.280 ;
        RECT 27.330 3.670 29.710 4.280 ;
        RECT 30.550 3.670 32.930 4.280 ;
        RECT 33.770 3.670 36.150 4.280 ;
        RECT 36.990 3.670 39.370 4.280 ;
        RECT 40.210 3.670 42.590 4.280 ;
        RECT 43.430 3.670 45.810 4.280 ;
        RECT 46.650 3.670 49.030 4.280 ;
        RECT 49.870 3.670 52.250 4.280 ;
        RECT 53.090 3.670 55.470 4.280 ;
        RECT 56.310 3.670 58.690 4.280 ;
        RECT 59.530 3.670 61.910 4.280 ;
        RECT 62.750 3.670 65.130 4.280 ;
        RECT 65.970 3.670 68.350 4.280 ;
        RECT 69.190 3.670 71.570 4.280 ;
        RECT 72.410 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.010 4.280 ;
        RECT 78.850 3.670 81.230 4.280 ;
        RECT 82.070 3.670 84.450 4.280 ;
        RECT 85.290 3.670 87.670 4.280 ;
        RECT 88.510 3.670 90.890 4.280 ;
        RECT 91.730 3.670 94.110 4.280 ;
        RECT 94.950 3.670 97.330 4.280 ;
        RECT 98.170 3.670 100.550 4.280 ;
        RECT 101.390 3.670 103.770 4.280 ;
        RECT 104.610 3.670 106.990 4.280 ;
        RECT 107.830 3.670 110.210 4.280 ;
        RECT 111.050 3.670 113.430 4.280 ;
        RECT 114.270 3.670 116.650 4.280 ;
        RECT 117.490 3.670 119.905 4.280 ;
      LAYER met3 ;
        RECT 7.425 10.715 119.925 111.685 ;
      LAYER met4 ;
        RECT 21.455 12.415 32.720 106.585 ;
        RECT 35.120 12.415 46.925 106.585 ;
        RECT 49.325 12.415 61.125 106.585 ;
        RECT 63.525 12.415 75.330 106.585 ;
        RECT 77.730 12.415 89.530 106.585 ;
        RECT 91.930 12.415 99.985 106.585 ;
  END
END tt2_tholin_namebadge
END LIBRARY

