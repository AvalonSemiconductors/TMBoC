magic
tech sky130B
magscale 1 2
timestamp 1680261785
<< nwell >>
rect 1066 27461 28926 27782
rect 1066 26373 28926 26939
rect 1066 25285 28926 25851
rect 1066 24197 28926 24763
rect 1066 23109 28926 23675
rect 1066 22021 28926 22587
rect 1066 20933 28926 21499
rect 1066 19845 28926 20411
rect 1066 18757 28926 19323
rect 1066 17669 28926 18235
rect 1066 16581 28926 17147
rect 1066 15493 28926 16059
rect 1066 14405 28926 14971
rect 1066 13317 28926 13883
rect 1066 12229 28926 12795
rect 1066 11141 28926 11707
rect 1066 10053 28926 10619
rect 1066 8965 28926 9531
rect 1066 7877 28926 8443
rect 1066 6789 28926 7355
rect 1066 5701 28926 6267
rect 1066 4613 28926 5179
rect 1066 3525 28926 4091
rect 1066 2437 28926 3003
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 1104 2128 29048 27792
<< metal2 >>
rect 2042 29200 2098 30000
rect 5722 29200 5778 30000
rect 9402 29200 9458 30000
rect 13082 29200 13138 30000
rect 16762 29200 16818 30000
rect 20442 29200 20498 30000
rect 24122 29200 24178 30000
rect 27802 29200 27858 30000
<< obsm2 >>
rect 1584 29144 1986 29322
rect 2154 29144 5666 29322
rect 5834 29144 9346 29322
rect 9514 29144 13026 29322
rect 13194 29144 16706 29322
rect 16874 29144 20386 29322
rect 20554 29144 24066 29322
rect 24234 29144 27746 29322
rect 27914 29144 29042 29322
rect 1584 2139 29042 29144
<< metal3 >>
rect 29200 27752 30000 27872
rect 29200 24080 30000 24200
rect 29200 20408 30000 20528
rect 29200 16736 30000 16856
rect 29200 13064 30000 13184
rect 29200 9392 30000 9512
rect 29200 5720 30000 5840
rect 29200 2048 30000 2168
<< obsm3 >>
rect 4419 27672 29120 27845
rect 4419 24280 29378 27672
rect 4419 24000 29120 24280
rect 4419 20608 29378 24000
rect 4419 20328 29120 20608
rect 4419 16936 29378 20328
rect 4419 16656 29120 16936
rect 4419 13264 29378 16656
rect 4419 12984 29120 13264
rect 4419 9592 29378 12984
rect 4419 9312 29120 9592
rect 4419 5920 29378 9312
rect 4419 5640 29120 5920
rect 4419 2248 29378 5640
rect 4419 2143 29120 2248
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< labels >>
rlabel metal2 s 2042 29200 2098 30000 6 clk
port 1 nsew signal input
rlabel metal2 s 9402 29200 9458 30000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 13082 29200 13138 30000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 16762 29200 16818 30000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 20442 29200 20498 30000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 24122 29200 24178 30000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 27802 29200 27858 30000 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 29200 2048 30000 2168 6 io_out[0]
port 8 nsew signal output
rlabel metal3 s 29200 5720 30000 5840 6 io_out[1]
port 9 nsew signal output
rlabel metal3 s 29200 9392 30000 9512 6 io_out[2]
port 10 nsew signal output
rlabel metal3 s 29200 13064 30000 13184 6 io_out[3]
port 11 nsew signal output
rlabel metal3 s 29200 16736 30000 16856 6 io_out[4]
port 12 nsew signal output
rlabel metal3 s 29200 20408 30000 20528 6 io_out[5]
port 13 nsew signal output
rlabel metal3 s 29200 24080 30000 24200 6 io_out[6]
port 14 nsew signal output
rlabel metal3 s 29200 27752 30000 27872 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 5722 29200 5778 30000 6 rst
port 16 nsew signal input
rlabel metal4 s 4417 2128 4737 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1880304
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/TBB1143/runs/23_03_31_13_18/results/signoff/tholin_avalonsemi_tbb1143.magic.gds
string GDS_START 469992
<< end >>

