// This is the unpowered netlist.
module wrapped_as2650 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [7:0] io_in;
 output [26:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.sense ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \lfsr[0] ;
 wire \lfsr[10] ;
 wire \lfsr[11] ;
 wire \lfsr[12] ;
 wire \lfsr[13] ;
 wire \lfsr[14] ;
 wire \lfsr[15] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \lfsr[8] ;
 wire \lfsr[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__A (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__B (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__C (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A3 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__B (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__C_N (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__B (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__S (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__B (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__B (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__A_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__C (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__C (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__C (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__C (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A (.DIODE(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A (.DIODE(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A (.DIODE(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__B (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__C (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__B (.DIODE(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__B (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__C (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__C (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__D (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__C (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__D (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A2 (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A3 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B2 (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__D (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__B (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__B (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__B (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A_N (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A_N (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__C (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__B (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__C (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A2 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__S1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__B (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__B (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__B (.DIODE(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__C_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__B (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__B (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__B1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A_N (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__B (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__B1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__S1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__B (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A2 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A2 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A_N (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__B (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A_N (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__B (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A2 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A (.DIODE(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__B (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A (.DIODE(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__B (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A2 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__B (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__B (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A2 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A3 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B1 (.DIODE(_2925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__B (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__C1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__D1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__C1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__B2 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__S (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A1 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A2 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__B (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A0 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A1 (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__S (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A0 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__B1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(_2874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A2 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A1 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A2 (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__B1 (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__B1 (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A2 (.DIODE(_2986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A2 (.DIODE(_2987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__B2 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A2 (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B2 (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__C (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__C (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B1 (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__B2 (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A2 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A2 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A1 (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__C1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A1 (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A1 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B (.DIODE(_0334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A1 (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B1 (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A0 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__S1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__C (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B2 (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B1 (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__S (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__C1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A1 (.DIODE(_2925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__C1 (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A0 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A2 (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B1 (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__S1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B2 (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__D (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A2 (.DIODE(_2958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A2 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A2 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B1 (.DIODE(_2925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B1 (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__B2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__C1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A2 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A2 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A2 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__C1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__C (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__S (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B1 (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__S0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A2 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A2 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A1 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A0 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__C1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A1 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A2 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__C1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B2 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A1 (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B2 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__C (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A (.DIODE(_2945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A2 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A2 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B2 (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A2 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__S (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__C1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A1 (.DIODE(_2925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__C1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A2 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A1 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A2 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A1 (.DIODE(_2909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B1 (.DIODE(_2930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__B2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__B1 (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A2 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A3 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A1 (.DIODE(_2915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A2 (.DIODE(_0552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A2 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__C (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__C (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__C (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A0 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__S (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__S (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__C (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A0 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__S (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B1 (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A0 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B1 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A1 (.DIODE(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A1 (.DIODE(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B2 (.DIODE(\as2650.pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A1 (.DIODE(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B2 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B2 (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__C (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__C (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A1 (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A2 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A (.DIODE(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A1 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A1 (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A2 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__C (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A0 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A1 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(_2986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B1 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A0 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A1 (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A1 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B1 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A1 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A2 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A0 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__B (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A1 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A1 (.DIODE(_0552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A1 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A0 (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__C (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__C (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__C (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A3 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__C_N (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__D1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__C1 (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__D1 (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__S (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__C (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__C (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__B (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__S (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__S (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B (.DIODE(_2986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__C (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__D (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A1 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A2 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B1 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__C (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__D (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A3 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__C1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__D (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(_2804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__C_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__D_N (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__C (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A3 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__C (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__B (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__B (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__C (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B (.DIODE(_2767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__C (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__C (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__B (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__S (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__C1 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__C (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__D (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B1 (.DIODE(_0543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__C1 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__C (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__D (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A1 (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A2 (.DIODE(_2651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B2 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__B1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B1 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A (.DIODE(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__B2 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A1 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A1 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(\as2650.psu[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A2 (.DIODE(_2651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(\as2650.psu[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A2 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B2 (.DIODE(\as2650.psu[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__B1 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B1 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B2 (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A3 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A2 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__S (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__C1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__S (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B2 (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__S (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A0 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A2 (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__C (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__D_N (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A2 (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A2 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__C (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A1_N (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A1_N (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__C (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__D (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__C (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__D (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A1_N (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__D (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__B2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A1_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A1_N (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A1 (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B1 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__C1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__D (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__B2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__C (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A1_N (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A2 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A2 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A2 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__B (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__C (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A0 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A1 (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(\as2650.sense ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A1 (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A2 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A2 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A2 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A2 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__C (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B1 (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__C (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B1 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B1_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__C1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__D (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A2 (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A1 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__D (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__B1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A2 (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__D1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A_N (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__C (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__B1 (.DIODE(_2651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A1 (.DIODE(_2651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A2 (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A3 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__C (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A2 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B2 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A2 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__B (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B2 (.DIODE(_2651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__B1 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__B2 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__C1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__B (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__B (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A2 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1_N (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A2_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__B (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B1 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__B (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__C (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__B1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__B2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B2 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A2 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B2 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__B (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__B (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A2 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B1 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1_N (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B2 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B2 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B2 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1_N (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A1 (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A2 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__B (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A0 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__B (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1_N (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A1 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A2 (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__B1 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A1_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A2 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A2 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A2 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__B (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A0 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A0 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A2 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B2 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__C1 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__D1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A1_N (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A2_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__B (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__B (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__C1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__B (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B1 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__C1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B (.DIODE(_0552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B (.DIODE(_0552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B1 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B1 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__B1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A2 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__C1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B1 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B1 (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B2 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__B2 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__C1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__B2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__C1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__B1 (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A2 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__B1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A1_N (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B2 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B2 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__C1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B1 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A2 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__C1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__C1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A2 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A2 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__C1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__C1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__S (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A2 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A1_N (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A1_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A2_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A4 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__C1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__S (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A2 (.DIODE(_2744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__C (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A3 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B1 (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A2 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A2_N (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A2 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A2 (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A3 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A2 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A3 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__C (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B1 (.DIODE(_1397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A3 (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__C (.DIODE(_2727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A2 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__C1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A2 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__C1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A3 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A0 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A (.DIODE(\as2650.r0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__C1 (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__C (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A (.DIODE(_2937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A2_N (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A2 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A2 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__B2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2_N (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__C (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__C (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A3 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A_N (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__C (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A2 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__D1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A1 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A2 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__D1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A3 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__B1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A1 (.DIODE(_2737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A3 (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A3 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__C1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__C1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__C1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__S (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B2 (.DIODE(\as2650.sense ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__C1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A1 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__C1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__S (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A (.DIODE(_2635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__C (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__C1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__C (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__C (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(_2728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__C1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__C (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A3 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A2 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(_2001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B1 (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__B (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A0 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__S (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B2 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A2 (.DIODE(_2018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B1 (.DIODE(_2852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B1 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__C1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(\as2650.pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A0 (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__C1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B2 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B (.DIODE(_0303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__C1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B1 (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B2 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A0 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__S (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(_1397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B1 (.DIODE(_2075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B2 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__C1 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(_2096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B2 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__C1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__C1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A1 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B1 (.DIODE(_2124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A0 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__S (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A1 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A2 (.DIODE(_2132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__C1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A2 (.DIODE(_2132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B2 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B2 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__C1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A0 (.DIODE(\as2650.addr_buff[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__S (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1_N (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A2 (.DIODE(_2168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__C1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B1_N (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B (.DIODE(_2168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__S (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1_N (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A2_N (.DIODE(_2183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__C1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A0 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B1 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A2 (.DIODE(_2194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B (.DIODE(_2208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B2 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B1 (.DIODE(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A_N (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__C_N (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B (.DIODE(_2208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__C1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A2 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__C1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B2 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1_N (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A2_N (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B2 (.DIODE(_2993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__B1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__S (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A (.DIODE(\as2650.pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A2_N (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__D1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_0340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A0 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A1 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__C1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A1 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B1 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__C1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A3 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A3 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(\as2650.pc[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__C1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A (.DIODE(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__B (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__C (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__C1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__C1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(\as2650.pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A2 (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__C1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A0 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(_2912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B1 (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B1 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A3 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__B1 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(\as2650.psu[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A2 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A2 (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__C1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__C1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A3 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A3 (.DIODE(_2865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__D1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__C1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B (.DIODE(_2986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A0 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A2 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A2 (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(_2001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__C1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A2 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__C1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__B1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A0 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A2 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A2 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__B1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A2 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__C1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A2 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__C1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__C1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B1 (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A0 (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A1 (.DIODE(\as2650.psu[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A2 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B1 (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__C1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A2 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A0 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A2 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A (.DIODE(\as2650.psu[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A1 (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__C1 (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A2 (.DIODE(_2096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B1 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A2 (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__C1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A2 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__B (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A0 (.DIODE(_2124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A0 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A2 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B1 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__C1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A0 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__B1 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A2 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__C1 (.DIODE(_2792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__B2 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A0 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_0552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B (.DIODE(_2183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B2 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A2 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B2 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__C1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A2 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__C (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A0 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__C (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A1 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A1 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__S (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A3 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B2 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(_2987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(_0334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A1 (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A1 (.DIODE(_2935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1 (.DIODE(_2987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(_0334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A2 (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A0 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A1 (.DIODE(_2629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A2 (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A0 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(_2507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A1 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__C1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B1 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(_0399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__C1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B1 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__C1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__B1 (.DIODE(_2515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__C1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A0 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A1 (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A2 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__C_N (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__C (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A2 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__C1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__C1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__B1 (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B1 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A2 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__B (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A1 (.DIODE(_2986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__B1_N (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A2 (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2_N (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B1 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A1 (.DIODE(\as2650.carry ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__B2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A3 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A2 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B1 (.DIODE(_2567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__S (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__B1 (.DIODE(_2567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__S (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A2 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__B1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B1 (.DIODE(_2567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__C (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__C1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A3 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A0 (.DIODE(\as2650.psu[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A2 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__B1 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A2 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__B1 (.DIODE(\as2650.psl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A3 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__C1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B1 (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1_N (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__C1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__B1 (.DIODE(\as2650.psu[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B1 (.DIODE(\as2650.psu[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__CLK (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__CLK (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(_2852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(_2852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(\as2650.psu[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(\as2650.psu[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(\as2650.r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(\as2650.r0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(\as2650.r0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(\as2650.pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(\as2650.pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(\as2650.pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(\as2650.pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(\as2650.addr_buff[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_1397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkinv_2 _3001_ (.A(\as2650.psl[1] ),
    .Y(_2623_));
 sky130_fd_sc_hd__clkinv_4 _3002_ (.A(net223),
    .Y(_2624_));
 sky130_fd_sc_hd__inv_2 _3003_ (.A(\as2650.overflow ),
    .Y(_2625_));
 sky130_fd_sc_hd__inv_2 _3004_ (.A(net224),
    .Y(_2626_));
 sky130_fd_sc_hd__clkinv_4 _3005_ (.A(net228),
    .Y(_2627_));
 sky130_fd_sc_hd__inv_2 _3006_ (.A(net241),
    .Y(_2628_));
 sky130_fd_sc_hd__inv_2 _3007_ (.A(net267),
    .Y(_2629_));
 sky130_fd_sc_hd__inv_2 _3008_ (.A(net271),
    .Y(_2630_));
 sky130_fd_sc_hd__inv_2 _3009_ (.A(net274),
    .Y(_2631_));
 sky130_fd_sc_hd__clkinv_4 _3010_ (.A(net281),
    .Y(_2632_));
 sky130_fd_sc_hd__inv_4 _3011_ (.A(net283),
    .Y(_2633_));
 sky130_fd_sc_hd__inv_4 _3012_ (.A(\as2650.pc[2] ),
    .Y(_2634_));
 sky130_fd_sc_hd__clkinv_4 _3013_ (.A(net286),
    .Y(_2635_));
 sky130_fd_sc_hd__inv_4 _3014_ (.A(net295),
    .Y(_2636_));
 sky130_fd_sc_hd__inv_6 _3015_ (.A(\as2650.cycle[7] ),
    .Y(_2637_));
 sky130_fd_sc_hd__inv_2 _3016_ (.A(net293),
    .Y(_2638_));
 sky130_fd_sc_hd__inv_2 _3017_ (.A(\as2650.idx_ctrl[1] ),
    .Y(_2639_));
 sky130_fd_sc_hd__clkinv_4 _3018_ (.A(\as2650.idx_ctrl[0] ),
    .Y(_2640_));
 sky130_fd_sc_hd__clkinv_2 _3019_ (.A(net24),
    .Y(net10));
 sky130_fd_sc_hd__inv_2 _3020_ (.A(\as2650.psl[7] ),
    .Y(_2641_));
 sky130_fd_sc_hd__inv_2 _3021_ (.A(\as2650.psl[6] ),
    .Y(_2642_));
 sky130_fd_sc_hd__inv_2 _3022_ (.A(net306),
    .Y(_2643_));
 sky130_fd_sc_hd__inv_2 _3023_ (.A(net304),
    .Y(_2644_));
 sky130_fd_sc_hd__inv_2 _3024_ (.A(net237),
    .Y(_2645_));
 sky130_fd_sc_hd__inv_4 _3025_ (.A(net230),
    .Y(_2646_));
 sky130_fd_sc_hd__inv_8 _3026_ (.A(net299),
    .Y(_2647_));
 sky130_fd_sc_hd__inv_4 _3027_ (.A(net309),
    .Y(_2648_));
 sky130_fd_sc_hd__inv_4 _3028_ (.A(net324),
    .Y(_2649_));
 sky130_fd_sc_hd__clkinv_4 _3029_ (.A(net326),
    .Y(_2650_));
 sky130_fd_sc_hd__clkinv_4 _3030_ (.A(net349),
    .Y(_2651_));
 sky130_fd_sc_hd__inv_4 _3031_ (.A(net346),
    .Y(_2652_));
 sky130_fd_sc_hd__clkinv_2 _3032_ (.A(net342),
    .Y(_2653_));
 sky130_fd_sc_hd__inv_8 _3033_ (.A(net341),
    .Y(_2654_));
 sky130_fd_sc_hd__inv_6 _3034_ (.A(net339),
    .Y(_2655_));
 sky130_fd_sc_hd__inv_2 _3035_ (.A(\as2650.holding_reg[4] ),
    .Y(_2656_));
 sky130_fd_sc_hd__inv_2 _3036_ (.A(net336),
    .Y(_2657_));
 sky130_fd_sc_hd__clkinv_4 _3037_ (.A(net334),
    .Y(_2658_));
 sky130_fd_sc_hd__inv_2 _3038_ (.A(\as2650.holding_reg[7] ),
    .Y(_2659_));
 sky130_fd_sc_hd__inv_2 _3039_ (.A(net310),
    .Y(_2660_));
 sky130_fd_sc_hd__inv_2 _3040_ (.A(\as2650.addr_buff[1] ),
    .Y(_2661_));
 sky130_fd_sc_hd__inv_2 _3041_ (.A(\as2650.addr_buff[4] ),
    .Y(_2662_));
 sky130_fd_sc_hd__inv_2 _3042_ (.A(\lfsr[0] ),
    .Y(_2663_));
 sky130_fd_sc_hd__nor2_4 _3043_ (.A(net216),
    .B(net213),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(net235),
    .B(net230),
    .Y(_2665_));
 sky130_fd_sc_hd__or4_4 _3045_ (.A(\as2650.cycle[7] ),
    .B(\as2650.cycle[6] ),
    .C(\as2650.cycle[5] ),
    .D(\as2650.cycle[4] ),
    .X(_2666_));
 sky130_fd_sc_hd__or4b_4 _3046_ (.A(net289),
    .B(net217),
    .C(net290),
    .D_N(net291),
    .X(_2667_));
 sky130_fd_sc_hd__nor3_4 _3047_ (.A(net289),
    .B(net290),
    .C(_2666_),
    .Y(_2668_));
 sky130_fd_sc_hd__or3_4 _3048_ (.A(net289),
    .B(net290),
    .C(_2666_),
    .X(_2669_));
 sky130_fd_sc_hd__nor2_4 _3049_ (.A(_2666_),
    .B(_2667_),
    .Y(_2670_));
 sky130_fd_sc_hd__or2_2 _3050_ (.A(_2666_),
    .B(_2667_),
    .X(_2671_));
 sky130_fd_sc_hd__and2b_4 _3051_ (.A_N(net298),
    .B(net297),
    .X(_2672_));
 sky130_fd_sc_hd__nand2b_4 _3052_ (.A_N(net298),
    .B(net297),
    .Y(_2673_));
 sky130_fd_sc_hd__and2_4 _3053_ (.A(net308),
    .B(net304),
    .X(_2674_));
 sky130_fd_sc_hd__nand2_1 _3054_ (.A(net308),
    .B(net304),
    .Y(_2675_));
 sky130_fd_sc_hd__and3_4 _3055_ (.A(net173),
    .B(_2672_),
    .C(net209),
    .X(_2676_));
 sky130_fd_sc_hd__or3_4 _3056_ (.A(net210),
    .B(_2673_),
    .C(net208),
    .X(_2677_));
 sky130_fd_sc_hd__and2_1 _3057_ (.A(net301),
    .B(_2676_),
    .X(_2678_));
 sky130_fd_sc_hd__nand2_2 _3058_ (.A(net301),
    .B(_2676_),
    .Y(_2679_));
 sky130_fd_sc_hd__nor2_8 _3059_ (.A(net160),
    .B(net97),
    .Y(_2680_));
 sky130_fd_sc_hd__nand2_2 _3060_ (.A(net159),
    .B(net100),
    .Y(_2681_));
 sky130_fd_sc_hd__or3b_4 _3061_ (.A(_2666_),
    .B(net289),
    .C_N(net290),
    .X(_2682_));
 sky130_fd_sc_hd__nor2_2 _3062_ (.A(net291),
    .B(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__or2_4 _3063_ (.A(net291),
    .B(net293),
    .X(_2684_));
 sky130_fd_sc_hd__or3b_4 _3064_ (.A(net290),
    .B(_2666_),
    .C_N(net289),
    .X(_2685_));
 sky130_fd_sc_hd__nor2_2 _3065_ (.A(net291),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__or2_2 _3066_ (.A(net291),
    .B(_2685_),
    .X(_2687_));
 sky130_fd_sc_hd__nor2_2 _3067_ (.A(_2684_),
    .B(_2685_),
    .Y(_2688_));
 sky130_fd_sc_hd__or3b_4 _3068_ (.A(_2684_),
    .B(\as2650.cycle[3] ),
    .C_N(net290),
    .X(_2689_));
 sky130_fd_sc_hd__nor2_8 _3069_ (.A(_2666_),
    .B(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__or2_2 _3070_ (.A(_2666_),
    .B(_2689_),
    .X(_2691_));
 sky130_fd_sc_hd__nor2_8 _3071_ (.A(_2682_),
    .B(_2684_),
    .Y(_2692_));
 sky130_fd_sc_hd__or2_4 _3072_ (.A(_2682_),
    .B(_2684_),
    .X(_2693_));
 sky130_fd_sc_hd__nand2_4 _3073_ (.A(net157),
    .B(net149),
    .Y(_2694_));
 sky130_fd_sc_hd__o32a_1 _3074_ (.A1(net100),
    .A2(_2688_),
    .A3(_2694_),
    .B1(_2681_),
    .B2(_2683_),
    .X(_2695_));
 sky130_fd_sc_hd__nor2_8 _3075_ (.A(net301),
    .B(net172),
    .Y(_2696_));
 sky130_fd_sc_hd__or2_2 _3076_ (.A(net301),
    .B(net172),
    .X(_2697_));
 sky130_fd_sc_hd__and2_2 _3077_ (.A(net292),
    .B(_2668_),
    .X(_2698_));
 sky130_fd_sc_hd__nand2_2 _3078_ (.A(net292),
    .B(_2668_),
    .Y(_2699_));
 sky130_fd_sc_hd__nor2_2 _3079_ (.A(net293),
    .B(net141),
    .Y(_2700_));
 sky130_fd_sc_hd__nand2_1 _3080_ (.A(net217),
    .B(net143),
    .Y(_2701_));
 sky130_fd_sc_hd__nor2_2 _3081_ (.A(net146),
    .B(net93),
    .Y(_2702_));
 sky130_fd_sc_hd__nand2_2 _3082_ (.A(net291),
    .B(net217),
    .Y(_2703_));
 sky130_fd_sc_hd__nor2_1 _3083_ (.A(_2669_),
    .B(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__or2_4 _3084_ (.A(_2669_),
    .B(_2703_),
    .X(_2705_));
 sky130_fd_sc_hd__or3_2 _3085_ (.A(_2695_),
    .B(_2696_),
    .C(net94),
    .X(_2706_));
 sky130_fd_sc_hd__or4_4 _3086_ (.A(net289),
    .B(net290),
    .C(net291),
    .D(net217),
    .X(_2707_));
 sky130_fd_sc_hd__or3b_4 _3087_ (.A(\as2650.cycle[5] ),
    .B(\as2650.cycle[4] ),
    .C_N(\as2650.cycle[6] ),
    .X(_2708_));
 sky130_fd_sc_hd__nor2_4 _3088_ (.A(_2707_),
    .B(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__or2_4 _3089_ (.A(_2707_),
    .B(_2708_),
    .X(_2710_));
 sky130_fd_sc_hd__nor2_4 _3090_ (.A(_2637_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_1 _3091_ (.A(\as2650.cycle[7] ),
    .B(_2709_),
    .Y(_2712_));
 sky130_fd_sc_hd__or3_4 _3092_ (.A(net289),
    .B(net290),
    .C(_2684_),
    .X(_2713_));
 sky130_fd_sc_hd__nor2_2 _3093_ (.A(_2708_),
    .B(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__or2_4 _3094_ (.A(_2708_),
    .B(_2713_),
    .X(_2715_));
 sky130_fd_sc_hd__nor2_8 _3095_ (.A(\as2650.cycle[7] ),
    .B(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__nand2_2 _3096_ (.A(_2637_),
    .B(net131),
    .Y(_2717_));
 sky130_fd_sc_hd__nor2_8 _3097_ (.A(net85),
    .B(_2716_),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2_4 _3098_ (.A(net84),
    .B(_2717_),
    .Y(_2719_));
 sky130_fd_sc_hd__or4_4 _3099_ (.A(_2637_),
    .B(\as2650.cycle[5] ),
    .C(\as2650.cycle[4] ),
    .D(_2713_),
    .X(_2720_));
 sky130_fd_sc_hd__or3b_1 _3100_ (.A(_2686_),
    .B(_2694_),
    .C_N(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__or2_1 _3101_ (.A(_2719_),
    .B(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__nor2_4 _3102_ (.A(net229),
    .B(net137),
    .Y(_2723_));
 sky130_fd_sc_hd__nand2_2 _3103_ (.A(net212),
    .B(net133),
    .Y(_2724_));
 sky130_fd_sc_hd__a32o_1 _3104_ (.A1(net84),
    .A2(_2722_),
    .A3(net81),
    .B1(_2706_),
    .B2(net173),
    .X(_2725_));
 sky130_fd_sc_hd__nor2_8 _3105_ (.A(net292),
    .B(_2669_),
    .Y(_2726_));
 sky130_fd_sc_hd__nor2_8 _3106_ (.A(_2666_),
    .B(_2707_),
    .Y(_2727_));
 sky130_fd_sc_hd__or2_4 _3107_ (.A(_2666_),
    .B(_2707_),
    .X(_2728_));
 sky130_fd_sc_hd__nor2_2 _3108_ (.A(net230),
    .B(_2687_),
    .Y(_2729_));
 sky130_fd_sc_hd__nor2_1 _3109_ (.A(_2727_),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__nor2_4 _3110_ (.A(_2669_),
    .B(_2684_),
    .Y(_2731_));
 sky130_fd_sc_hd__or2_4 _3111_ (.A(_2669_),
    .B(_2684_),
    .X(_2732_));
 sky130_fd_sc_hd__nand2_4 _3112_ (.A(net213),
    .B(net161),
    .Y(_2733_));
 sky130_fd_sc_hd__nand2_1 _3113_ (.A(net129),
    .B(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__or3_2 _3114_ (.A(_2727_),
    .B(_2729_),
    .C(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__nor2_2 _3115_ (.A(\as2650.cycle[6] ),
    .B(_2720_),
    .Y(_2736_));
 sky130_fd_sc_hd__or2_4 _3116_ (.A(\as2650.cycle[6] ),
    .B(_2720_),
    .X(_2737_));
 sky130_fd_sc_hd__nor2_2 _3117_ (.A(net230),
    .B(_2731_),
    .Y(_2738_));
 sky130_fd_sc_hd__nand2_2 _3118_ (.A(net212),
    .B(net129),
    .Y(_2739_));
 sky130_fd_sc_hd__nand2_2 _3119_ (.A(net79),
    .B(_2738_),
    .Y(_2740_));
 sky130_fd_sc_hd__nor2_8 _3120_ (.A(net303),
    .B(net157),
    .Y(_2741_));
 sky130_fd_sc_hd__or2_4 _3121_ (.A(net301),
    .B(net157),
    .X(_2742_));
 sky130_fd_sc_hd__nand2_2 _3122_ (.A(net144),
    .B(net77),
    .Y(_2743_));
 sky130_fd_sc_hd__nor2_8 _3123_ (.A(_2696_),
    .B(_2741_),
    .Y(_2744_));
 sky130_fd_sc_hd__or2_4 _3124_ (.A(net294),
    .B(net322),
    .X(_2745_));
 sky130_fd_sc_hd__a31o_1 _3125_ (.A1(net145),
    .A2(net132),
    .A3(net77),
    .B1(net210),
    .X(_2746_));
 sky130_fd_sc_hd__nand3_1 _3126_ (.A(_2689_),
    .B(_2740_),
    .C(_2746_),
    .Y(_2747_));
 sky130_fd_sc_hd__or4b_4 _3127_ (.A(_2735_),
    .B(net206),
    .C(_2747_),
    .D_N(_2725_),
    .X(_2748_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(net349),
    .A1(net310),
    .S(_2748_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(net346),
    .A1(\as2650.addr_buff[1] ),
    .S(_2748_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(net342),
    .A1(\as2650.addr_buff[2] ),
    .S(_2748_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(net341),
    .A1(\as2650.addr_buff[3] ),
    .S(_2748_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(net339),
    .A1(\as2650.addr_buff[4] ),
    .S(_2748_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(net337),
    .A1(\as2650.addr_buff[5] ),
    .S(_2748_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(net335),
    .A1(\as2650.addr_buff[6] ),
    .S(_2748_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(net328),
    .A1(net309),
    .S(_2748_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_4 _3136_ (.A(net307),
    .B(net304),
    .Y(_2749_));
 sky130_fd_sc_hd__or2_1 _3137_ (.A(net308),
    .B(net304),
    .X(_2750_));
 sky130_fd_sc_hd__nor2_1 _3138_ (.A(net223),
    .B(net205),
    .Y(_2751_));
 sky130_fd_sc_hd__nand2_1 _3139_ (.A(_2624_),
    .B(net203),
    .Y(_2752_));
 sky130_fd_sc_hd__or2_4 _3140_ (.A(net206),
    .B(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__and2b_4 _3141_ (.A_N(net297),
    .B(\as2650.ins_reg[6] ),
    .X(_2754_));
 sky130_fd_sc_hd__nand2b_4 _3142_ (.A_N(net297),
    .B(\as2650.ins_reg[6] ),
    .Y(_2755_));
 sky130_fd_sc_hd__nor2_8 _3143_ (.A(net300),
    .B(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_8 _3144_ (.A(_2647_),
    .B(_2754_),
    .Y(_2757_));
 sky130_fd_sc_hd__and3b_4 _3145_ (.A_N(net302),
    .B(net234),
    .C(_2756_),
    .X(_2758_));
 sky130_fd_sc_hd__or3_4 _3146_ (.A(net302),
    .B(net213),
    .C(_2757_),
    .X(_2759_));
 sky130_fd_sc_hd__nor2_1 _3147_ (.A(net302),
    .B(net237),
    .Y(_2760_));
 sky130_fd_sc_hd__or2_1 _3148_ (.A(net302),
    .B(net236),
    .X(_2761_));
 sky130_fd_sc_hd__or3_4 _3149_ (.A(net237),
    .B(net90),
    .C(net128),
    .X(_2762_));
 sky130_fd_sc_hd__nand2_8 _3150_ (.A(net298),
    .B(net297),
    .Y(_2763_));
 sky130_fd_sc_hd__or2_4 _3151_ (.A(net299),
    .B(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__nor2_4 _3152_ (.A(net230),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__or2_4 _3153_ (.A(net231),
    .B(_2764_),
    .X(_2766_));
 sky130_fd_sc_hd__nor2_4 _3154_ (.A(net200),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__nand2_1 _3155_ (.A(net202),
    .B(_2765_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand2_4 _3156_ (.A(net233),
    .B(net298),
    .Y(_2769_));
 sky130_fd_sc_hd__and3_4 _3157_ (.A(net234),
    .B(net298),
    .C(net297),
    .X(_2770_));
 sky130_fd_sc_hd__nor2_8 _3158_ (.A(net214),
    .B(_2764_),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_4 _3159_ (.A(_2647_),
    .B(_2770_),
    .Y(_2772_));
 sky130_fd_sc_hd__nor2_4 _3160_ (.A(net302),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__or2_2 _3161_ (.A(net303),
    .B(_2772_),
    .X(_2774_));
 sky130_fd_sc_hd__nor2_1 _3162_ (.A(net199),
    .B(_2772_),
    .Y(_2775_));
 sky130_fd_sc_hd__or2_4 _3163_ (.A(net199),
    .B(_2772_),
    .X(_2776_));
 sky130_fd_sc_hd__nor3_2 _3164_ (.A(net91),
    .B(_2753_),
    .C(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(net233),
    .B(net206),
    .Y(_2778_));
 sky130_fd_sc_hd__or2_4 _3166_ (.A(net233),
    .B(net206),
    .X(_2779_));
 sky130_fd_sc_hd__nor2_8 _3167_ (.A(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_2780_));
 sky130_fd_sc_hd__nand2_1 _3168_ (.A(_2648_),
    .B(net85),
    .Y(_2781_));
 sky130_fd_sc_hd__nor2_4 _3169_ (.A(\as2650.cycle[7] ),
    .B(_2710_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_8 _3170_ (.A(_2637_),
    .B(_2709_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor2_8 _3171_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_2784_));
 sky130_fd_sc_hd__or2_1 _3172_ (.A(\as2650.idx_ctrl[1] ),
    .B(\as2650.idx_ctrl[0] ),
    .X(_2785_));
 sky130_fd_sc_hd__nor2_1 _3173_ (.A(_2779_),
    .B(_2784_),
    .Y(_2786_));
 sky130_fd_sc_hd__nand2_1 _3174_ (.A(_2778_),
    .B(net197),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2_8 _3175_ (.A(net231),
    .B(net299),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_4 _3176_ (.A(net302),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__or2_4 _3177_ (.A(net302),
    .B(_2788_),
    .X(_2790_));
 sky130_fd_sc_hd__nor2_4 _3178_ (.A(net297),
    .B(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__or2_4 _3179_ (.A(\as2650.ins_reg[7] ),
    .B(_2790_),
    .X(_2792_));
 sky130_fd_sc_hd__nor2_2 _3180_ (.A(net236),
    .B(net213),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_8 _3181_ (.A(net215),
    .B(net233),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _3182_ (.A(net216),
    .B(net126),
    .Y(_2795_));
 sky130_fd_sc_hd__or2_4 _3183_ (.A(net158),
    .B(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__nor2_1 _3184_ (.A(_2753_),
    .B(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__or2_4 _3185_ (.A(_2753_),
    .B(_2796_),
    .X(_2798_));
 sky130_fd_sc_hd__nor2_4 _3186_ (.A(_2647_),
    .B(_2763_),
    .Y(_2799_));
 sky130_fd_sc_hd__nand2_1 _3187_ (.A(net204),
    .B(net198),
    .Y(_2800_));
 sky130_fd_sc_hd__or4_1 _3188_ (.A(net151),
    .B(net197),
    .C(_2799_),
    .D(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__or2_4 _3189_ (.A(net223),
    .B(net206),
    .X(_2802_));
 sky130_fd_sc_hd__nand2_4 _3190_ (.A(net205),
    .B(net202),
    .Y(_2803_));
 sky130_fd_sc_hd__nor2_8 _3191_ (.A(net298),
    .B(\as2650.ins_reg[7] ),
    .Y(_2804_));
 sky130_fd_sc_hd__nand2_1 _3192_ (.A(net233),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__or2_4 _3193_ (.A(net299),
    .B(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__nor2_2 _3194_ (.A(_2803_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__or2_2 _3195_ (.A(_2803_),
    .B(_2806_),
    .X(_2808_));
 sky130_fd_sc_hd__or3_4 _3196_ (.A(net214),
    .B(net300),
    .C(_2673_),
    .X(_2809_));
 sky130_fd_sc_hd__nand2_4 _3197_ (.A(net306),
    .B(_2644_),
    .Y(_2810_));
 sky130_fd_sc_hd__or3_1 _3198_ (.A(net198),
    .B(_2809_),
    .C(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__and2_2 _3199_ (.A(net73),
    .B(net124),
    .X(_2812_));
 sky130_fd_sc_hd__nand2_8 _3200_ (.A(net74),
    .B(net125),
    .Y(_2813_));
 sky130_fd_sc_hd__or3_4 _3201_ (.A(net90),
    .B(_2802_),
    .C(_2812_),
    .X(_2814_));
 sky130_fd_sc_hd__nand2_4 _3202_ (.A(net216),
    .B(net96),
    .Y(_2815_));
 sky130_fd_sc_hd__or3_2 _3203_ (.A(_2753_),
    .B(net127),
    .C(_2815_),
    .X(_2816_));
 sky130_fd_sc_hd__inv_2 _3204_ (.A(net57),
    .Y(_2817_));
 sky130_fd_sc_hd__or4_4 _3205_ (.A(net91),
    .B(net205),
    .C(_2768_),
    .D(_2802_),
    .X(_2818_));
 sky130_fd_sc_hd__nor2_8 _3206_ (.A(net309),
    .B(_2780_),
    .Y(_2819_));
 sky130_fd_sc_hd__or2_4 _3207_ (.A(net309),
    .B(_2780_),
    .X(_2820_));
 sky130_fd_sc_hd__or4_4 _3208_ (.A(net83),
    .B(_2752_),
    .C(_2779_),
    .D(_2820_),
    .X(_2821_));
 sky130_fd_sc_hd__or3_1 _3209_ (.A(_2752_),
    .B(_2783_),
    .C(_2787_),
    .X(_2822_));
 sky130_fd_sc_hd__and4_1 _3210_ (.A(_2798_),
    .B(_2818_),
    .C(_2821_),
    .D(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__nor2_4 _3211_ (.A(_2753_),
    .B(_2762_),
    .Y(_2824_));
 sky130_fd_sc_hd__or2_4 _3212_ (.A(_2753_),
    .B(_2762_),
    .X(_2825_));
 sky130_fd_sc_hd__nor2_4 _3213_ (.A(net215),
    .B(net89),
    .Y(_2826_));
 sky130_fd_sc_hd__nand2_8 _3214_ (.A(net237),
    .B(net93),
    .Y(_2827_));
 sky130_fd_sc_hd__or2_2 _3215_ (.A(_2799_),
    .B(_2800_),
    .X(_2828_));
 sky130_fd_sc_hd__or4_1 _3216_ (.A(net233),
    .B(net150),
    .C(net196),
    .D(_2828_),
    .X(_2829_));
 sky130_fd_sc_hd__o32a_1 _3217_ (.A1(_2753_),
    .A2(_2769_),
    .A3(_2827_),
    .B1(_2829_),
    .B2(_2802_),
    .X(_2830_));
 sky130_fd_sc_hd__and4_4 _3218_ (.A(net57),
    .B(_2823_),
    .C(_2825_),
    .D(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__or2_4 _3219_ (.A(net304),
    .B(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__inv_2 _3220_ (.A(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__or4_4 _3221_ (.A(net233),
    .B(net147),
    .C(net197),
    .D(_2828_),
    .X(_2834_));
 sky130_fd_sc_hd__nor2_4 _3222_ (.A(_2802_),
    .B(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__or2_4 _3223_ (.A(_2802_),
    .B(_2834_),
    .X(_2836_));
 sky130_fd_sc_hd__nor2_1 _3224_ (.A(net134),
    .B(_2802_),
    .Y(_2837_));
 sky130_fd_sc_hd__and3_1 _3225_ (.A(net203),
    .B(_2775_),
    .C(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__and4_4 _3226_ (.A(net85),
    .B(_2751_),
    .C(_2778_),
    .D(_2819_),
    .X(_2839_));
 sky130_fd_sc_hd__and3_4 _3227_ (.A(_2751_),
    .B(_2782_),
    .C(_2786_),
    .X(_2840_));
 sky130_fd_sc_hd__or3_4 _3228_ (.A(_2752_),
    .B(_2783_),
    .C(_2787_),
    .X(_2841_));
 sky130_fd_sc_hd__and3_4 _3229_ (.A(net203),
    .B(_2767_),
    .C(_2837_),
    .X(_2842_));
 sky130_fd_sc_hd__and3_4 _3230_ (.A(net318),
    .B(_2814_),
    .C(_2832_),
    .X(_2843_));
 sky130_fd_sc_hd__nand3_4 _3231_ (.A(net321),
    .B(_2814_),
    .C(_2832_),
    .Y(_2844_));
 sky130_fd_sc_hd__nor2_2 _3232_ (.A(net89),
    .B(net73),
    .Y(_2845_));
 sky130_fd_sc_hd__or3_4 _3233_ (.A(net90),
    .B(_2802_),
    .C(net73),
    .X(_2846_));
 sky130_fd_sc_hd__nor2_4 _3234_ (.A(net224),
    .B(net225),
    .Y(_2847_));
 sky130_fd_sc_hd__or2_2 _3235_ (.A(net224),
    .B(net225),
    .X(_2848_));
 sky130_fd_sc_hd__nor2_8 _3236_ (.A(net228),
    .B(_2847_),
    .Y(_2849_));
 sky130_fd_sc_hd__nand2_8 _3237_ (.A(net227),
    .B(net195),
    .Y(_2850_));
 sky130_fd_sc_hd__and3_1 _3238_ (.A(net228),
    .B(\as2650.stack[3][8] ),
    .C(net195),
    .X(_2851_));
 sky130_fd_sc_hd__or2_4 _3239_ (.A(_2626_),
    .B(net225),
    .X(_2852_));
 sky130_fd_sc_hd__nand2_1 _3240_ (.A(_2626_),
    .B(net225),
    .Y(_2853_));
 sky130_fd_sc_hd__nand2_4 _3241_ (.A(net224),
    .B(net225),
    .Y(_2854_));
 sky130_fd_sc_hd__and2_1 _3242_ (.A(net193),
    .B(net192),
    .X(_2855_));
 sky130_fd_sc_hd__nand2_1 _3243_ (.A(net193),
    .B(net192),
    .Y(_2856_));
 sky130_fd_sc_hd__o22a_1 _3244_ (.A1(\as2650.stack[0][8] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[1][8] ),
    .X(_2857_));
 sky130_fd_sc_hd__and2b_4 _3245_ (.A_N(_2849_),
    .B(_2850_),
    .X(_2858_));
 sky130_fd_sc_hd__nand2b_4 _3246_ (.A_N(_2849_),
    .B(_2850_),
    .Y(_2859_));
 sky130_fd_sc_hd__o221a_1 _3247_ (.A1(_2849_),
    .A2(_2851_),
    .B1(net191),
    .B2(\as2650.stack[2][8] ),
    .C1(_2857_),
    .X(_2860_));
 sky130_fd_sc_hd__o22a_1 _3248_ (.A1(\as2650.stack[7][8] ),
    .A2(net194),
    .B1(net192),
    .B2(\as2650.stack[6][8] ),
    .X(_2861_));
 sky130_fd_sc_hd__o22a_1 _3249_ (.A1(\as2650.stack[4][8] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[5][8] ),
    .X(_2862_));
 sky130_fd_sc_hd__a31o_4 _3250_ (.A1(net123),
    .A2(_2861_),
    .A3(_2862_),
    .B1(_2860_),
    .X(_2863_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(_2629_),
    .B(_2846_),
    .Y(_2864_));
 sky130_fd_sc_hd__or2_4 _3252_ (.A(_2803_),
    .B(_2809_),
    .X(_2865_));
 sky130_fd_sc_hd__nor3_2 _3253_ (.A(net90),
    .B(_2802_),
    .C(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__or3_4 _3254_ (.A(net90),
    .B(_2802_),
    .C(_2865_),
    .X(_2867_));
 sky130_fd_sc_hd__nand2_4 _3255_ (.A(_2814_),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__o211a_1 _3256_ (.A1(_2846_),
    .A2(_2863_),
    .B1(_2864_),
    .C1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__nor2_1 _3257_ (.A(_2624_),
    .B(net205),
    .Y(_2870_));
 sky130_fd_sc_hd__nand2_2 _3258_ (.A(net223),
    .B(net203),
    .Y(_2871_));
 sky130_fd_sc_hd__mux4_2 _3259_ (.A0(\as2650.r123[1][0] ),
    .A1(\as2650.r123[0][0] ),
    .A2(\as2650.r123_2[1][0] ),
    .A3(\as2650.r123_2[0][0] ),
    .S0(net307),
    .S1(net220),
    .X(_2872_));
 sky130_fd_sc_hd__mux2_8 _3260_ (.A0(\as2650.r123[2][0] ),
    .A1(\as2650.r123_2[2][0] ),
    .S(net221),
    .X(_2873_));
 sky130_fd_sc_hd__and2_4 _3261_ (.A(net209),
    .B(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__nand2_4 _3262_ (.A(net209),
    .B(_2873_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor3b_4 _3263_ (.A(net308),
    .B(\as2650.ins_reg[1] ),
    .C_N(net266),
    .Y(_2876_));
 sky130_fd_sc_hd__a31oi_4 _3264_ (.A1(net207),
    .A2(net204),
    .A3(_2872_),
    .B1(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__a31o_4 _3265_ (.A1(net207),
    .A2(net204),
    .A3(_2872_),
    .B1(_2876_),
    .X(_2878_));
 sky130_fd_sc_hd__nor2_8 _3266_ (.A(_2874_),
    .B(_2878_),
    .Y(_2879_));
 sky130_fd_sc_hd__nand2_8 _3267_ (.A(_2875_),
    .B(_2877_),
    .Y(_2880_));
 sky130_fd_sc_hd__xnor2_4 _3268_ (.A(_2770_),
    .B(net121),
    .Y(_2881_));
 sky130_fd_sc_hd__nor2_1 _3269_ (.A(net58),
    .B(_2881_),
    .Y(_2882_));
 sky130_fd_sc_hd__mux4_2 _3270_ (.A0(\as2650.r123[1][1] ),
    .A1(\as2650.r123[0][1] ),
    .A2(\as2650.r123_2[1][1] ),
    .A3(\as2650.r123_2[0][1] ),
    .S0(net307),
    .S1(net222),
    .X(_2883_));
 sky130_fd_sc_hd__and3_1 _3271_ (.A(net208),
    .B(net204),
    .C(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__mux2_8 _3272_ (.A0(\as2650.r123[2][1] ),
    .A1(\as2650.r123_2[2][1] ),
    .S(net221),
    .X(_2885_));
 sky130_fd_sc_hd__a22o_2 _3273_ (.A1(net263),
    .A2(net205),
    .B1(_2885_),
    .B2(net209),
    .X(_2886_));
 sky130_fd_sc_hd__or2_4 _3274_ (.A(_2884_),
    .B(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__a211o_1 _3275_ (.A1(net347),
    .A2(net58),
    .B1(_2824_),
    .C1(_2882_),
    .X(_2888_));
 sky130_fd_sc_hd__o211a_1 _3276_ (.A1(_2825_),
    .A2(net119),
    .B1(_2888_),
    .C1(net57),
    .X(_2889_));
 sky130_fd_sc_hd__nand2b_2 _3277_ (.A_N(\as2650.carry ),
    .B(\as2650.psl[3] ),
    .Y(_2890_));
 sky130_fd_sc_hd__mux2_4 _3278_ (.A0(\as2650.r123[2][7] ),
    .A1(\as2650.r123_2[2][7] ),
    .S(net221),
    .X(_2891_));
 sky130_fd_sc_hd__a22o_4 _3279_ (.A1(net241),
    .A2(net205),
    .B1(_2891_),
    .B2(net209),
    .X(_2892_));
 sky130_fd_sc_hd__mux2_8 _3280_ (.A0(\as2650.r123[0][7] ),
    .A1(\as2650.r123_2[0][7] ),
    .S(net220),
    .X(_2893_));
 sky130_fd_sc_hd__mux4_1 _3281_ (.A0(\as2650.r123[1][7] ),
    .A1(\as2650.r123[0][7] ),
    .A2(\as2650.r123_2[1][7] ),
    .A3(\as2650.r123_2[0][7] ),
    .S0(net307),
    .S1(net220),
    .X(_2894_));
 sky130_fd_sc_hd__and3_4 _3282_ (.A(net207),
    .B(net203),
    .C(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__nor2_8 _3283_ (.A(_2892_),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__or2_4 _3284_ (.A(_2892_),
    .B(_2895_),
    .X(_2897_));
 sky130_fd_sc_hd__nand2_2 _3285_ (.A(\as2650.psl[3] ),
    .B(\as2650.carry ),
    .Y(_2898_));
 sky130_fd_sc_hd__o21a_2 _3286_ (.A1(\as2650.psl[3] ),
    .A2(_2897_),
    .B1(_2890_),
    .X(_2899_));
 sky130_fd_sc_hd__inv_2 _3287_ (.A(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__a211o_1 _3288_ (.A1(_2777_),
    .A2(_2899_),
    .B1(_2889_),
    .C1(_2842_),
    .X(_2901_));
 sky130_fd_sc_hd__o211a_1 _3289_ (.A1(net266),
    .A2(_2818_),
    .B1(_2821_),
    .C1(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__nand2b_4 _3290_ (.A_N(\as2650.addr_buff[6] ),
    .B(\as2650.addr_buff[5] ),
    .Y(_2903_));
 sky130_fd_sc_hd__nand2b_4 _3291_ (.A_N(\as2650.addr_buff[5] ),
    .B(\as2650.addr_buff[6] ),
    .Y(_2904_));
 sky130_fd_sc_hd__nand2_8 _3292_ (.A(_2903_),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_4 _3293_ (.A(_2879_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__a211o_1 _3294_ (.A1(_2839_),
    .A2(_2906_),
    .B1(_2902_),
    .C1(_2840_),
    .X(_2907_));
 sky130_fd_sc_hd__nor2_1 _3295_ (.A(\as2650.idx_ctrl[1] ),
    .B(_2640_),
    .Y(_2908_));
 sky130_fd_sc_hd__nand2_8 _3296_ (.A(_2639_),
    .B(\as2650.idx_ctrl[0] ),
    .Y(_2909_));
 sky130_fd_sc_hd__nand2_8 _3297_ (.A(\as2650.idx_ctrl[1] ),
    .B(_2640_),
    .Y(_2910_));
 sky130_fd_sc_hd__nand2_8 _3298_ (.A(_2909_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__xnor2_4 _3299_ (.A(_2879_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__o21a_1 _3300_ (.A1(_2841_),
    .A2(_2912_),
    .B1(_2907_),
    .X(_2913_));
 sky130_fd_sc_hd__and2_4 _3301_ (.A(net299),
    .B(_2804_),
    .X(_2914_));
 sky130_fd_sc_hd__nand2_8 _3302_ (.A(net299),
    .B(_2804_),
    .Y(_2915_));
 sky130_fd_sc_hd__and2_1 _3303_ (.A(\as2650.holding_reg[0] ),
    .B(net121),
    .X(_2916_));
 sky130_fd_sc_hd__or2_1 _3304_ (.A(\as2650.holding_reg[0] ),
    .B(net202),
    .X(_2917_));
 sky130_fd_sc_hd__o31a_4 _3305_ (.A1(net199),
    .A2(_2874_),
    .A3(_2878_),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__nor2_1 _3306_ (.A(\as2650.holding_reg[0] ),
    .B(net199),
    .Y(_2919_));
 sky130_fd_sc_hd__a31o_4 _3307_ (.A1(net199),
    .A2(_2875_),
    .A3(_2877_),
    .B1(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__inv_2 _3308_ (.A(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__and2_1 _3309_ (.A(_2918_),
    .B(_2920_),
    .X(_2922_));
 sky130_fd_sc_hd__xor2_4 _3310_ (.A(_2918_),
    .B(_2920_),
    .X(_2923_));
 sky130_fd_sc_hd__inv_2 _3311_ (.A(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__nor2_4 _3312_ (.A(net299),
    .B(_2673_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_2 _3313_ (.A(_2647_),
    .B(_2672_),
    .Y(_2926_));
 sky130_fd_sc_hd__o21ai_1 _3314_ (.A1(_2898_),
    .A2(_2923_),
    .B1(_2925_),
    .Y(_2927_));
 sky130_fd_sc_hd__a21oi_1 _3315_ (.A1(_2898_),
    .A2(_2923_),
    .B1(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_1 _3316_ (.A(_2890_),
    .B(_2923_),
    .Y(_2929_));
 sky130_fd_sc_hd__nand2_4 _3317_ (.A(net300),
    .B(_2672_),
    .Y(_2930_));
 sky130_fd_sc_hd__o2111a_1 _3318_ (.A1(_2890_),
    .A2(_2923_),
    .B1(_2929_),
    .C1(_2672_),
    .D1(net300),
    .X(_2931_));
 sky130_fd_sc_hd__a221o_1 _3319_ (.A1(_2673_),
    .A2(_2918_),
    .B1(_2921_),
    .B2(_2754_),
    .C1(_2756_),
    .X(_2932_));
 sky130_fd_sc_hd__o32a_1 _3320_ (.A1(_2928_),
    .A2(_2931_),
    .A3(_2932_),
    .B1(_2916_),
    .B2(_2757_),
    .X(_2933_));
 sky130_fd_sc_hd__mux2_8 _3321_ (.A0(_2924_),
    .A1(_2933_),
    .S(_2915_),
    .X(_2934_));
 sky130_fd_sc_hd__mux2_4 _3322_ (.A0(_2913_),
    .A1(_2934_),
    .S(_2835_),
    .X(_2935_));
 sky130_fd_sc_hd__a211o_1 _3323_ (.A1(_2833_),
    .A2(_2935_),
    .B1(_2869_),
    .C1(_2843_),
    .X(_2936_));
 sky130_fd_sc_hd__nand2_4 _3324_ (.A(_2812_),
    .B(_2865_),
    .Y(_2937_));
 sky130_fd_sc_hd__o21a_1 _3325_ (.A1(\as2650.r123[0][0] ),
    .A2(_2844_),
    .B1(_2936_),
    .X(_0008_));
 sky130_fd_sc_hd__and3_1 _3326_ (.A(net228),
    .B(\as2650.stack[3][9] ),
    .C(net195),
    .X(_2938_));
 sky130_fd_sc_hd__o22a_1 _3327_ (.A1(\as2650.stack[0][9] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[1][9] ),
    .X(_2939_));
 sky130_fd_sc_hd__o221a_2 _3328_ (.A1(\as2650.stack[2][9] ),
    .A2(net191),
    .B1(_2938_),
    .B2(_2849_),
    .C1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__mux4_2 _3329_ (.A0(\as2650.stack[7][9] ),
    .A1(\as2650.stack[4][9] ),
    .A2(\as2650.stack[5][9] ),
    .A3(\as2650.stack[6][9] ),
    .S0(net224),
    .S1(net225),
    .X(_2941_));
 sky130_fd_sc_hd__a21oi_4 _3330_ (.A1(net123),
    .A2(_2941_),
    .B1(_2940_),
    .Y(_2942_));
 sky130_fd_sc_hd__inv_2 _3331_ (.A(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o221a_1 _3332_ (.A1(net264),
    .A2(net75),
    .B1(_2846_),
    .B2(_2943_),
    .C1(_2868_),
    .X(_2944_));
 sky130_fd_sc_hd__nor2_8 _3333_ (.A(_2763_),
    .B(_2788_),
    .Y(_2945_));
 sky130_fd_sc_hd__mux2_4 _3334_ (.A0(_2771_),
    .A1(_2945_),
    .S(_2879_),
    .X(_2946_));
 sky130_fd_sc_hd__xor2_4 _3335_ (.A(net119),
    .B(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__mux2_8 _3336_ (.A0(\as2650.r123[2][2] ),
    .A1(\as2650.r123_2[2][2] ),
    .S(net221),
    .X(_2948_));
 sky130_fd_sc_hd__mux2_2 _3337_ (.A0(\as2650.r123[0][2] ),
    .A1(\as2650.r123_2[0][2] ),
    .S(net221),
    .X(_2949_));
 sky130_fd_sc_hd__mux4_1 _3338_ (.A0(\as2650.r123[1][2] ),
    .A1(\as2650.r123[0][2] ),
    .A2(\as2650.r123_2[1][2] ),
    .A3(\as2650.r123_2[0][2] ),
    .S0(net307),
    .S1(net222),
    .X(_2950_));
 sky130_fd_sc_hd__and3_1 _3339_ (.A(net207),
    .B(net203),
    .C(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__a221o_2 _3340_ (.A1(net258),
    .A2(net205),
    .B1(_2948_),
    .B2(net209),
    .C1(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__or2_1 _3341_ (.A(net58),
    .B(_2947_),
    .X(_2953_));
 sky130_fd_sc_hd__o211a_1 _3342_ (.A1(net346),
    .A2(_2798_),
    .B1(_2825_),
    .C1(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__a211o_1 _3343_ (.A1(_2824_),
    .A2(net116),
    .B1(_2954_),
    .C1(_2817_),
    .X(_2955_));
 sky130_fd_sc_hd__o211a_1 _3344_ (.A1(net57),
    .A2(net121),
    .B1(_2955_),
    .C1(_2818_),
    .X(_2956_));
 sky130_fd_sc_hd__a21o_1 _3345_ (.A1(net263),
    .A2(_2842_),
    .B1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__o22a_4 _3346_ (.A1(_2874_),
    .A2(_2878_),
    .B1(_2884_),
    .B2(_2886_),
    .X(_2958_));
 sky130_fd_sc_hd__nor2_1 _3347_ (.A(_2880_),
    .B(net119),
    .Y(_2959_));
 sky130_fd_sc_hd__xnor2_4 _3348_ (.A(net121),
    .B(net119),
    .Y(_2960_));
 sky130_fd_sc_hd__a21bo_2 _3349_ (.A1(net121),
    .A2(_2903_),
    .B1_N(_2904_),
    .X(_2961_));
 sky130_fd_sc_hd__xnor2_4 _3350_ (.A(_2960_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(_2957_),
    .A1(_2962_),
    .S(_2839_),
    .X(_2963_));
 sky130_fd_sc_hd__o21a_2 _3352_ (.A1(_2879_),
    .A2(_2908_),
    .B1(_2910_),
    .X(_2964_));
 sky130_fd_sc_hd__xor2_4 _3353_ (.A(_2960_),
    .B(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__o21a_1 _3354_ (.A1(_2841_),
    .A2(_2965_),
    .B1(_2836_),
    .X(_2966_));
 sky130_fd_sc_hd__o21ai_1 _3355_ (.A1(_2840_),
    .A2(_2963_),
    .B1(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__and2_4 _3356_ (.A(\as2650.holding_reg[1] ),
    .B(net120),
    .X(_2968_));
 sky130_fd_sc_hd__nor2_4 _3357_ (.A(\as2650.holding_reg[1] ),
    .B(net120),
    .Y(_2969_));
 sky130_fd_sc_hd__nor2_8 _3358_ (.A(_2968_),
    .B(_2969_),
    .Y(_2970_));
 sky130_fd_sc_hd__o2bb2a_2 _3359_ (.A1_N(_2890_),
    .A2_N(_2923_),
    .B1(_2916_),
    .B2(_2920_),
    .X(_2971_));
 sky130_fd_sc_hd__or2_1 _3360_ (.A(_2970_),
    .B(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__nand2_1 _3361_ (.A(_2970_),
    .B(_2971_),
    .Y(_2973_));
 sky130_fd_sc_hd__a21o_1 _3362_ (.A1(_2972_),
    .A2(_2973_),
    .B1(_2930_),
    .X(_2974_));
 sky130_fd_sc_hd__o21bai_4 _3363_ (.A1(_2898_),
    .A2(_2923_),
    .B1_N(_2916_),
    .Y(_2975_));
 sky130_fd_sc_hd__xor2_1 _3364_ (.A(_2970_),
    .B(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__nand2_2 _3365_ (.A(net300),
    .B(_2754_),
    .Y(_2977_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(\as2650.holding_reg[1] ),
    .A1(net120),
    .S(net201),
    .X(_2978_));
 sky130_fd_sc_hd__o22a_1 _3367_ (.A1(_2926_),
    .A2(_2976_),
    .B1(_2978_),
    .B2(_2672_),
    .X(_2979_));
 sky130_fd_sc_hd__a21oi_1 _3368_ (.A1(net300),
    .A2(_2969_),
    .B1(_2755_),
    .Y(_2980_));
 sky130_fd_sc_hd__a31o_1 _3369_ (.A1(_2974_),
    .A2(_2977_),
    .A3(_2979_),
    .B1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__o21a_4 _3370_ (.A1(_2757_),
    .A2(_2968_),
    .B1(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__or2_2 _3371_ (.A(\as2650.holding_reg[1] ),
    .B(net199),
    .X(_2983_));
 sky130_fd_sc_hd__o21ai_4 _3372_ (.A1(net201),
    .A2(net120),
    .B1(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__or2_4 _3373_ (.A(_2915_),
    .B(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__xnor2_4 _3374_ (.A(_2982_),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__a21bo_4 _3375_ (.A1(_2835_),
    .A2(_2986_),
    .B1_N(_2967_),
    .X(_2987_));
 sky130_fd_sc_hd__a211o_1 _3376_ (.A1(_2833_),
    .A2(_2987_),
    .B1(_2944_),
    .C1(_2843_),
    .X(_2988_));
 sky130_fd_sc_hd__o21a_1 _3377_ (.A1(\as2650.r123[0][1] ),
    .A2(_2844_),
    .B1(_2988_),
    .X(_0009_));
 sky130_fd_sc_hd__and3_1 _3378_ (.A(net228),
    .B(\as2650.stack[3][10] ),
    .C(net195),
    .X(_2989_));
 sky130_fd_sc_hd__o22a_1 _3379_ (.A1(\as2650.stack[0][10] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[1][10] ),
    .X(_2990_));
 sky130_fd_sc_hd__o221a_1 _3380_ (.A1(\as2650.stack[2][10] ),
    .A2(net191),
    .B1(_2989_),
    .B2(_2849_),
    .C1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__mux4_1 _3381_ (.A0(\as2650.stack[7][10] ),
    .A1(\as2650.stack[4][10] ),
    .A2(\as2650.stack[5][10] ),
    .A3(\as2650.stack[6][10] ),
    .S0(net224),
    .S1(net225),
    .X(_2992_));
 sky130_fd_sc_hd__a21o_2 _3382_ (.A1(net122),
    .A2(_2992_),
    .B1(_2991_),
    .X(_2993_));
 sky130_fd_sc_hd__o221a_1 _3383_ (.A1(net259),
    .A2(net75),
    .B1(_2846_),
    .B2(_2993_),
    .C1(_2868_),
    .X(_2994_));
 sky130_fd_sc_hd__or2_1 _3384_ (.A(_2843_),
    .B(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__a22o_2 _3385_ (.A1(_2771_),
    .A2(_2958_),
    .B1(_2959_),
    .B2(_2945_),
    .X(_2996_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(net115),
    .B(_2958_),
    .Y(_2997_));
 sky130_fd_sc_hd__and3_2 _3387_ (.A(_2771_),
    .B(net114),
    .C(_2958_),
    .X(_2998_));
 sky130_fd_sc_hd__nor3_4 _3388_ (.A(net121),
    .B(net120),
    .C(net114),
    .Y(_2999_));
 sky130_fd_sc_hd__xnor2_4 _3389_ (.A(net114),
    .B(_2996_),
    .Y(_3000_));
 sky130_fd_sc_hd__inv_2 _3390_ (.A(_3000_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _3391_ (.A(net58),
    .B(_3000_),
    .Y(_0301_));
 sky130_fd_sc_hd__a211o_1 _3392_ (.A1(net344),
    .A2(net58),
    .B1(_2824_),
    .C1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_4 _3393_ (.A0(\as2650.r123[2][3] ),
    .A1(\as2650.r123_2[2][3] ),
    .S(net221),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_2 _3394_ (.A0(\as2650.r123[0][3] ),
    .A1(\as2650.r123_2[0][3] ),
    .S(net220),
    .X(_0304_));
 sky130_fd_sc_hd__mux4_1 _3395_ (.A0(\as2650.r123[1][3] ),
    .A1(\as2650.r123[0][3] ),
    .A2(\as2650.r123_2[1][3] ),
    .A3(\as2650.r123_2[0][3] ),
    .S0(net307),
    .S1(net220),
    .X(_0305_));
 sky130_fd_sc_hd__and3_1 _3396_ (.A(net207),
    .B(net203),
    .C(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_2 _3397_ (.A1(net255),
    .A2(net205),
    .B1(_0303_),
    .B2(net209),
    .C1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _3398_ (.A(_2825_),
    .B(net113),
    .X(_0308_));
 sky130_fd_sc_hd__o21a_1 _3399_ (.A1(net121),
    .A2(net120),
    .B1(net114),
    .X(_0309_));
 sky130_fd_sc_hd__xor2_2 _3400_ (.A(net114),
    .B(_2958_),
    .X(_0310_));
 sky130_fd_sc_hd__o32a_1 _3401_ (.A1(_2904_),
    .A2(_2999_),
    .A3(_0309_),
    .B1(_0310_),
    .B2(_2903_),
    .X(_0311_));
 sky130_fd_sc_hd__o21a_4 _3402_ (.A1(_2905_),
    .A2(net114),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a32o_1 _3403_ (.A1(net57),
    .A2(_0302_),
    .A3(_0308_),
    .B1(_2838_),
    .B2(net119),
    .X(_0313_));
 sky130_fd_sc_hd__o221a_1 _3404_ (.A1(net258),
    .A2(_2818_),
    .B1(_2842_),
    .B2(_0313_),
    .C1(_2821_),
    .X(_0314_));
 sky130_fd_sc_hd__or3_1 _3405_ (.A(_2910_),
    .B(_2999_),
    .C(_0309_),
    .X(_0315_));
 sky130_fd_sc_hd__o221a_4 _3406_ (.A1(_2911_),
    .A2(net114),
    .B1(_0310_),
    .B2(_2909_),
    .C1(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a211o_1 _3407_ (.A1(_2839_),
    .A2(_0312_),
    .B1(_0314_),
    .C1(_2840_),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _3408_ (.A1(_2841_),
    .A2(_0316_),
    .B1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_2 _3409_ (.A(\as2650.holding_reg[2] ),
    .B(net116),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_2 _3410_ (.A(\as2650.holding_reg[2] ),
    .B(net116),
    .Y(_0320_));
 sky130_fd_sc_hd__nor2_2 _3411_ (.A(_0319_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _3412_ (.A(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__o22ai_4 _3413_ (.A1(_2970_),
    .A2(_2971_),
    .B1(_2984_),
    .B2(_2968_),
    .Y(_0323_));
 sky130_fd_sc_hd__xnor2_1 _3414_ (.A(_0321_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_2 _3415_ (.A1(_2970_),
    .A2(_2975_),
    .B1(_2968_),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_1 _3416_ (.A(_0321_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\as2650.holding_reg[2] ),
    .A1(net116),
    .S(net201),
    .X(_0327_));
 sky130_fd_sc_hd__o221a_1 _3418_ (.A1(_2926_),
    .A2(_0326_),
    .B1(_0327_),
    .B2(_2672_),
    .C1(_2977_),
    .X(_0328_));
 sky130_fd_sc_hd__o21ai_1 _3419_ (.A1(_2930_),
    .A2(_0324_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__o211a_1 _3420_ (.A1(_2977_),
    .A2(_0320_),
    .B1(_0329_),
    .C1(_2757_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_1 _3421_ (.A(_2757_),
    .B(_0319_),
    .Y(_0331_));
 sky130_fd_sc_hd__or3_2 _3422_ (.A(_2914_),
    .B(_0330_),
    .C(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__o21ai_4 _3423_ (.A1(_2915_),
    .A2(_0322_),
    .B1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__mux2_4 _3424_ (.A0(_0318_),
    .A1(_0333_),
    .S(_2835_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _3425_ (.A(_2833_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o22a_1 _3426_ (.A1(\as2650.r123[0][2] ),
    .A2(_2844_),
    .B1(_2995_),
    .B2(_0335_),
    .X(_0010_));
 sky130_fd_sc_hd__o22a_1 _3427_ (.A1(\as2650.stack[3][11] ),
    .A2(net194),
    .B1(net165),
    .B2(\as2650.stack[1][11] ),
    .X(_0336_));
 sky130_fd_sc_hd__o221a_2 _3428_ (.A1(\as2650.stack[0][11] ),
    .A2(net169),
    .B1(net191),
    .B2(\as2650.stack[2][11] ),
    .C1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o221a_1 _3429_ (.A1(\as2650.stack[4][11] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[5][11] ),
    .C1(net122),
    .X(_0338_));
 sky130_fd_sc_hd__o221a_2 _3430_ (.A1(\as2650.stack[7][11] ),
    .A2(net194),
    .B1(net192),
    .B2(\as2650.stack[6][11] ),
    .C1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__a21oi_4 _3431_ (.A1(_2859_),
    .A2(_0337_),
    .B1(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _3432_ (.A(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__o221a_1 _3433_ (.A1(net256),
    .A2(net75),
    .B1(_2846_),
    .B2(_0341_),
    .C1(_2868_),
    .X(_0342_));
 sky130_fd_sc_hd__a21oi_4 _3434_ (.A1(_2945_),
    .A2(_2999_),
    .B1(_2998_),
    .Y(_0343_));
 sky130_fd_sc_hd__xnor2_4 _3435_ (.A(net111),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__or2_1 _3436_ (.A(net58),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o211a_1 _3437_ (.A1(net340),
    .A2(_2798_),
    .B1(_2825_),
    .C1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_8 _3438_ (.A0(\as2650.r123[2][4] ),
    .A1(\as2650.r123_2[2][4] ),
    .S(net221),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_4 _3439_ (.A1(net253),
    .A2(net205),
    .B1(_0347_),
    .B2(net209),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_2 _3440_ (.A0(\as2650.r123[0][4] ),
    .A1(\as2650.r123_2[0][4] ),
    .S(net221),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _3441_ (.A0(\as2650.r123[1][4] ),
    .A1(\as2650.r123[0][4] ),
    .A2(\as2650.r123_2[1][4] ),
    .A3(\as2650.r123_2[0][4] ),
    .S0(net307),
    .S1(net221),
    .X(_0350_));
 sky130_fd_sc_hd__and3_4 _3442_ (.A(net207),
    .B(net203),
    .C(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_8 _3443_ (.A(_0348_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_4 _3444_ (.A(_0348_),
    .B(_0351_),
    .X(_0353_));
 sky130_fd_sc_hd__o21ai_1 _3445_ (.A1(_2825_),
    .A2(net110),
    .B1(net57),
    .Y(_0354_));
 sky130_fd_sc_hd__o22a_1 _3446_ (.A1(_2816_),
    .A2(net115),
    .B1(_0346_),
    .B2(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(_0355_),
    .A1(net255),
    .S(_2842_),
    .X(_0356_));
 sky130_fd_sc_hd__xnor2_2 _3448_ (.A(_2997_),
    .B(net111),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_1 _3449_ (.A(net114),
    .B(net112),
    .X(_0358_));
 sky130_fd_sc_hd__nor4_4 _3450_ (.A(_2880_),
    .B(net119),
    .C(net114),
    .D(net111),
    .Y(_0359_));
 sky130_fd_sc_hd__o31a_1 _3451_ (.A1(_2880_),
    .A2(net119),
    .A3(net115),
    .B1(net111),
    .X(_0360_));
 sky130_fd_sc_hd__or3_1 _3452_ (.A(_2904_),
    .B(_0359_),
    .C(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__o221a_4 _3453_ (.A1(_2905_),
    .A2(net111),
    .B1(_0357_),
    .B2(_2903_),
    .C1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__or3_1 _3454_ (.A(_2910_),
    .B(_0359_),
    .C(_0360_),
    .X(_0363_));
 sky130_fd_sc_hd__o221a_4 _3455_ (.A1(_2911_),
    .A2(net111),
    .B1(_0357_),
    .B2(_2909_),
    .C1(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _3456_ (.A(\as2650.holding_reg[3] ),
    .B(net112),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _3457_ (.A(\as2650.holding_reg[3] ),
    .B(net112),
    .Y(_0366_));
 sky130_fd_sc_hd__or2_1 _3458_ (.A(\as2650.holding_reg[3] ),
    .B(net112),
    .X(_0367_));
 sky130_fd_sc_hd__and2_4 _3459_ (.A(_0366_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(\as2650.holding_reg[2] ),
    .A1(net116),
    .S(net199),
    .X(_0369_));
 sky130_fd_sc_hd__o2bb2a_1 _3461_ (.A1_N(_0322_),
    .A2_N(_0323_),
    .B1(_0327_),
    .B2(_0320_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _3462_ (.A(_0368_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a21oi_1 _3463_ (.A1(_0368_),
    .A2(_0370_),
    .B1(_2930_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_1 _3464_ (.A(_0320_),
    .B(_0325_),
    .Y(_0373_));
 sky130_fd_sc_hd__nor2_1 _3465_ (.A(_0319_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__xnor2_1 _3466_ (.A(_0368_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__mux2_4 _3467_ (.A0(\as2650.holding_reg[3] ),
    .A1(net112),
    .S(net199),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(\as2650.holding_reg[3] ),
    .A1(net112),
    .S(net201),
    .X(_0377_));
 sky130_fd_sc_hd__a221o_1 _3469_ (.A1(_2754_),
    .A2(_0376_),
    .B1(_0377_),
    .B2(_2673_),
    .C1(_2756_),
    .X(_0378_));
 sky130_fd_sc_hd__a21o_1 _3470_ (.A1(_2925_),
    .A2(_0375_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__a21o_1 _3471_ (.A1(_0371_),
    .A2(_0372_),
    .B1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o211a_1 _3472_ (.A1(_2757_),
    .A2(_0365_),
    .B1(_0380_),
    .C1(_2915_),
    .X(_0381_));
 sky130_fd_sc_hd__a21oi_4 _3473_ (.A1(_2914_),
    .A2(_0368_),
    .B1(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(_0356_),
    .A1(_0362_),
    .S(_2839_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(_0364_),
    .A1(_0383_),
    .S(_2841_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _3476_ (.A(_2836_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__o21ai_4 _3477_ (.A1(_2836_),
    .A2(_0382_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a211o_1 _3478_ (.A1(_2833_),
    .A2(_0386_),
    .B1(_0342_),
    .C1(_2843_),
    .X(_0387_));
 sky130_fd_sc_hd__o21a_1 _3479_ (.A1(\as2650.r123[0][3] ),
    .A2(_2844_),
    .B1(_0387_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _3480_ (.A(net228),
    .B(\as2650.stack[3][12] ),
    .C(net195),
    .X(_0388_));
 sky130_fd_sc_hd__o22a_1 _3481_ (.A1(\as2650.stack[0][12] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[1][12] ),
    .X(_0389_));
 sky130_fd_sc_hd__o221a_1 _3482_ (.A1(\as2650.stack[2][12] ),
    .A2(net191),
    .B1(_0388_),
    .B2(_2849_),
    .C1(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__mux4_1 _3483_ (.A0(\as2650.stack[7][12] ),
    .A1(\as2650.stack[4][12] ),
    .A2(\as2650.stack[5][12] ),
    .A3(\as2650.stack[6][12] ),
    .S0(net224),
    .S1(net226),
    .X(_0391_));
 sky130_fd_sc_hd__a21o_2 _3484_ (.A1(net123),
    .A2(_0391_),
    .B1(_0390_),
    .X(_0392_));
 sky130_fd_sc_hd__o221a_1 _3485_ (.A1(net252),
    .A2(net75),
    .B1(_2846_),
    .B2(_0392_),
    .C1(_2868_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_4 _3486_ (.A0(\as2650.r123[2][5] ),
    .A1(\as2650.r123_2[2][5] ),
    .S(net220),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_4 _3487_ (.A1(net248),
    .A2(_2749_),
    .B1(_0394_),
    .B2(_2674_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_8 _3488_ (.A0(\as2650.r123[0][5] ),
    .A1(\as2650.r123_2[0][5] ),
    .S(net220),
    .X(_0396_));
 sky130_fd_sc_hd__mux4_1 _3489_ (.A0(\as2650.r123[1][5] ),
    .A1(\as2650.r123[0][5] ),
    .A2(\as2650.r123_2[1][5] ),
    .A3(\as2650.r123_2[0][5] ),
    .S0(net307),
    .S1(net220),
    .X(_0397_));
 sky130_fd_sc_hd__and3_4 _3490_ (.A(net207),
    .B(net203),
    .C(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_8 _3491_ (.A(_0395_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__or2_2 _3492_ (.A(_0395_),
    .B(_0398_),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_2 _3493_ (.A1(_2998_),
    .A2(net111),
    .B1(_0359_),
    .B2(_2945_),
    .X(_0401_));
 sky130_fd_sc_hd__xnor2_4 _3494_ (.A(net110),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__or2_1 _3495_ (.A(_2797_),
    .B(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _3496_ (.A1(_2655_),
    .A2(net58),
    .B1(_2824_),
    .Y(_0404_));
 sky130_fd_sc_hd__a22o_1 _3497_ (.A1(_2824_),
    .A2(net109),
    .B1(_0403_),
    .B2(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(net111),
    .A1(_0405_),
    .S(net57),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(_0406_),
    .A1(net253),
    .S(_2842_),
    .X(_0407_));
 sky130_fd_sc_hd__and4_2 _3500_ (.A(net114),
    .B(_2958_),
    .C(net113),
    .D(_0353_),
    .X(_0408_));
 sky130_fd_sc_hd__a31o_1 _3501_ (.A1(net115),
    .A2(_2958_),
    .A3(net112),
    .B1(_0353_),
    .X(_0409_));
 sky130_fd_sc_hd__nand2b_1 _3502_ (.A_N(_0408_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2b_1 _3503_ (.A_N(_2903_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_2 _3504_ (.A(net110),
    .B(_0359_),
    .Y(_0412_));
 sky130_fd_sc_hd__o221a_4 _3505_ (.A1(_2905_),
    .A2(_0353_),
    .B1(_0412_),
    .B2(_2904_),
    .C1(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(_0407_),
    .A1(_0413_),
    .S(_2839_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _3507_ (.A(_2908_),
    .B(_0410_),
    .Y(_0415_));
 sky130_fd_sc_hd__o221a_4 _3508_ (.A1(_2911_),
    .A2(_0353_),
    .B1(_0412_),
    .B2(_2910_),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_2 _3509_ (.A0(_2656_),
    .A1(net110),
    .S(net200),
    .X(_0417_));
 sky130_fd_sc_hd__inv_2 _3510_ (.A(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_2 _3511_ (.A(_2915_),
    .B(_0417_),
    .Y(_0419_));
 sky130_fd_sc_hd__nor2_4 _3512_ (.A(_2656_),
    .B(net110),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2_1 _3513_ (.A(\as2650.holding_reg[4] ),
    .B(_0353_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_4 _3514_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__o31a_2 _3515_ (.A1(_0319_),
    .A2(_0365_),
    .A3(_0373_),
    .B1(_0367_),
    .X(_0423_));
 sky130_fd_sc_hd__nand2_1 _3516_ (.A(_0422_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21a_1 _3517_ (.A1(_0422_),
    .A2(_0423_),
    .B1(_2925_),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _3518_ (.A(_0366_),
    .B(_0376_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21o_1 _3519_ (.A1(_0371_),
    .A2(_0426_),
    .B1(_0422_),
    .X(_0427_));
 sky130_fd_sc_hd__a31o_1 _3520_ (.A1(_0371_),
    .A2(_0422_),
    .A3(_0426_),
    .B1(_2930_),
    .X(_0428_));
 sky130_fd_sc_hd__and2b_1 _3521_ (.A_N(_0428_),
    .B(_0427_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(\as2650.holding_reg[4] ),
    .A1(_0353_),
    .S(net201),
    .X(_0430_));
 sky130_fd_sc_hd__a221o_1 _3523_ (.A1(_2754_),
    .A2(_0418_),
    .B1(_0430_),
    .B2(_2673_),
    .C1(_2756_),
    .X(_0431_));
 sky130_fd_sc_hd__a211o_1 _3524_ (.A1(_0424_),
    .A2(_0425_),
    .B1(_0429_),
    .C1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__o21ai_4 _3525_ (.A1(_2757_),
    .A2(_0420_),
    .B1(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__xnor2_4 _3526_ (.A(_0419_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__a21o_1 _3527_ (.A1(_2840_),
    .A2(_0416_),
    .B1(_2835_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _3528_ (.A1(_2841_),
    .A2(_0414_),
    .B1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__o21a_4 _3529_ (.A1(_2836_),
    .A2(_0434_),
    .B1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a211o_1 _3530_ (.A1(_2833_),
    .A2(_0437_),
    .B1(_0393_),
    .C1(_2843_),
    .X(_0438_));
 sky130_fd_sc_hd__o21a_1 _3531_ (.A1(\as2650.r123[0][4] ),
    .A2(_2844_),
    .B1(_0438_),
    .X(_0012_));
 sky130_fd_sc_hd__o22a_1 _3532_ (.A1(\as2650.stack[3][13] ),
    .A2(net194),
    .B1(net191),
    .B2(\as2650.stack[2][13] ),
    .X(_0439_));
 sky130_fd_sc_hd__o221a_1 _3533_ (.A1(\as2650.stack[0][13] ),
    .A2(net170),
    .B1(net166),
    .B2(\as2650.stack[1][13] ),
    .C1(_2859_),
    .X(_0440_));
 sky130_fd_sc_hd__o22a_1 _3534_ (.A1(\as2650.stack[7][13] ),
    .A2(net194),
    .B1(net192),
    .B2(\as2650.stack[6][13] ),
    .X(_0441_));
 sky130_fd_sc_hd__o221a_1 _3535_ (.A1(\as2650.stack[4][13] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[5][13] ),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_4 _3536_ (.A1(_0439_),
    .A2(_0440_),
    .B1(_0442_),
    .B2(net123),
    .X(_0443_));
 sky130_fd_sc_hd__o221a_1 _3537_ (.A1(net249),
    .A2(net75),
    .B1(_2846_),
    .B2(_0443_),
    .C1(_2868_),
    .X(_0444_));
 sky130_fd_sc_hd__and2_2 _3538_ (.A(net108),
    .B(_0408_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _3539_ (.A(net108),
    .B(_0408_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_1 _3540_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__or2_1 _3541_ (.A(_2909_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__and3_2 _3542_ (.A(net110),
    .B(_0359_),
    .C(_0399_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _3543_ (.A1(net110),
    .A2(_0359_),
    .B1(_0399_),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_2 _3544_ (.A(_0449_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__o221a_4 _3545_ (.A1(_2911_),
    .A2(net108),
    .B1(_0451_),
    .B2(_2910_),
    .C1(_0448_),
    .X(_0452_));
 sky130_fd_sc_hd__and3_1 _3546_ (.A(_2945_),
    .B(net110),
    .C(_0359_),
    .X(_0453_));
 sky130_fd_sc_hd__a21o_2 _3547_ (.A1(_2771_),
    .A2(_0408_),
    .B1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__xnor2_4 _3548_ (.A(net108),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _3549_ (.A(net336),
    .B(_2798_),
    .Y(_0456_));
 sky130_fd_sc_hd__a211o_1 _3550_ (.A1(_2798_),
    .A2(_0455_),
    .B1(_0456_),
    .C1(_2824_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_4 _3551_ (.A0(\as2650.r123[2][6] ),
    .A1(\as2650.r123_2[2][6] ),
    .S(net221),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_4 _3552_ (.A1(net245),
    .A2(_2749_),
    .B1(_0458_),
    .B2(_2674_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_2 _3553_ (.A0(\as2650.r123[0][6] ),
    .A1(\as2650.r123_2[0][6] ),
    .S(net220),
    .X(_0460_));
 sky130_fd_sc_hd__mux4_1 _3554_ (.A0(\as2650.r123[1][6] ),
    .A1(\as2650.r123[0][6] ),
    .A2(\as2650.r123_2[1][6] ),
    .A3(\as2650.r123_2[0][6] ),
    .S0(net307),
    .S1(net222),
    .X(_0461_));
 sky130_fd_sc_hd__and3_4 _3555_ (.A(net207),
    .B(net203),
    .C(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_8 _3556_ (.A(_0459_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__or2_4 _3557_ (.A(_0459_),
    .B(_0462_),
    .X(_0464_));
 sky130_fd_sc_hd__o211a_1 _3558_ (.A1(_2825_),
    .A2(_0463_),
    .B1(_0457_),
    .C1(net57),
    .X(_0465_));
 sky130_fd_sc_hd__a21oi_1 _3559_ (.A1(_2777_),
    .A2(_0352_),
    .B1(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(_0466_),
    .A1(net248),
    .S(_2842_),
    .X(_0467_));
 sky130_fd_sc_hd__or2_1 _3561_ (.A(_2903_),
    .B(_0447_),
    .X(_0468_));
 sky130_fd_sc_hd__o221a_4 _3562_ (.A1(_2905_),
    .A2(net108),
    .B1(_0451_),
    .B2(_2904_),
    .C1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(_0467_),
    .A1(_0469_),
    .S(_2839_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(_0452_),
    .A1(_0470_),
    .S(_2841_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_2 _3565_ (.A(\as2650.holding_reg[5] ),
    .B(net108),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _3566_ (.A(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_2 _3567_ (.A(\as2650.holding_reg[5] ),
    .B(net108),
    .Y(_0474_));
 sky130_fd_sc_hd__nor2_4 _3568_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__a21oi_2 _3569_ (.A1(_0422_),
    .A2(_0423_),
    .B1(_0420_),
    .Y(_0476_));
 sky130_fd_sc_hd__xor2_1 _3570_ (.A(_0475_),
    .B(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__or2_1 _3571_ (.A(_0417_),
    .B(_0420_),
    .X(_0478_));
 sky130_fd_sc_hd__and3_1 _3572_ (.A(_0427_),
    .B(_0475_),
    .C(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__a21o_1 _3573_ (.A1(_0427_),
    .A2(_0478_),
    .B1(_0475_),
    .X(_0480_));
 sky130_fd_sc_hd__or3b_1 _3574_ (.A(_2930_),
    .B(_0479_),
    .C_N(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__or2_1 _3575_ (.A(\as2650.holding_reg[5] ),
    .B(net199),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_1 _3576_ (.A1(net201),
    .A2(net108),
    .B1(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o21ai_1 _3577_ (.A1(net201),
    .A2(net108),
    .B1(_0482_),
    .Y(_0484_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\as2650.holding_reg[5] ),
    .A1(net108),
    .S(net201),
    .X(_0485_));
 sky130_fd_sc_hd__a221oi_2 _3579_ (.A1(_2754_),
    .A2(_0483_),
    .B1(_0485_),
    .B2(_2673_),
    .C1(_2756_),
    .Y(_0486_));
 sky130_fd_sc_hd__o211a_1 _3580_ (.A1(_2926_),
    .A2(_0477_),
    .B1(_0481_),
    .C1(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a21o_1 _3581_ (.A1(_2756_),
    .A2(_0472_),
    .B1(_2914_),
    .X(_0488_));
 sky130_fd_sc_hd__a2bb2o_4 _3582_ (.A1_N(_0487_),
    .A2_N(_0488_),
    .B1(_2914_),
    .B2(_0475_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_4 _3583_ (.A0(_0471_),
    .A1(_0489_),
    .S(_2835_),
    .X(_0490_));
 sky130_fd_sc_hd__a211o_1 _3584_ (.A1(_2833_),
    .A2(_0490_),
    .B1(_0444_),
    .C1(_2843_),
    .X(_0491_));
 sky130_fd_sc_hd__o21a_1 _3585_ (.A1(\as2650.r123[0][5] ),
    .A2(_2844_),
    .B1(_0491_),
    .X(_0013_));
 sky130_fd_sc_hd__o22a_1 _3586_ (.A1(\as2650.stack[7][14] ),
    .A2(net194),
    .B1(net191),
    .B2(\as2650.stack[6][14] ),
    .X(_0492_));
 sky130_fd_sc_hd__o221a_1 _3587_ (.A1(\as2650.stack[4][14] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[5][14] ),
    .C1(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__o22a_1 _3588_ (.A1(\as2650.stack[3][14] ),
    .A2(net194),
    .B1(net191),
    .B2(\as2650.stack[2][14] ),
    .X(_0494_));
 sky130_fd_sc_hd__o221a_1 _3589_ (.A1(\as2650.stack[0][14] ),
    .A2(net169),
    .B1(net165),
    .B2(\as2650.stack[1][14] ),
    .C1(_2859_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_4 _3590_ (.A1(net123),
    .A2(_0493_),
    .B1(_0494_),
    .B2(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__o221a_1 _3591_ (.A1(net244),
    .A2(net75),
    .B1(_2846_),
    .B2(_0496_),
    .C1(_2868_),
    .X(_0497_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(_2843_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__and3_2 _3593_ (.A(net109),
    .B(_0408_),
    .C(net107),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_1 _3594_ (.A(_0445_),
    .B(net107),
    .Y(_0500_));
 sky130_fd_sc_hd__a21oi_1 _3595_ (.A1(_2771_),
    .A2(_0445_),
    .B1(net107),
    .Y(_0501_));
 sky130_fd_sc_hd__a22o_1 _3596_ (.A1(_2945_),
    .A2(_0449_),
    .B1(_0499_),
    .B2(_2771_),
    .X(_0502_));
 sky130_fd_sc_hd__and3_1 _3597_ (.A(net110),
    .B(_0399_),
    .C(_0463_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_2 _3598_ (.A(_0359_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__and3_1 _3599_ (.A(_2945_),
    .B(_0359_),
    .C(_0503_),
    .X(_0505_));
 sky130_fd_sc_hd__o21ba_2 _3600_ (.A1(_0501_),
    .A2(_0502_),
    .B1_N(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_1 _3601_ (.A(net58),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__a211o_1 _3602_ (.A1(net334),
    .A2(_2797_),
    .B1(_2824_),
    .C1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__o211a_1 _3603_ (.A1(_2825_),
    .A2(_2897_),
    .B1(_0508_),
    .C1(net57),
    .X(_0509_));
 sky130_fd_sc_hd__a211o_1 _3604_ (.A1(_2838_),
    .A2(net109),
    .B1(_0509_),
    .C1(_2842_),
    .X(_0510_));
 sky130_fd_sc_hd__o211a_1 _3605_ (.A1(net245),
    .A2(_2818_),
    .B1(_2821_),
    .C1(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__nor2_2 _3606_ (.A(_0499_),
    .B(_0500_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_1 _3607_ (.A(_0449_),
    .B(_0463_),
    .Y(_0513_));
 sky130_fd_sc_hd__or2_1 _3608_ (.A(_2904_),
    .B(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__o221a_4 _3609_ (.A1(_2905_),
    .A2(net106),
    .B1(_0512_),
    .B2(_2903_),
    .C1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__a211o_2 _3610_ (.A1(_2839_),
    .A2(_0515_),
    .B1(_0511_),
    .C1(_2840_),
    .X(_0516_));
 sky130_fd_sc_hd__or2_1 _3611_ (.A(_2910_),
    .B(_0513_),
    .X(_0517_));
 sky130_fd_sc_hd__o221a_4 _3612_ (.A1(_2911_),
    .A2(net107),
    .B1(_0512_),
    .B2(_2909_),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__o211ai_4 _3613_ (.A1(_2841_),
    .A2(_0518_),
    .B1(_0516_),
    .C1(_2836_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_2 _3614_ (.A(\as2650.holding_reg[6] ),
    .B(net106),
    .Y(_0520_));
 sky130_fd_sc_hd__or2_1 _3615_ (.A(\as2650.holding_reg[6] ),
    .B(net106),
    .X(_0521_));
 sky130_fd_sc_hd__and2_1 _3616_ (.A(_0520_),
    .B(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nand2_2 _3617_ (.A(_0520_),
    .B(_0521_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_0472_),
    .B(_0483_),
    .Y(_0524_));
 sky130_fd_sc_hd__and3_1 _3619_ (.A(_0480_),
    .B(_0522_),
    .C(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__a21oi_2 _3620_ (.A1(_0480_),
    .A2(_0524_),
    .B1(_0522_),
    .Y(_0526_));
 sky130_fd_sc_hd__or3_1 _3621_ (.A(_2930_),
    .B(_0525_),
    .C(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__o21ai_2 _3622_ (.A1(_0474_),
    .A2(_0476_),
    .B1(_0472_),
    .Y(_0528_));
 sky130_fd_sc_hd__xnor2_1 _3623_ (.A(_0523_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__mux2_2 _3624_ (.A0(\as2650.holding_reg[6] ),
    .A1(net106),
    .S(net198),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _3625_ (.A0(\as2650.holding_reg[6] ),
    .A1(net106),
    .S(net201),
    .X(_0531_));
 sky130_fd_sc_hd__a221o_1 _3626_ (.A1(_2754_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_2673_),
    .C1(_2756_),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _3627_ (.A1(_2925_),
    .A2(_0529_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(_2756_),
    .A2(_0520_),
    .B1(_0527_),
    .B2(_0533_),
    .C1(_2914_),
    .X(_0534_));
 sky130_fd_sc_hd__o21a_4 _3629_ (.A1(_2915_),
    .A2(_0523_),
    .B1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o21ai_4 _3630_ (.A1(_2836_),
    .A2(_0535_),
    .B1(_0519_),
    .Y(_0536_));
 sky130_fd_sc_hd__and2_1 _3631_ (.A(_2833_),
    .B(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__o22a_1 _3632_ (.A1(\as2650.r123[0][6] ),
    .A2(_2844_),
    .B1(_0498_),
    .B2(_0537_),
    .X(_0014_));
 sky130_fd_sc_hd__a31o_1 _3633_ (.A1(net241),
    .A2(net74),
    .A3(_2868_),
    .B1(_2843_),
    .X(_0538_));
 sky130_fd_sc_hd__a31o_2 _3634_ (.A1(_2771_),
    .A2(_0445_),
    .A3(net107),
    .B1(_0505_),
    .X(_0539_));
 sky130_fd_sc_hd__xnor2_4 _3635_ (.A(net118),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nor2_1 _3636_ (.A(net58),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__a211o_1 _3637_ (.A1(net331),
    .A2(net58),
    .B1(_2824_),
    .C1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__o21a_2 _3638_ (.A1(\as2650.psl[3] ),
    .A2(net121),
    .B1(_2890_),
    .X(_0543_));
 sky130_fd_sc_hd__o211a_1 _3639_ (.A1(_2825_),
    .A2(_0543_),
    .B1(_0542_),
    .C1(net57),
    .X(_0544_));
 sky130_fd_sc_hd__a211o_1 _3640_ (.A1(_2777_),
    .A2(net107),
    .B1(_0544_),
    .C1(_2842_),
    .X(_0545_));
 sky130_fd_sc_hd__o21a_1 _3641_ (.A1(net241),
    .A2(_2818_),
    .B1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__xnor2_2 _3642_ (.A(_2896_),
    .B(_0499_),
    .Y(_0547_));
 sky130_fd_sc_hd__xnor2_2 _3643_ (.A(_2897_),
    .B(_0504_),
    .Y(_0548_));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(net118),
    .B(_2905_),
    .X(_0549_));
 sky130_fd_sc_hd__o221a_4 _3645_ (.A1(_2903_),
    .A2(_0547_),
    .B1(_0548_),
    .B2(_2904_),
    .C1(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or2_1 _3646_ (.A(net118),
    .B(_2911_),
    .X(_0551_));
 sky130_fd_sc_hd__o221a_4 _3647_ (.A1(_2909_),
    .A2(_0547_),
    .B1(_0548_),
    .B2(_2910_),
    .C1(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(\as2650.holding_reg[7] ),
    .B(net118),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_2 _3649_ (.A(_2659_),
    .B(_2896_),
    .Y(_0554_));
 sky130_fd_sc_hd__and2_2 _3650_ (.A(_0553_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_2 _3651_ (.A(_0553_),
    .B(_0554_),
    .Y(_0556_));
 sky130_fd_sc_hd__and2_1 _3652_ (.A(_0520_),
    .B(_0530_),
    .X(_0557_));
 sky130_fd_sc_hd__or3_1 _3653_ (.A(_0526_),
    .B(_0555_),
    .C(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o21ai_1 _3654_ (.A1(_0526_),
    .A2(_0557_),
    .B1(_0555_),
    .Y(_0559_));
 sky130_fd_sc_hd__a21o_1 _3655_ (.A1(_0558_),
    .A2(_0559_),
    .B1(_2930_),
    .X(_0560_));
 sky130_fd_sc_hd__a21boi_1 _3656_ (.A1(_0522_),
    .A2(_0528_),
    .B1_N(_0520_),
    .Y(_0561_));
 sky130_fd_sc_hd__xnor2_1 _3657_ (.A(_0556_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(_2659_),
    .A1(_2896_),
    .S(net201),
    .X(_0563_));
 sky130_fd_sc_hd__o221a_1 _3659_ (.A1(_2926_),
    .A2(_0562_),
    .B1(_0563_),
    .B2(_2672_),
    .C1(_2977_),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _3660_ (.A1(net300),
    .A2(_0554_),
    .B1(_2755_),
    .Y(_0565_));
 sky130_fd_sc_hd__a21oi_1 _3661_ (.A1(_0560_),
    .A2(_0564_),
    .B1(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__a31o_1 _3662_ (.A1(\as2650.holding_reg[7] ),
    .A2(_2756_),
    .A3(net118),
    .B1(_2914_),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_4 _3663_ (.A1(_2915_),
    .A2(_0555_),
    .B1(_0566_),
    .B2(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__o221a_1 _3664_ (.A1(_2839_),
    .A2(_0546_),
    .B1(_0550_),
    .B2(_2821_),
    .C1(_2822_),
    .X(_0569_));
 sky130_fd_sc_hd__a211o_1 _3665_ (.A1(_2840_),
    .A2(_0552_),
    .B1(_0569_),
    .C1(_2835_),
    .X(_0570_));
 sky130_fd_sc_hd__o21a_4 _3666_ (.A1(_2836_),
    .A2(_0568_),
    .B1(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _3667_ (.A1(_2833_),
    .A2(_0571_),
    .B1(_0538_),
    .X(_0572_));
 sky130_fd_sc_hd__o21a_1 _3668_ (.A1(\as2650.r123[0][7] ),
    .A2(_2844_),
    .B1(_0572_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_4 _3669_ (.A(net217),
    .B(_2687_),
    .Y(_0573_));
 sky130_fd_sc_hd__nor2_8 _3670_ (.A(net309),
    .B(net149),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_4 _3671_ (.A(_2648_),
    .B(net153),
    .Y(_0575_));
 sky130_fd_sc_hd__nor2_2 _3672_ (.A(net148),
    .B(_0573_),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_1 _3673_ (.A(_0573_),
    .B(_0574_),
    .Y(_0577_));
 sky130_fd_sc_hd__o22a_1 _3674_ (.A1(net328),
    .A2(net77),
    .B1(_0577_),
    .B2(net101),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_4 _3675_ (.A(net215),
    .B(net146),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_2 _3676_ (.A(net237),
    .B(net145),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2b_2 _3677_ (.A_N(_2788_),
    .B(_2763_),
    .Y(_0581_));
 sky130_fd_sc_hd__or3_1 _3678_ (.A(_0578_),
    .B(_0580_),
    .C(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or3_1 _3679_ (.A(_2647_),
    .B(net98),
    .C(net149),
    .X(_0583_));
 sky130_fd_sc_hd__a21o_4 _3680_ (.A1(_0582_),
    .A2(_0583_),
    .B1(net206),
    .X(_0584_));
 sky130_fd_sc_hd__or3_4 _3681_ (.A(net219),
    .B(net170),
    .C(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__nor3_4 _3682_ (.A(net198),
    .B(_2806_),
    .C(_2810_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_8 _3683_ (.A(net93),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_2 _3684_ (.A(_2745_),
    .B(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__or3_4 _3685_ (.A(net219),
    .B(net166),
    .C(net55),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _3686_ (.A0(net288),
    .A1(\as2650.stack[5][0] ),
    .S(_0585_),
    .X(_0590_));
 sky130_fd_sc_hd__nand2_4 _3687_ (.A(net139),
    .B(_0586_),
    .Y(_0591_));
 sky130_fd_sc_hd__mux2_1 _3688_ (.A0(net265),
    .A1(_0590_),
    .S(_0589_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(net285),
    .A1(\as2650.stack[5][1] ),
    .S(_0585_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(net261),
    .A1(_0592_),
    .S(_0589_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(\as2650.pc[2] ),
    .A1(\as2650.stack[5][2] ),
    .S(_0585_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(net257),
    .A1(_0593_),
    .S(_0589_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(net283),
    .A1(\as2650.stack[5][3] ),
    .S(_0585_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(net254),
    .A1(_0594_),
    .S(_0589_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _3695_ (.A0(net281),
    .A1(\as2650.stack[5][4] ),
    .S(_0585_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _3696_ (.A0(net251),
    .A1(_0595_),
    .S(_0589_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(net280),
    .A1(\as2650.stack[5][5] ),
    .S(_0585_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _3698_ (.A0(net247),
    .A1(_0596_),
    .S(_0589_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _3699_ (.A0(net277),
    .A1(\as2650.stack[5][6] ),
    .S(_0585_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _3700_ (.A0(net243),
    .A1(_0597_),
    .S(_0589_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(net275),
    .A1(\as2650.stack[5][7] ),
    .S(_0585_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(net239),
    .A1(_0598_),
    .S(_0589_),
    .X(_0023_));
 sky130_fd_sc_hd__nor3_4 _3703_ (.A(_2627_),
    .B(net166),
    .C(net49),
    .Y(_0599_));
 sky130_fd_sc_hd__or3_4 _3704_ (.A(net219),
    .B(net166),
    .C(net49),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_8 _3705_ (.A(_0589_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_8 _3706_ (.A(_2802_),
    .B(_0587_),
    .Y(_0602_));
 sky130_fd_sc_hd__or2_4 _3707_ (.A(_2624_),
    .B(net206),
    .X(_0603_));
 sky130_fd_sc_hd__nor3_4 _3708_ (.A(_2624_),
    .B(_2745_),
    .C(_0591_),
    .Y(_0604_));
 sky130_fd_sc_hd__mux2_8 _3709_ (.A0(\as2650.r123[0][0] ),
    .A1(\as2650.r123_2[0][0] ),
    .S(net220),
    .X(_0605_));
 sky130_fd_sc_hd__o22a_1 _3710_ (.A1(net274),
    .A2(_0604_),
    .B1(_0605_),
    .B2(net55),
    .X(_0606_));
 sky130_fd_sc_hd__a21o_4 _3711_ (.A1(\as2650.r123[0][0] ),
    .A2(_0602_),
    .B1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _3712_ (.A0(\as2650.stack[6][8] ),
    .A1(_0607_),
    .S(_0601_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_8 _3713_ (.A0(\as2650.r123[0][1] ),
    .A1(\as2650.r123_2[0][1] ),
    .S(net222),
    .X(_0608_));
 sky130_fd_sc_hd__o22a_1 _3714_ (.A1(net273),
    .A2(_0604_),
    .B1(_0608_),
    .B2(net55),
    .X(_0609_));
 sky130_fd_sc_hd__a21o_4 _3715_ (.A1(\as2650.r123[0][1] ),
    .A2(_0602_),
    .B1(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _3716_ (.A0(\as2650.stack[6][9] ),
    .A1(_0610_),
    .S(_0601_),
    .X(_0025_));
 sky130_fd_sc_hd__o22a_1 _3717_ (.A1(net187),
    .A2(net55),
    .B1(_0604_),
    .B2(net272),
    .X(_0611_));
 sky130_fd_sc_hd__a21o_4 _3718_ (.A1(\as2650.r123[0][2] ),
    .A2(_0602_),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(\as2650.stack[6][10] ),
    .A1(_0612_),
    .S(_0601_),
    .X(_0026_));
 sky130_fd_sc_hd__o22a_1 _3720_ (.A1(net185),
    .A2(net55),
    .B1(_0604_),
    .B2(\as2650.pc[11] ),
    .X(_0613_));
 sky130_fd_sc_hd__a21o_4 _3721_ (.A1(\as2650.r123[0][3] ),
    .A2(_0602_),
    .B1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _3722_ (.A0(\as2650.stack[6][11] ),
    .A1(_0614_),
    .S(_0601_),
    .X(_0027_));
 sky130_fd_sc_hd__o22a_1 _3723_ (.A1(net183),
    .A2(net56),
    .B1(_0604_),
    .B2(net269),
    .X(_0615_));
 sky130_fd_sc_hd__a21o_4 _3724_ (.A1(\as2650.r123[0][4] ),
    .A2(_0602_),
    .B1(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _3725_ (.A0(\as2650.stack[6][12] ),
    .A1(_0616_),
    .S(_0601_),
    .X(_0028_));
 sky130_fd_sc_hd__o22a_1 _3726_ (.A1(_0396_),
    .A2(_0588_),
    .B1(_0604_),
    .B2(\as2650.pc[13] ),
    .X(_0617_));
 sky130_fd_sc_hd__a21o_4 _3727_ (.A1(\as2650.r123[0][5] ),
    .A2(_0602_),
    .B1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(\as2650.stack[6][13] ),
    .A1(_0618_),
    .S(_0601_),
    .X(_0029_));
 sky130_fd_sc_hd__o22a_1 _3729_ (.A1(net179),
    .A2(_0588_),
    .B1(_0604_),
    .B2(\as2650.pc[14] ),
    .X(_0619_));
 sky130_fd_sc_hd__a21o_4 _3730_ (.A1(\as2650.r123[0][6] ),
    .A2(_0602_),
    .B1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(\as2650.stack[6][14] ),
    .A1(_0620_),
    .S(_0601_),
    .X(_0030_));
 sky130_fd_sc_hd__nor2_1 _3732_ (.A(_2624_),
    .B(net90),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _3733_ (.A(_2745_),
    .B(_2871_),
    .Y(_0622_));
 sky130_fd_sc_hd__or2_4 _3734_ (.A(_2745_),
    .B(_2871_),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _3735_ (.A(_2796_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__or2_2 _3736_ (.A(_2796_),
    .B(_0623_),
    .X(_0625_));
 sky130_fd_sc_hd__nor2_2 _3737_ (.A(_2762_),
    .B(_0623_),
    .Y(_0626_));
 sky130_fd_sc_hd__or2_4 _3738_ (.A(_2762_),
    .B(_0623_),
    .X(_0627_));
 sky130_fd_sc_hd__or3_4 _3739_ (.A(net127),
    .B(_2815_),
    .C(_0623_),
    .X(_0628_));
 sky130_fd_sc_hd__and4_4 _3740_ (.A(net86),
    .B(_2778_),
    .C(_2819_),
    .D(_2870_),
    .X(_0629_));
 sky130_fd_sc_hd__or4_4 _3741_ (.A(net83),
    .B(_2779_),
    .C(_2820_),
    .D(_2871_),
    .X(_0630_));
 sky130_fd_sc_hd__or4_2 _3742_ (.A(net237),
    .B(net134),
    .C(net128),
    .D(_0623_),
    .X(_0631_));
 sky130_fd_sc_hd__and3_4 _3743_ (.A(net139),
    .B(_2767_),
    .C(_0622_),
    .X(_0632_));
 sky130_fd_sc_hd__or3_4 _3744_ (.A(net134),
    .B(_2768_),
    .C(_0623_),
    .X(_0633_));
 sky130_fd_sc_hd__and3_4 _3745_ (.A(net139),
    .B(_2775_),
    .C(_0622_),
    .X(_0634_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__or2_4 _3747_ (.A(_2834_),
    .B(_0603_),
    .X(_0636_));
 sky130_fd_sc_hd__clkinv_2 _3748_ (.A(net60),
    .Y(_0637_));
 sky130_fd_sc_hd__and3_4 _3749_ (.A(_2782_),
    .B(_2786_),
    .C(_2870_),
    .X(_0638_));
 sky130_fd_sc_hd__or3_4 _3750_ (.A(_2783_),
    .B(_2787_),
    .C(_2871_),
    .X(_0639_));
 sky130_fd_sc_hd__and4_1 _3751_ (.A(_0630_),
    .B(_0635_),
    .C(net60),
    .D(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__o311a_1 _3752_ (.A1(_2769_),
    .A2(_2827_),
    .A3(_0623_),
    .B1(_0625_),
    .C1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_2 _3753_ (.A(_0631_),
    .B(_0633_),
    .C(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_4 _3754_ (.A(\as2650.ins_reg[1] ),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_1 _3755_ (.A(_2881_),
    .B(net54),
    .Y(_0644_));
 sky130_fd_sc_hd__a211o_1 _3756_ (.A1(net347),
    .A2(net54),
    .B1(_0626_),
    .C1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__o211a_1 _3757_ (.A1(net119),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__a211o_1 _3758_ (.A1(_2899_),
    .A2(_0634_),
    .B1(_0646_),
    .C1(_0632_),
    .X(_0647_));
 sky130_fd_sc_hd__o211a_1 _3759_ (.A1(net266),
    .A2(_0633_),
    .B1(_0647_),
    .C1(_0630_),
    .X(_0648_));
 sky130_fd_sc_hd__a211o_1 _3760_ (.A1(_2906_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__o21ai_1 _3761_ (.A1(_2912_),
    .A2(_0639_),
    .B1(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(_2934_),
    .B(net60),
    .Y(_0651_));
 sky130_fd_sc_hd__a21o_2 _3763_ (.A1(_0636_),
    .A2(_0650_),
    .B1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__nor2_1 _3764_ (.A(_0643_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__or3_4 _3765_ (.A(net135),
    .B(net74),
    .C(_0603_),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_2 _3766_ (.A(net223),
    .B(net139),
    .Y(_0655_));
 sky130_fd_sc_hd__a31o_1 _3767_ (.A1(_2636_),
    .A2(_2813_),
    .A3(_0621_),
    .B1(net325),
    .X(_0656_));
 sky130_fd_sc_hd__inv_2 _3768_ (.A(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__and4_1 _3769_ (.A(_2636_),
    .B(net318),
    .C(_2813_),
    .D(_0621_),
    .X(_0658_));
 sky130_fd_sc_hd__o221a_1 _3770_ (.A1(net267),
    .A2(net76),
    .B1(_2863_),
    .B2(_0654_),
    .C1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__and2_4 _3771_ (.A(_0643_),
    .B(_0657_),
    .X(_0660_));
 sky130_fd_sc_hd__and4b_4 _3772_ (.A_N(_0655_),
    .B(_2813_),
    .C(net318),
    .D(net218),
    .X(_0661_));
 sky130_fd_sc_hd__a211o_1 _3773_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_0660_),
    .B1(_0659_),
    .C1(_0653_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _3774_ (.A0(net346),
    .A1(_2947_),
    .S(_0625_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(net117),
    .A1(_0662_),
    .S(_0631_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _3776_ (.A0(_2880_),
    .A1(_0663_),
    .S(_0635_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(net263),
    .A1(_0664_),
    .S(_0633_),
    .X(_0665_));
 sky130_fd_sc_hd__a21o_1 _3778_ (.A1(_2962_),
    .A2(_0629_),
    .B1(_0638_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _3779_ (.A1(_0630_),
    .A2(_0665_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__o21a_1 _3780_ (.A1(_2965_),
    .A2(_0639_),
    .B1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or2_2 _3781_ (.A(_2986_),
    .B(net60),
    .X(_0669_));
 sky130_fd_sc_hd__o21ai_4 _3782_ (.A1(_0637_),
    .A2(_0668_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _3783_ (.A(_0643_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__o221a_1 _3784_ (.A1(net263),
    .A2(net76),
    .B1(_2943_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0672_));
 sky130_fd_sc_hd__a211o_1 _3785_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_0660_),
    .B1(_0671_),
    .C1(_0672_),
    .X(_0032_));
 sky130_fd_sc_hd__nor2_1 _3786_ (.A(_3000_),
    .B(net54),
    .Y(_0673_));
 sky130_fd_sc_hd__a211o_1 _3787_ (.A1(net344),
    .A2(net54),
    .B1(_0626_),
    .C1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__o211a_1 _3788_ (.A1(net111),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_1 _3789_ (.A1(net119),
    .A2(_0634_),
    .B1(_0675_),
    .C1(_0632_),
    .X(_0676_));
 sky130_fd_sc_hd__o211a_1 _3790_ (.A1(net258),
    .A2(_0633_),
    .B1(_0676_),
    .C1(_0630_),
    .X(_0677_));
 sky130_fd_sc_hd__a211o_1 _3791_ (.A1(_0312_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__o21ai_1 _3792_ (.A1(_0316_),
    .A2(_0639_),
    .B1(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nor2_1 _3793_ (.A(_0333_),
    .B(_0636_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21o_2 _3794_ (.A1(_0636_),
    .A2(_0679_),
    .B1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__nor2_1 _3795_ (.A(_0643_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o221a_1 _3796_ (.A1(net259),
    .A2(net75),
    .B1(_2993_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0683_));
 sky130_fd_sc_hd__a211o_1 _3797_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_0660_),
    .B1(_0682_),
    .C1(_0683_),
    .X(_0033_));
 sky130_fd_sc_hd__nor2_1 _3798_ (.A(_0344_),
    .B(net54),
    .Y(_0684_));
 sky130_fd_sc_hd__a211o_1 _3799_ (.A1(_2654_),
    .A2(net54),
    .B1(_0626_),
    .C1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o211a_1 _3800_ (.A1(_0352_),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_1 _3801_ (.A(net115),
    .B(_0628_),
    .Y(_0687_));
 sky130_fd_sc_hd__o21ai_1 _3802_ (.A1(_0686_),
    .A2(_0687_),
    .B1(_0633_),
    .Y(_0688_));
 sky130_fd_sc_hd__o211a_1 _3803_ (.A1(net255),
    .A2(_0633_),
    .B1(_0688_),
    .C1(_0630_),
    .X(_0689_));
 sky130_fd_sc_hd__a211o_1 _3804_ (.A1(_0362_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__o21ai_1 _3805_ (.A1(_0364_),
    .A2(_0639_),
    .B1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__mux2_4 _3806_ (.A0(_0382_),
    .A1(_0691_),
    .S(net60),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_1 _3807_ (.A(_0643_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__o221a_1 _3808_ (.A1(net256),
    .A2(net75),
    .B1(_0341_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0694_));
 sky130_fd_sc_hd__a211o_1 _3809_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_0660_),
    .B1(_0693_),
    .C1(_0694_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(net339),
    .A1(_0402_),
    .S(_0625_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(net109),
    .A1(_0695_),
    .S(_0631_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _3812_ (.A0(net111),
    .A1(_0696_),
    .S(_0635_),
    .X(_0697_));
 sky130_fd_sc_hd__or2_1 _3813_ (.A(_0632_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__o211a_1 _3814_ (.A1(net253),
    .A2(_0633_),
    .B1(_0698_),
    .C1(_0630_),
    .X(_0699_));
 sky130_fd_sc_hd__a211o_1 _3815_ (.A1(_0413_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _3816_ (.A(_0416_),
    .B(_0639_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _3817_ (.A1(_0700_),
    .A2(_0701_),
    .B1(_0637_),
    .X(_0702_));
 sky130_fd_sc_hd__o21ai_4 _3818_ (.A1(_0434_),
    .A2(net60),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _3819_ (.A(_0643_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__o221a_1 _3820_ (.A1(net252),
    .A2(net75),
    .B1(_0392_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0705_));
 sky130_fd_sc_hd__a211o_1 _3821_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_0660_),
    .B1(_0704_),
    .C1(_0705_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _3822_ (.A(_0455_),
    .B(net54),
    .Y(_0706_));
 sky130_fd_sc_hd__a211o_1 _3823_ (.A1(net336),
    .A2(net54),
    .B1(_0626_),
    .C1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__o211a_1 _3824_ (.A1(net107),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__a211o_1 _3825_ (.A1(_0353_),
    .A2(_0634_),
    .B1(_0708_),
    .C1(_0632_),
    .X(_0709_));
 sky130_fd_sc_hd__o211a_1 _3826_ (.A1(net248),
    .A2(_0633_),
    .B1(_0709_),
    .C1(_0630_),
    .X(_0710_));
 sky130_fd_sc_hd__a211o_1 _3827_ (.A1(_0469_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__o21ai_1 _3828_ (.A1(_0452_),
    .A2(_0639_),
    .B1(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2_1 _3829_ (.A(_0489_),
    .B(net60),
    .Y(_0713_));
 sky130_fd_sc_hd__a21o_2 _3830_ (.A1(net60),
    .A2(_0712_),
    .B1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _3831_ (.A(_0643_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__o221a_1 _3832_ (.A1(net248),
    .A2(net75),
    .B1(_0443_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0716_));
 sky130_fd_sc_hd__a211o_1 _3833_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_0660_),
    .B1(_0715_),
    .C1(_0716_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_1 _3834_ (.A(_0506_),
    .B(_0624_),
    .Y(_0717_));
 sky130_fd_sc_hd__a211o_1 _3835_ (.A1(net334),
    .A2(_0624_),
    .B1(_0626_),
    .C1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__o211a_1 _3836_ (.A1(_2897_),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__a211o_1 _3837_ (.A1(net109),
    .A2(_0634_),
    .B1(_0719_),
    .C1(_0632_),
    .X(_0720_));
 sky130_fd_sc_hd__o211a_1 _3838_ (.A1(net245),
    .A2(_0633_),
    .B1(_0720_),
    .C1(_0630_),
    .X(_0721_));
 sky130_fd_sc_hd__a211o_1 _3839_ (.A1(_0515_),
    .A2(_0629_),
    .B1(_0638_),
    .C1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__o21ai_1 _3840_ (.A1(_0518_),
    .A2(_0639_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__mux2_4 _3841_ (.A0(_0535_),
    .A1(_0723_),
    .S(net60),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(_0643_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o221a_1 _3843_ (.A1(net245),
    .A2(net76),
    .B1(_0496_),
    .B2(_0654_),
    .C1(_0661_),
    .X(_0726_));
 sky130_fd_sc_hd__a211o_1 _3844_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_0660_),
    .B1(_0725_),
    .C1(_0726_),
    .X(_0037_));
 sky130_fd_sc_hd__nor2_1 _3845_ (.A(_0540_),
    .B(net54),
    .Y(_0727_));
 sky130_fd_sc_hd__a211o_1 _3846_ (.A1(net331),
    .A2(net54),
    .B1(_0626_),
    .C1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__o211a_1 _3847_ (.A1(_0543_),
    .A2(_0627_),
    .B1(_0628_),
    .C1(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__a211o_1 _3848_ (.A1(net107),
    .A2(_0634_),
    .B1(_0729_),
    .C1(_0632_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(_2628_),
    .B(_0632_),
    .Y(_0731_));
 sky130_fd_sc_hd__a21o_1 _3850_ (.A1(_0730_),
    .A2(_0731_),
    .B1(_0629_),
    .X(_0732_));
 sky130_fd_sc_hd__o211a_1 _3851_ (.A1(_0550_),
    .A2(_0630_),
    .B1(_0639_),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__a211o_1 _3852_ (.A1(_0552_),
    .A2(_0638_),
    .B1(_0733_),
    .C1(_0637_),
    .X(_0734_));
 sky130_fd_sc_hd__o21a_2 _3853_ (.A1(_0568_),
    .A2(net60),
    .B1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__a32o_1 _3854_ (.A1(net242),
    .A2(_0654_),
    .A3(_0661_),
    .B1(_0657_),
    .B2(\as2650.r123_2[0][7] ),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(_0735_),
    .A1(_0736_),
    .S(_0643_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_2 _3856_ (.A(net303),
    .B(net234),
    .C(_2804_),
    .X(_0737_));
 sky130_fd_sc_hd__nand3_4 _3857_ (.A(net302),
    .B(net234),
    .C(_2804_),
    .Y(_0738_));
 sky130_fd_sc_hd__xor2_1 _3858_ (.A(\as2650.psl[7] ),
    .B(net304),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_1 _3859_ (.A(\as2650.psl[6] ),
    .B(net305),
    .Y(_0740_));
 sky130_fd_sc_hd__or2_1 _3860_ (.A(\as2650.psl[6] ),
    .B(net305),
    .X(_0741_));
 sky130_fd_sc_hd__a21oi_2 _3861_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0739_),
    .Y(_0742_));
 sky130_fd_sc_hd__or2_4 _3862_ (.A(net209),
    .B(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _3863_ (.A(net217),
    .B(net143),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a31o_1 _3864_ (.A1(net299),
    .A2(net136),
    .A3(_0743_),
    .B1(_0738_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_1 _3865_ (.A(_2789_),
    .B(net163),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_4 _3866_ (.A(_2790_),
    .B(_0738_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_2 _3867_ (.A(_2758_),
    .B(_2773_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_2 _3868_ (.A(net128),
    .B(net127),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_2 _3869_ (.A(net304),
    .B(net202),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_4 _3870_ (.A(_2806_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__or2_2 _3871_ (.A(_2806_),
    .B(_0750_),
    .X(_0752_));
 sky130_fd_sc_hd__or2_1 _3872_ (.A(_0586_),
    .B(_0751_),
    .X(_0753_));
 sky130_fd_sc_hd__or2_2 _3873_ (.A(net306),
    .B(_0750_),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_2 _3874_ (.A(_2809_),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor2_1 _3875_ (.A(_0753_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__or3b_1 _3876_ (.A(net88),
    .B(_2937_),
    .C_N(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_4 _3877_ (.A(net305),
    .B(_0752_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand2_2 _3878_ (.A(_2643_),
    .B(_0751_),
    .Y(_0759_));
 sky130_fd_sc_hd__or2_4 _3879_ (.A(_2726_),
    .B(_2794_),
    .X(_0760_));
 sky130_fd_sc_hd__and2_4 _3880_ (.A(net302),
    .B(net216),
    .X(_0761_));
 sky130_fd_sc_hd__or3b_4 _3881_ (.A(_2755_),
    .B(_2788_),
    .C_N(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_2 _3882_ (.A(_2810_),
    .B(net105),
    .Y(_0763_));
 sky130_fd_sc_hd__or2_4 _3883_ (.A(_2810_),
    .B(net105),
    .X(_0764_));
 sky130_fd_sc_hd__a2111o_1 _3884_ (.A1(net161),
    .A2(_0763_),
    .B1(_0760_),
    .C1(net70),
    .D1(_2789_),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _3885_ (.A(net209),
    .B(net105),
    .Y(_0766_));
 sky130_fd_sc_hd__or4_2 _3886_ (.A(net158),
    .B(_0747_),
    .C(net70),
    .D(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__or4b_1 _3887_ (.A(net294),
    .B(net142),
    .C(_0765_),
    .D_N(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a2111oi_1 _3888_ (.A1(net95),
    .A2(_0751_),
    .B1(_0768_),
    .C1(_2937_),
    .D1(_0586_),
    .Y(_0769_));
 sky130_fd_sc_hd__o311a_1 _3889_ (.A1(_0747_),
    .A2(net70),
    .A3(_0757_),
    .B1(_0769_),
    .C1(_0745_),
    .X(_0770_));
 sky130_fd_sc_hd__or3_2 _3890_ (.A(_2937_),
    .B(_0753_),
    .C(_0755_),
    .X(_0771_));
 sky130_fd_sc_hd__or4_1 _3891_ (.A(net87),
    .B(_2789_),
    .C(net163),
    .D(net70),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_4 _3892_ (.A(_2806_),
    .B(_0754_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor3_1 _3893_ (.A(net134),
    .B(_2806_),
    .C(_0750_),
    .Y(_0774_));
 sky130_fd_sc_hd__or2_4 _3894_ (.A(net204),
    .B(net105),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _3895_ (.A0(\as2650.psu[5] ),
    .A1(_0775_),
    .S(net337),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _3896_ (.A0(net250),
    .A1(_0776_),
    .S(net132),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _3897_ (.A(_0738_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21oi_1 _3898_ (.A1(_0770_),
    .A2(_0778_),
    .B1(net322),
    .Y(_0779_));
 sky130_fd_sc_hd__o21a_1 _3899_ (.A1(\as2650.psu[5] ),
    .A2(_0770_),
    .B1(_0779_),
    .X(_0039_));
 sky130_fd_sc_hd__nor3_4 _3900_ (.A(net219),
    .B(net170),
    .C(net55),
    .Y(_0780_));
 sky130_fd_sc_hd__or3_4 _3901_ (.A(net219),
    .B(net170),
    .C(net55),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_8 _3902_ (.A(_0585_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(\as2650.stack[5][8] ),
    .A1(_0607_),
    .S(_0782_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _3904_ (.A0(\as2650.stack[5][9] ),
    .A1(_0610_),
    .S(_0782_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _3905_ (.A0(\as2650.stack[5][10] ),
    .A1(_0612_),
    .S(_0782_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\as2650.stack[5][11] ),
    .A1(_0614_),
    .S(_0782_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(\as2650.stack[5][12] ),
    .A1(_0616_),
    .S(_0782_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(\as2650.stack[5][13] ),
    .A1(_0618_),
    .S(_0782_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _3909_ (.A0(\as2650.stack[5][14] ),
    .A1(_0620_),
    .S(_0782_),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_8 _3910_ (.A(_2850_),
    .B(_0584_),
    .Y(_0783_));
 sky130_fd_sc_hd__or2_4 _3911_ (.A(_2850_),
    .B(_0584_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_4 _3912_ (.A(_2850_),
    .B(net56),
    .Y(_0785_));
 sky130_fd_sc_hd__or2_4 _3913_ (.A(_2850_),
    .B(net56),
    .X(_0786_));
 sky130_fd_sc_hd__nand2_8 _3914_ (.A(_0784_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(\as2650.stack[4][8] ),
    .A1(_0607_),
    .S(_0787_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(\as2650.stack[4][9] ),
    .A1(_0610_),
    .S(_0787_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(\as2650.stack[4][10] ),
    .A1(_0612_),
    .S(_0787_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _3918_ (.A0(\as2650.stack[4][11] ),
    .A1(_0614_),
    .S(_0787_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(\as2650.stack[4][12] ),
    .A1(_0616_),
    .S(_0787_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(\as2650.stack[4][13] ),
    .A1(_0618_),
    .S(_0787_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(\as2650.stack[4][14] ),
    .A1(_0620_),
    .S(_0787_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _3922_ (.A0(_2659_),
    .A1(_2896_),
    .S(net200),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _3923_ (.A(_0523_),
    .B(_0556_),
    .Y(_0789_));
 sky130_fd_sc_hd__o22a_1 _3924_ (.A1(_2922_),
    .A2(_2970_),
    .B1(_2984_),
    .B2(_2968_),
    .X(_0790_));
 sky130_fd_sc_hd__or2_2 _3925_ (.A(_0321_),
    .B(_0368_),
    .X(_0791_));
 sky130_fd_sc_hd__or3_1 _3926_ (.A(_0320_),
    .B(_0327_),
    .C(_0368_),
    .X(_0792_));
 sky130_fd_sc_hd__o211a_1 _3927_ (.A1(_0790_),
    .A2(_0791_),
    .B1(_0792_),
    .C1(_0426_),
    .X(_0793_));
 sky130_fd_sc_hd__o21a_1 _3928_ (.A1(_0422_),
    .A2(_0793_),
    .B1(_0478_),
    .X(_0794_));
 sky130_fd_sc_hd__o21a_1 _3929_ (.A1(_0475_),
    .A2(_0794_),
    .B1(_0524_),
    .X(_0795_));
 sky130_fd_sc_hd__o2bb2a_1 _3930_ (.A1_N(_0554_),
    .A2_N(_0563_),
    .B1(_0789_),
    .B2(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_2623_),
    .B(_0555_),
    .Y(_0797_));
 sky130_fd_sc_hd__a21bo_1 _3932_ (.A1(_0556_),
    .A2(_0557_),
    .B1_N(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(_0797_),
    .A1(_0798_),
    .S(_0796_),
    .X(_0799_));
 sky130_fd_sc_hd__a21o_1 _3934_ (.A1(_2799_),
    .A2(_0799_),
    .B1(net95),
    .X(_0800_));
 sky130_fd_sc_hd__or4_1 _3935_ (.A(net95),
    .B(_2970_),
    .C(_0422_),
    .D(_0475_),
    .X(_0801_));
 sky130_fd_sc_hd__o41a_1 _3936_ (.A1(_2924_),
    .A2(_0789_),
    .A3(_0791_),
    .A4(_0801_),
    .B1(_0800_),
    .X(_0802_));
 sky130_fd_sc_hd__or4_1 _3937_ (.A(_2934_),
    .B(_2986_),
    .C(_0333_),
    .D(_0434_),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_0489_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__a31o_1 _3939_ (.A1(_0382_),
    .A2(_0535_),
    .A3(_0804_),
    .B1(_0568_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _3940_ (.A(_2799_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__and3_4 _3941_ (.A(net214),
    .B(_2647_),
    .C(_2804_),
    .X(_0807_));
 sky130_fd_sc_hd__or4_1 _3942_ (.A(net243),
    .B(net247),
    .C(net251),
    .D(net254),
    .X(_0808_));
 sky130_fd_sc_hd__or4_1 _3943_ (.A(net260),
    .B(net264),
    .C(net265),
    .D(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_2628_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nor2_1 _3945_ (.A(_0807_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__a311o_1 _3946_ (.A1(_2896_),
    .A2(_0504_),
    .A3(_0807_),
    .B1(_0811_),
    .C1(net134),
    .X(_0812_));
 sky130_fd_sc_hd__o211a_1 _3947_ (.A1(_0802_),
    .A2(_0806_),
    .B1(_0812_),
    .C1(net214),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_8 _3948_ (.A(net237),
    .B(net163),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_2 _3949_ (.A(net215),
    .B(_0738_),
    .Y(_0815_));
 sky130_fd_sc_hd__and4_2 _3950_ (.A(net142),
    .B(_2790_),
    .C(net71),
    .D(_0814_),
    .X(_0816_));
 sky130_fd_sc_hd__nor3_4 _3951_ (.A(net208),
    .B(net198),
    .C(_2809_),
    .Y(_0817_));
 sky130_fd_sc_hd__or4bb_1 _3952_ (.A(_2794_),
    .B(_2804_),
    .C_N(net125),
    .D_N(_2865_),
    .X(_0818_));
 sky130_fd_sc_hd__nor2_2 _3953_ (.A(_0772_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__nor2_2 _3954_ (.A(_0771_),
    .B(_0817_),
    .Y(_0820_));
 sky130_fd_sc_hd__or4_1 _3955_ (.A(net133),
    .B(_0747_),
    .C(net70),
    .D(_0818_),
    .X(_0821_));
 sky130_fd_sc_hd__a22oi_4 _3956_ (.A1(net229),
    .A2(_0816_),
    .B1(_0819_),
    .B2(_0820_),
    .Y(_0822_));
 sky130_fd_sc_hd__nor2_2 _3957_ (.A(_2766_),
    .B(_2803_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_8 _3958_ (.A(net230),
    .B(net87),
    .Y(_0824_));
 sky130_fd_sc_hd__a22o_1 _3959_ (.A1(net96),
    .A2(_0823_),
    .B1(net59),
    .B2(net198),
    .X(_0825_));
 sky130_fd_sc_hd__or3_2 _3960_ (.A(net231),
    .B(_2757_),
    .C(_2803_),
    .X(_0826_));
 sky130_fd_sc_hd__nand2_1 _3961_ (.A(net136),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__a31o_2 _3962_ (.A1(net216),
    .A2(net158),
    .A3(net126),
    .B1(_0825_),
    .X(_0828_));
 sky130_fd_sc_hd__or2_4 _3963_ (.A(net87),
    .B(_0826_),
    .X(_0829_));
 sky130_fd_sc_hd__nor2_8 _3964_ (.A(net238),
    .B(_0738_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_2 _3965_ (.A(net215),
    .B(net163),
    .Y(_0831_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(net138),
    .B(_0755_),
    .Y(_0832_));
 sky130_fd_sc_hd__or3b_2 _3967_ (.A(_2937_),
    .B(_0586_),
    .C_N(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__or3_2 _3968_ (.A(net231),
    .B(net153),
    .C(net143),
    .X(_0834_));
 sky130_fd_sc_hd__and3_1 _3969_ (.A(_2728_),
    .B(_2733_),
    .C(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_4 _3970_ (.A(net297),
    .B(_2789_),
    .Y(_0836_));
 sky130_fd_sc_hd__or2_2 _3971_ (.A(net236),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nand2_2 _3972_ (.A(net234),
    .B(net134),
    .Y(_0838_));
 sky130_fd_sc_hd__o31a_1 _3973_ (.A1(net236),
    .A2(net136),
    .A3(net71),
    .B1(_0837_),
    .X(_0839_));
 sky130_fd_sc_hd__and3b_1 _3974_ (.A_N(_0767_),
    .B(_2647_),
    .C(net171),
    .X(_0840_));
 sky130_fd_sc_hd__or3_4 _3975_ (.A(net305),
    .B(net158),
    .C(net105),
    .X(_0841_));
 sky130_fd_sc_hd__nor2_2 _3976_ (.A(net294),
    .B(_2727_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(net218),
    .B(_2728_),
    .Y(_0843_));
 sky130_fd_sc_hd__or2_2 _3978_ (.A(net132),
    .B(_0826_),
    .X(_0844_));
 sky130_fd_sc_hd__and3_1 _3979_ (.A(net103),
    .B(_0842_),
    .C(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__or4_1 _3980_ (.A(net231),
    .B(_2767_),
    .C(_0807_),
    .D(_0827_),
    .X(_0846_));
 sky130_fd_sc_hd__and4b_1 _3981_ (.A_N(_2734_),
    .B(_0834_),
    .C(_0841_),
    .D(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__and3_1 _3982_ (.A(net210),
    .B(_0845_),
    .C(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__and3_1 _3983_ (.A(_0822_),
    .B(_0839_),
    .C(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__or4b_4 _3984_ (.A(_0828_),
    .B(_0833_),
    .C(_0840_),
    .D_N(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__a211o_1 _3985_ (.A1(_2900_),
    .A2(_0449_),
    .B1(net107),
    .C1(net127),
    .X(_0851_));
 sky130_fd_sc_hd__or4b_1 _3986_ (.A(net119),
    .B(net118),
    .C(_0358_),
    .D_N(_0503_),
    .X(_0852_));
 sky130_fd_sc_hd__or3b_1 _3987_ (.A(net128),
    .B(_0543_),
    .C_N(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(_2642_),
    .A1(_2644_),
    .S(net334),
    .X(_0854_));
 sky130_fd_sc_hd__a21oi_1 _3989_ (.A1(_0751_),
    .A2(_0810_),
    .B1(net91),
    .Y(_0855_));
 sky130_fd_sc_hd__o21ai_1 _3990_ (.A1(net243),
    .A2(_0751_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__o41a_1 _3991_ (.A1(_2643_),
    .A2(net95),
    .A3(net105),
    .A4(_0854_),
    .B1(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__o211a_1 _3992_ (.A1(_0749_),
    .A2(_0857_),
    .B1(_0853_),
    .C1(_2792_),
    .X(_0858_));
 sky130_fd_sc_hd__nand2_1 _3993_ (.A(_0851_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(net331),
    .B(net126),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(net234),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_2658_),
    .B(net126),
    .Y(_0862_));
 sky130_fd_sc_hd__or4_1 _3997_ (.A(net344),
    .B(net340),
    .C(net339),
    .D(net336),
    .X(_0863_));
 sky130_fd_sc_hd__or4_1 _3998_ (.A(net347),
    .B(net346),
    .C(_0862_),
    .D(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__and3b_1 _3999_ (.A_N(_0861_),
    .B(_0864_),
    .C(_0859_),
    .X(_0865_));
 sky130_fd_sc_hd__a21oi_1 _4000_ (.A1(_2642_),
    .A2(_0850_),
    .B1(net325),
    .Y(_0866_));
 sky130_fd_sc_hd__o31a_1 _4001_ (.A1(_0813_),
    .A2(_0850_),
    .A3(_0865_),
    .B1(_0866_),
    .X(_0054_));
 sky130_fd_sc_hd__o221a_1 _4002_ (.A1(net127),
    .A2(net106),
    .B1(_0543_),
    .B2(net128),
    .C1(_2792_),
    .X(_0867_));
 sky130_fd_sc_hd__and4_2 _4003_ (.A(net233),
    .B(net300),
    .C(_2672_),
    .D(_0761_),
    .X(_0868_));
 sky130_fd_sc_hd__o22a_1 _4004_ (.A1(\as2650.carry ),
    .A2(_2651_),
    .B1(_2654_),
    .B2(\as2650.psl[3] ),
    .X(_0869_));
 sky130_fd_sc_hd__o22a_1 _4005_ (.A1(\as2650.psl[1] ),
    .A2(_2652_),
    .B1(_2658_),
    .B2(\as2650.psl[6] ),
    .X(_0870_));
 sky130_fd_sc_hd__o221a_1 _4006_ (.A1(net223),
    .A2(_2655_),
    .B1(_2657_),
    .B2(\as2650.psl[5] ),
    .C1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__o221a_1 _4007_ (.A1(\as2650.psl[7] ),
    .A2(net312),
    .B1(_2653_),
    .B2(\as2650.overflow ),
    .C1(_0869_),
    .X(_0872_));
 sky130_fd_sc_hd__nand2_1 _4008_ (.A(\as2650.ins_reg[0] ),
    .B(_0868_),
    .Y(_0873_));
 sky130_fd_sc_hd__and4_1 _4009_ (.A(net305),
    .B(_0868_),
    .C(_0871_),
    .D(_0872_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(net347),
    .B(_2879_),
    .Y(_0875_));
 sky130_fd_sc_hd__o221a_1 _4011_ (.A1(_2654_),
    .A2(net113),
    .B1(net109),
    .B2(_2657_),
    .C1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__o22a_1 _4012_ (.A1(_2653_),
    .A2(net117),
    .B1(_0353_),
    .B2(_2655_),
    .X(_0877_));
 sky130_fd_sc_hd__o221a_1 _4013_ (.A1(_2652_),
    .A2(_2887_),
    .B1(net106),
    .B2(_2658_),
    .C1(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__o2111a_1 _4014_ (.A1(_2650_),
    .A2(net118),
    .B1(_0873_),
    .C1(_0876_),
    .D1(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _4015_ (.A1(_2643_),
    .A2(_0868_),
    .B1(_0874_),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__o22a_1 _4016_ (.A1(\as2650.psu[0] ),
    .A2(_2651_),
    .B1(_2658_),
    .B2(net29),
    .X(_0881_));
 sky130_fd_sc_hd__o221a_1 _4017_ (.A1(\as2650.psu[3] ),
    .A2(_2654_),
    .B1(_2655_),
    .B2(\as2650.psu[4] ),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__o221a_1 _4018_ (.A1(\as2650.psu[7] ),
    .A2(_2650_),
    .B1(_2657_),
    .B2(\as2650.psu[5] ),
    .C1(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__o221a_1 _4019_ (.A1(net226),
    .A2(_2652_),
    .B1(_2653_),
    .B2(\as2650.psu[2] ),
    .C1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__or3b_1 _4020_ (.A(net305),
    .B(_0884_),
    .C_N(_0868_),
    .X(_0885_));
 sky130_fd_sc_hd__o211a_1 _4021_ (.A1(net208),
    .A2(net105),
    .B1(_0880_),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or4_1 _4022_ (.A(\as2650.psl[7] ),
    .B(net331),
    .C(net208),
    .D(_0762_),
    .X(_0887_));
 sky130_fd_sc_hd__or3b_1 _4023_ (.A(_0763_),
    .B(_0886_),
    .C_N(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__o31a_1 _4024_ (.A1(_2641_),
    .A2(net331),
    .A3(_0764_),
    .B1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__nor2_1 _4025_ (.A(net96),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__a211o_1 _4026_ (.A1(net239),
    .A2(net96),
    .B1(_0749_),
    .C1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__a21o_1 _4027_ (.A1(_0867_),
    .A2(_0891_),
    .B1(_0861_),
    .X(_0892_));
 sky130_fd_sc_hd__o21ba_1 _4028_ (.A1(_2799_),
    .A2(_0568_),
    .B1_N(_0800_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(net242),
    .A1(net118),
    .S(_0807_),
    .X(_0894_));
 sky130_fd_sc_hd__a211o_1 _4030_ (.A1(net138),
    .A2(_0894_),
    .B1(_0893_),
    .C1(net234),
    .X(_0895_));
 sky130_fd_sc_hd__a21oi_1 _4031_ (.A1(_0892_),
    .A2(_0895_),
    .B1(_0850_),
    .Y(_0896_));
 sky130_fd_sc_hd__a211oi_1 _4032_ (.A1(_2641_),
    .A2(_0850_),
    .B1(_0896_),
    .C1(net325),
    .Y(_0055_));
 sky130_fd_sc_hd__or2_4 _4033_ (.A(net227),
    .B(net190),
    .X(_0897_));
 sky130_fd_sc_hd__or2_4 _4034_ (.A(net56),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_2 _4035_ (.A(net49),
    .B(_0897_),
    .Y(_0899_));
 sky130_fd_sc_hd__or2_4 _4036_ (.A(net49),
    .B(_0897_),
    .X(_0900_));
 sky130_fd_sc_hd__nand2_8 _4037_ (.A(_0898_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(\as2650.stack[3][8] ),
    .A1(_0607_),
    .S(_0901_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(\as2650.stack[3][9] ),
    .A1(_0610_),
    .S(_0901_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(\as2650.stack[3][10] ),
    .A1(_0612_),
    .S(_0901_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(\as2650.stack[3][11] ),
    .A1(_0614_),
    .S(_0901_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(\as2650.stack[3][12] ),
    .A1(_0616_),
    .S(_0901_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(\as2650.stack[3][13] ),
    .A1(_0618_),
    .S(_0901_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(\as2650.stack[3][14] ),
    .A1(_0620_),
    .S(_0901_),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _4045_ (.A1(net312),
    .A2(net161),
    .B1(net145),
    .B2(_2728_),
    .X(_0902_));
 sky130_fd_sc_hd__or4_4 _4046_ (.A(net217),
    .B(_2669_),
    .C(net206),
    .D(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__nor2_4 _4047_ (.A(_2728_),
    .B(net206),
    .Y(_0904_));
 sky130_fd_sc_hd__nor3_1 _4048_ (.A(net211),
    .B(_2727_),
    .C(_0903_),
    .Y(_0905_));
 sky130_fd_sc_hd__a221o_1 _4049_ (.A1(net306),
    .A2(_0903_),
    .B1(_0904_),
    .B2(net349),
    .C1(_0905_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(net346),
    .A1(net173),
    .S(_2728_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(_0906_),
    .A1(net304),
    .S(_0903_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _4052_ (.A1(net302),
    .A2(_0903_),
    .B1(_0904_),
    .B2(net344),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4053_ (.A0(net299),
    .A1(net337),
    .S(_0904_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _4054_ (.A1(\as2650.ins_reg[6] ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(net335),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _4055_ (.A1(net297),
    .A2(_0903_),
    .B1(_0904_),
    .B2(net328),
    .X(_0068_));
 sky130_fd_sc_hd__or3_4 _4056_ (.A(net227),
    .B(net164),
    .C(net49),
    .X(_0907_));
 sky130_fd_sc_hd__nor3_2 _4057_ (.A(net227),
    .B(net164),
    .C(net56),
    .Y(_0908_));
 sky130_fd_sc_hd__or3_4 _4058_ (.A(net227),
    .B(net164),
    .C(net56),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_8 _4059_ (.A(_0907_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(\as2650.stack[2][8] ),
    .A1(_0607_),
    .S(_0910_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4061_ (.A0(\as2650.stack[2][9] ),
    .A1(_0610_),
    .S(_0910_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(\as2650.stack[2][10] ),
    .A1(_0612_),
    .S(_0910_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(\as2650.stack[2][11] ),
    .A1(_0614_),
    .S(_0910_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(\as2650.stack[2][12] ),
    .A1(_0616_),
    .S(_0910_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(\as2650.stack[2][13] ),
    .A1(_0618_),
    .S(_0910_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(\as2650.stack[2][14] ),
    .A1(_0620_),
    .S(_0910_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_4 _4067_ (.A(net307),
    .B(_0642_),
    .X(_0911_));
 sky130_fd_sc_hd__inv_2 _4068_ (.A(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_1 _4069_ (.A(_0652_),
    .B(_0911_),
    .Y(_0913_));
 sky130_fd_sc_hd__o31ai_4 _4070_ (.A1(net296),
    .A2(_2865_),
    .A3(_0655_),
    .B1(net318),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_8 _4071_ (.A(_0912_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor4b_4 _4072_ (.A(net90),
    .B(_0603_),
    .C(_0915_),
    .D_N(_2937_),
    .Y(_0916_));
 sky130_fd_sc_hd__a31o_1 _4073_ (.A1(net266),
    .A2(_0605_),
    .A3(net42),
    .B1(_0913_),
    .X(_0917_));
 sky130_fd_sc_hd__a21o_1 _4074_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_0915_),
    .B1(_0917_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_2 _4075_ (.A(net262),
    .B(net176),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _4076_ (.A(net266),
    .B(net174),
    .Y(_0919_));
 sky130_fd_sc_hd__and4_1 _4077_ (.A(net262),
    .B(net266),
    .C(net176),
    .D(net174),
    .X(_0920_));
 sky130_fd_sc_hd__a21oi_1 _4078_ (.A1(_0918_),
    .A2(_0919_),
    .B1(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__a2bb2o_1 _4079_ (.A1_N(_0670_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][1] ),
    .X(_0922_));
 sky130_fd_sc_hd__a21o_1 _4080_ (.A1(net42),
    .A2(_0921_),
    .B1(_0922_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _4081_ (.A1(net258),
    .A2(net176),
    .B1(net174),
    .B2(net263),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_2 _4082_ (.A(net258),
    .B(net174),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_4 _4083_ (.A(_0918_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__or2_1 _4084_ (.A(_0918_),
    .B(_0924_),
    .X(_0926_));
 sky130_fd_sc_hd__and4_4 _4085_ (.A(net268),
    .B(net186),
    .C(_0923_),
    .D(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__a22oi_1 _4086_ (.A1(net266),
    .A2(net186),
    .B1(_0923_),
    .B2(_0926_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _4087_ (.A(_0927_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand2_2 _4088_ (.A(_0920_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__or2_1 _4089_ (.A(_0920_),
    .B(_0929_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _4090_ (.A(_0930_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__a2bb2o_1 _4091_ (.A1_N(_0681_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][2] ),
    .X(_0933_));
 sky130_fd_sc_hd__a21o_1 _4092_ (.A1(net42),
    .A2(_0932_),
    .B1(_0933_),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(net255),
    .B(net177),
    .Y(_0934_));
 sky130_fd_sc_hd__and4_1 _4094_ (.A(net255),
    .B(net258),
    .C(net177),
    .D(net175),
    .X(_0935_));
 sky130_fd_sc_hd__a21o_2 _4095_ (.A1(_0924_),
    .A2(_0934_),
    .B1(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__and4_1 _4096_ (.A(net263),
    .B(net266),
    .C(net186),
    .D(net184),
    .X(_0937_));
 sky130_fd_sc_hd__a22oi_1 _4097_ (.A1(net263),
    .A2(net187),
    .B1(net185),
    .B2(net267),
    .Y(_0938_));
 sky130_fd_sc_hd__or2_4 _4098_ (.A(_0937_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__xor2_4 _4099_ (.A(_0936_),
    .B(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__o21ai_4 _4100_ (.A1(_0925_),
    .A2(_0927_),
    .B1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__o31ai_4 _4101_ (.A1(_0925_),
    .A2(_0927_),
    .A3(_0940_),
    .B1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__or2_2 _4102_ (.A(_0930_),
    .B(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__xor2_2 _4103_ (.A(_0930_),
    .B(_0942_),
    .X(_0944_));
 sky130_fd_sc_hd__a2bb2o_1 _4104_ (.A1_N(_0692_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][3] ),
    .X(_0945_));
 sky130_fd_sc_hd__a21o_1 _4105_ (.A1(net41),
    .A2(_0944_),
    .B1(_0945_),
    .X(_0079_));
 sky130_fd_sc_hd__a21oi_1 _4106_ (.A1(net255),
    .A2(net174),
    .B1(_0937_),
    .Y(_0946_));
 sky130_fd_sc_hd__and3_1 _4107_ (.A(net255),
    .B(net174),
    .C(_0937_),
    .X(_0947_));
 sky130_fd_sc_hd__nor2_2 _4108_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2_1 _4109_ (.A(net253),
    .B(net176),
    .Y(_0949_));
 sky130_fd_sc_hd__xor2_2 _4110_ (.A(_0948_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_2 _4111_ (.A(net259),
    .B(net187),
    .Y(_0951_));
 sky130_fd_sc_hd__and4_1 _4112_ (.A(net262),
    .B(net267),
    .C(net185),
    .D(net183),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(net262),
    .A2(net185),
    .B1(net183),
    .B2(net267),
    .X(_0953_));
 sky130_fd_sc_hd__and2b_2 _4114_ (.A_N(_0952_),
    .B(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__xnor2_4 _4115_ (.A(_0951_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2b_4 _4116_ (.A_N(_0950_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__xnor2_1 _4117_ (.A(_0950_),
    .B(_0955_),
    .Y(_0957_));
 sky130_fd_sc_hd__o21bai_1 _4118_ (.A1(_0936_),
    .A2(_0939_),
    .B1_N(_0935_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_1 _4119_ (.A(_0957_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _4120_ (.A(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(_0957_),
    .B(_0958_),
    .Y(_0961_));
 sky130_fd_sc_hd__or2_1 _4122_ (.A(_0960_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__nor2_1 _4123_ (.A(_0941_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2_1 _4124_ (.A(_0943_),
    .B(_0962_),
    .Y(_0964_));
 sky130_fd_sc_hd__and2_1 _4125_ (.A(_0943_),
    .B(_0962_),
    .X(_0965_));
 sky130_fd_sc_hd__or2_1 _4126_ (.A(_0964_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__a21oi_1 _4127_ (.A1(_0941_),
    .A2(_0966_),
    .B1(_0963_),
    .Y(_0967_));
 sky130_fd_sc_hd__a2bb2o_1 _4128_ (.A1_N(_0703_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][4] ),
    .X(_0968_));
 sky130_fd_sc_hd__a21o_1 _4129_ (.A1(net41),
    .A2(_0967_),
    .B1(_0968_),
    .X(_0080_));
 sky130_fd_sc_hd__a31o_2 _4130_ (.A1(net253),
    .A2(net176),
    .A3(_0948_),
    .B1(_0947_),
    .X(_0969_));
 sky130_fd_sc_hd__and2_1 _4131_ (.A(net256),
    .B(net186),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _4132_ (.A1(net258),
    .A2(net185),
    .B1(net183),
    .B2(net262),
    .X(_0971_));
 sky130_fd_sc_hd__nand4_2 _4133_ (.A(net258),
    .B(net262),
    .C(net184),
    .D(net182),
    .Y(_0972_));
 sky130_fd_sc_hd__a21o_1 _4134_ (.A1(_0971_),
    .A2(_0972_),
    .B1(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__nand3_1 _4135_ (.A(_0970_),
    .B(_0971_),
    .C(_0972_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(net266),
    .B(net181),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__and3_2 _4138_ (.A(_0973_),
    .B(_0974_),
    .C(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a21oi_1 _4139_ (.A1(_0973_),
    .A2(_0974_),
    .B1(_0976_),
    .Y(_0978_));
 sky130_fd_sc_hd__or2_4 _4140_ (.A(_0977_),
    .B(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__nand2_2 _4141_ (.A(net248),
    .B(net176),
    .Y(_0980_));
 sky130_fd_sc_hd__a31o_4 _4142_ (.A1(net259),
    .A2(net187),
    .A3(_0953_),
    .B1(_0952_),
    .X(_0981_));
 sky130_fd_sc_hd__nand2_2 _4143_ (.A(net253),
    .B(net174),
    .Y(_0982_));
 sky130_fd_sc_hd__and3_1 _4144_ (.A(net253),
    .B(net174),
    .C(_0981_),
    .X(_0983_));
 sky130_fd_sc_hd__xnor2_4 _4145_ (.A(_0981_),
    .B(_0982_),
    .Y(_0984_));
 sky130_fd_sc_hd__xnor2_4 _4146_ (.A(_0980_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__and2b_2 _4147_ (.A_N(_0979_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__xnor2_4 _4148_ (.A(_0979_),
    .B(_0985_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2b_2 _4149_ (.A_N(_0956_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__xnor2_4 _4150_ (.A(_0956_),
    .B(_0987_),
    .Y(_0989_));
 sky130_fd_sc_hd__nand2_2 _4151_ (.A(_0969_),
    .B(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__xnor2_2 _4152_ (.A(_0969_),
    .B(_0989_),
    .Y(_0991_));
 sky130_fd_sc_hd__or2_2 _4153_ (.A(_0959_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_1 _4154_ (.A(_0959_),
    .B(_0991_),
    .Y(_0993_));
 sky130_fd_sc_hd__a2111o_4 _4155_ (.A1(_0941_),
    .A2(_0943_),
    .B1(_0960_),
    .C1(_0961_),
    .D1(_0991_),
    .X(_0994_));
 sky130_fd_sc_hd__a211o_1 _4156_ (.A1(_0992_),
    .A2(_0993_),
    .B1(_0963_),
    .C1(_0964_),
    .X(_0995_));
 sky130_fd_sc_hd__and2_1 _4157_ (.A(_0994_),
    .B(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__a2bb2o_1 _4158_ (.A1_N(_0714_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][5] ),
    .X(_0997_));
 sky130_fd_sc_hd__a21o_1 _4159_ (.A1(net42),
    .A2(_0996_),
    .B1(_0997_),
    .X(_0081_));
 sky130_fd_sc_hd__a31o_4 _4160_ (.A1(net248),
    .A2(net176),
    .A3(_0984_),
    .B1(_0983_),
    .X(_0998_));
 sky130_fd_sc_hd__a22o_1 _4161_ (.A1(net256),
    .A2(net184),
    .B1(net182),
    .B2(net258),
    .X(_0999_));
 sky130_fd_sc_hd__nand4_4 _4162_ (.A(net255),
    .B(net258),
    .C(net184),
    .D(net182),
    .Y(_1000_));
 sky130_fd_sc_hd__and2_1 _4163_ (.A(net253),
    .B(net186),
    .X(_1001_));
 sky130_fd_sc_hd__a21o_1 _4164_ (.A1(_0999_),
    .A2(_1000_),
    .B1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__nand3_2 _4165_ (.A(_0999_),
    .B(_1000_),
    .C(_1001_),
    .Y(_1003_));
 sky130_fd_sc_hd__a22oi_2 _4166_ (.A1(net262),
    .A2(net181),
    .B1(net179),
    .B2(net267),
    .Y(_1004_));
 sky130_fd_sc_hd__and4_2 _4167_ (.A(net262),
    .B(net267),
    .C(net181),
    .D(net179),
    .X(_1005_));
 sky130_fd_sc_hd__nor2_2 _4168_ (.A(_1004_),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand3_4 _4169_ (.A(_1002_),
    .B(_1003_),
    .C(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__a21o_2 _4170_ (.A1(_1002_),
    .A2(_1003_),
    .B1(_1006_),
    .X(_1008_));
 sky130_fd_sc_hd__nand3_4 _4171_ (.A(_0977_),
    .B(_1007_),
    .C(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a21o_1 _4172_ (.A1(_1007_),
    .A2(_1008_),
    .B1(_0977_),
    .X(_1010_));
 sky130_fd_sc_hd__nand2_2 _4173_ (.A(net245),
    .B(net176),
    .Y(_1011_));
 sky130_fd_sc_hd__a21bo_4 _4174_ (.A1(_0970_),
    .A2(_0971_),
    .B1_N(_0972_),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_2 _4175_ (.A(net248),
    .B(net174),
    .Y(_1013_));
 sky130_fd_sc_hd__and3_1 _4176_ (.A(net248),
    .B(net174),
    .C(_1012_),
    .X(_1014_));
 sky130_fd_sc_hd__xnor2_4 _4177_ (.A(_1012_),
    .B(_1013_),
    .Y(_1015_));
 sky130_fd_sc_hd__xnor2_4 _4178_ (.A(_1011_),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a21o_2 _4179_ (.A1(_1009_),
    .A2(_1010_),
    .B1(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__nand3_4 _4180_ (.A(_1009_),
    .B(_1010_),
    .C(_1016_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand3_4 _4181_ (.A(_0986_),
    .B(_1017_),
    .C(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__a21o_2 _4182_ (.A1(_1017_),
    .A2(_1018_),
    .B1(_0986_),
    .X(_1020_));
 sky130_fd_sc_hd__a21oi_4 _4183_ (.A1(_1019_),
    .A2(_1020_),
    .B1(_0998_),
    .Y(_1021_));
 sky130_fd_sc_hd__and3_2 _4184_ (.A(_0998_),
    .B(_1019_),
    .C(_1020_),
    .X(_1022_));
 sky130_fd_sc_hd__nand3_4 _4185_ (.A(_0998_),
    .B(_1019_),
    .C(_1020_),
    .Y(_1023_));
 sky130_fd_sc_hd__a211oi_4 _4186_ (.A1(_0988_),
    .A2(_0990_),
    .B1(_1021_),
    .C1(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__o211a_2 _4187_ (.A1(_1021_),
    .A2(_1022_),
    .B1(_0988_),
    .C1(_0990_),
    .X(_1025_));
 sky130_fd_sc_hd__a211oi_4 _4188_ (.A1(_0992_),
    .A2(_0994_),
    .B1(_1024_),
    .C1(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__o211a_1 _4189_ (.A1(_1024_),
    .A2(_1025_),
    .B1(_0992_),
    .C1(_0994_),
    .X(_1027_));
 sky130_fd_sc_hd__nor2_2 _4190_ (.A(_1026_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__a2bb2o_1 _4191_ (.A1_N(_0724_),
    .A2_N(_0911_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][6] ),
    .X(_1029_));
 sky130_fd_sc_hd__a21o_1 _4192_ (.A1(net42),
    .A2(_1028_),
    .B1(_1029_),
    .X(_0082_));
 sky130_fd_sc_hd__nor2_1 _4193_ (.A(_1024_),
    .B(_1026_),
    .Y(_1030_));
 sky130_fd_sc_hd__a31o_2 _4194_ (.A1(net245),
    .A2(net176),
    .A3(_1015_),
    .B1(_1014_),
    .X(_1031_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(net259),
    .B(net180),
    .Y(_1032_));
 sky130_fd_sc_hd__a22o_2 _4196_ (.A1(net267),
    .A2(_2893_),
    .B1(net179),
    .B2(net262),
    .X(_1033_));
 sky130_fd_sc_hd__nand4_4 _4197_ (.A(net262),
    .B(net267),
    .C(net188),
    .D(net178),
    .Y(_1034_));
 sky130_fd_sc_hd__a21bo_2 _4198_ (.A1(_1033_),
    .A2(_1034_),
    .B1_N(_1032_),
    .X(_1035_));
 sky130_fd_sc_hd__nand3b_4 _4199_ (.A_N(_1032_),
    .B(_1033_),
    .C(_1034_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand3_4 _4200_ (.A(_1005_),
    .B(_1035_),
    .C(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a21o_2 _4201_ (.A1(_1035_),
    .A2(_1036_),
    .B1(_1005_),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_2 _4202_ (.A(net248),
    .B(net186),
    .Y(_1039_));
 sky130_fd_sc_hd__a22oi_4 _4203_ (.A1(net252),
    .A2(net184),
    .B1(net182),
    .B2(net255),
    .Y(_1040_));
 sky130_fd_sc_hd__and4_2 _4204_ (.A(net252),
    .B(net256),
    .C(net184),
    .D(net182),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_4 _4205_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__and3_1 _4206_ (.A(net249),
    .B(net186),
    .C(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__xnor2_4 _4207_ (.A(_1039_),
    .B(_1042_),
    .Y(_1044_));
 sky130_fd_sc_hd__a21oi_4 _4208_ (.A1(_1037_),
    .A2(_1038_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__and3_2 _4209_ (.A(_1037_),
    .B(_1038_),
    .C(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__or3_4 _4210_ (.A(_1007_),
    .B(_1045_),
    .C(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__o21ai_4 _4211_ (.A1(_1045_),
    .A2(_1046_),
    .B1(_1007_),
    .Y(_1048_));
 sky130_fd_sc_hd__a21bo_1 _4212_ (.A1(_0999_),
    .A2(_1001_),
    .B1_N(_1000_),
    .X(_1049_));
 sky130_fd_sc_hd__nand2_1 _4213_ (.A(net245),
    .B(net175),
    .Y(_1050_));
 sky130_fd_sc_hd__and3_2 _4214_ (.A(net245),
    .B(net175),
    .C(_1049_),
    .X(_1051_));
 sky130_fd_sc_hd__xnor2_1 _4215_ (.A(_1049_),
    .B(_1050_),
    .Y(_1052_));
 sky130_fd_sc_hd__and3_2 _4216_ (.A(net241),
    .B(net177),
    .C(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__a21oi_1 _4217_ (.A1(net241),
    .A2(net177),
    .B1(_1052_),
    .Y(_1054_));
 sky130_fd_sc_hd__nor2_2 _4218_ (.A(_1053_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__a21oi_4 _4219_ (.A1(_1047_),
    .A2(_1048_),
    .B1(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__and3_2 _4220_ (.A(_1047_),
    .B(_1048_),
    .C(_1055_),
    .X(_1057_));
 sky130_fd_sc_hd__nand3_2 _4221_ (.A(_1047_),
    .B(_1048_),
    .C(_1055_),
    .Y(_1058_));
 sky130_fd_sc_hd__o211ai_4 _4222_ (.A1(_1056_),
    .A2(_1057_),
    .B1(_1009_),
    .C1(_1018_),
    .Y(_1059_));
 sky130_fd_sc_hd__a211o_2 _4223_ (.A1(_1009_),
    .A2(_1018_),
    .B1(_1056_),
    .C1(_1057_),
    .X(_1060_));
 sky130_fd_sc_hd__a21oi_4 _4224_ (.A1(_1059_),
    .A2(_1060_),
    .B1(_1031_),
    .Y(_1061_));
 sky130_fd_sc_hd__and3_2 _4225_ (.A(_1031_),
    .B(_1059_),
    .C(_1060_),
    .X(_1062_));
 sky130_fd_sc_hd__a211oi_4 _4226_ (.A1(_1019_),
    .A2(_1023_),
    .B1(_1061_),
    .C1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__a211o_1 _4227_ (.A1(_1019_),
    .A2(_1023_),
    .B1(_1061_),
    .C1(_1062_),
    .X(_1064_));
 sky130_fd_sc_hd__o211ai_2 _4228_ (.A1(_1061_),
    .A2(_1062_),
    .B1(_1019_),
    .C1(_1023_),
    .Y(_1065_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(_1064_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__o211a_2 _4230_ (.A1(_1024_),
    .A2(_1026_),
    .B1(_1064_),
    .C1(_1065_),
    .X(_1067_));
 sky130_fd_sc_hd__xor2_2 _4231_ (.A(_1030_),
    .B(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__a22o_1 _4232_ (.A1(_0735_),
    .A2(_0912_),
    .B1(_0915_),
    .B2(\as2650.r123_2[1][7] ),
    .X(_1069_));
 sky130_fd_sc_hd__a21o_1 _4233_ (.A1(net42),
    .A2(_1068_),
    .B1(_1069_),
    .X(_0083_));
 sky130_fd_sc_hd__or2_2 _4234_ (.A(net227),
    .B(net168),
    .X(_1070_));
 sky130_fd_sc_hd__nor2_2 _4235_ (.A(net49),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__or2_4 _4236_ (.A(net49),
    .B(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_1 _4237_ (.A(net56),
    .B(_1070_),
    .Y(_1073_));
 sky130_fd_sc_hd__or2_4 _4238_ (.A(net56),
    .B(_1070_),
    .X(_1074_));
 sky130_fd_sc_hd__nand2_8 _4239_ (.A(_1072_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(\as2650.stack[1][8] ),
    .A1(_0607_),
    .S(_1075_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(\as2650.stack[1][9] ),
    .A1(_0610_),
    .S(_1075_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(\as2650.stack[1][10] ),
    .A1(_0612_),
    .S(_1075_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(\as2650.stack[1][11] ),
    .A1(_0614_),
    .S(_1075_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(\as2650.stack[1][12] ),
    .A1(_0616_),
    .S(_1075_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(\as2650.stack[1][13] ),
    .A1(_0618_),
    .S(_1075_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(\as2650.stack[1][14] ),
    .A1(_0620_),
    .S(_1075_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_8 _4247_ (.A(net219),
    .B(net195),
    .Y(_1076_));
 sky130_fd_sc_hd__nor2_1 _4248_ (.A(net49),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__or2_4 _4249_ (.A(net49),
    .B(_1076_),
    .X(_1078_));
 sky130_fd_sc_hd__nor2_8 _4250_ (.A(net55),
    .B(_1076_),
    .Y(_1079_));
 sky130_fd_sc_hd__or2_4 _4251_ (.A(net55),
    .B(_1076_),
    .X(_1080_));
 sky130_fd_sc_hd__nand2_8 _4252_ (.A(_1078_),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(\as2650.stack[0][8] ),
    .A1(_0607_),
    .S(_1081_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(\as2650.stack[0][9] ),
    .A1(_0610_),
    .S(_1081_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(\as2650.stack[0][10] ),
    .A1(_0612_),
    .S(_1081_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\as2650.stack[0][11] ),
    .A1(_0614_),
    .S(_1081_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(\as2650.stack[0][12] ),
    .A1(_0616_),
    .S(_1081_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\as2650.stack[0][13] ),
    .A1(_0618_),
    .S(_1081_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(\as2650.stack[0][14] ),
    .A1(_0620_),
    .S(_1081_),
    .X(_0097_));
 sky130_fd_sc_hd__o211a_2 _4260_ (.A1(_1041_),
    .A2(_1043_),
    .B1(net241),
    .C1(net175),
    .X(_1082_));
 sky130_fd_sc_hd__a211oi_1 _4261_ (.A1(net241),
    .A2(net175),
    .B1(_1041_),
    .C1(_1043_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _4262_ (.A(_1082_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__a22oi_4 _4263_ (.A1(net249),
    .A2(net184),
    .B1(net182),
    .B2(net252),
    .Y(_1085_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(net249),
    .B(net182),
    .Y(_1086_));
 sky130_fd_sc_hd__and4_1 _4265_ (.A(net249),
    .B(net252),
    .C(net184),
    .D(net182),
    .X(_1087_));
 sky130_fd_sc_hd__or2_4 _4266_ (.A(_1085_),
    .B(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_4 _4267_ (.A(net244),
    .B(net186),
    .Y(_1089_));
 sky130_fd_sc_hd__xnor2_4 _4268_ (.A(_1088_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_2 _4269_ (.A(net259),
    .B(net188),
    .Y(_1091_));
 sky130_fd_sc_hd__and4_2 _4270_ (.A(net259),
    .B(net264),
    .C(net188),
    .D(net178),
    .X(_1092_));
 sky130_fd_sc_hd__a22oi_4 _4271_ (.A1(net264),
    .A2(_2893_),
    .B1(net178),
    .B2(net259),
    .Y(_1093_));
 sky130_fd_sc_hd__nor2_4 _4272_ (.A(_1092_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_2 _4273_ (.A(net256),
    .B(net180),
    .Y(_1095_));
 sky130_fd_sc_hd__xnor2_4 _4274_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__and2_2 _4275_ (.A(_1034_),
    .B(_1036_),
    .X(_1097_));
 sky130_fd_sc_hd__nand2b_1 _4276_ (.A_N(_1097_),
    .B(_1096_),
    .Y(_1098_));
 sky130_fd_sc_hd__xor2_4 _4277_ (.A(_1096_),
    .B(_1097_),
    .X(_1099_));
 sky130_fd_sc_hd__xor2_4 _4278_ (.A(_1090_),
    .B(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__a21boi_4 _4279_ (.A1(_1038_),
    .A2(_1044_),
    .B1_N(_1037_),
    .Y(_1101_));
 sky130_fd_sc_hd__and2b_1 _4280_ (.A_N(_1101_),
    .B(_1100_),
    .X(_1102_));
 sky130_fd_sc_hd__xnor2_2 _4281_ (.A(_1100_),
    .B(_1101_),
    .Y(_1103_));
 sky130_fd_sc_hd__and2_2 _4282_ (.A(_1084_),
    .B(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__nor2_2 _4283_ (.A(_1084_),
    .B(_1103_),
    .Y(_1105_));
 sky130_fd_sc_hd__a211o_2 _4284_ (.A1(_1047_),
    .A2(_1058_),
    .B1(_1104_),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__o211ai_4 _4285_ (.A1(_1104_),
    .A2(_1105_),
    .B1(_1047_),
    .C1(_1058_),
    .Y(_1107_));
 sky130_fd_sc_hd__o211ai_4 _4286_ (.A1(_1051_),
    .A2(_1053_),
    .B1(_1106_),
    .C1(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__a211o_2 _4287_ (.A1(_1106_),
    .A2(_1107_),
    .B1(_1051_),
    .C1(_1053_),
    .X(_1109_));
 sky130_fd_sc_hd__a21bo_2 _4288_ (.A1(_1031_),
    .A2(_1059_),
    .B1_N(_1060_),
    .X(_1110_));
 sky130_fd_sc_hd__nand3_4 _4289_ (.A(_1108_),
    .B(_1109_),
    .C(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__a21o_1 _4290_ (.A1(_1108_),
    .A2(_1109_),
    .B1(_1110_),
    .X(_1112_));
 sky130_fd_sc_hd__o211ai_4 _4291_ (.A1(_1063_),
    .A2(_1067_),
    .B1(_1111_),
    .C1(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__a211o_1 _4292_ (.A1(_1111_),
    .A2(_1112_),
    .B1(_1063_),
    .C1(_1067_),
    .X(_1114_));
 sky130_fd_sc_hd__and2_1 _4293_ (.A(_1113_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__or2_4 _4294_ (.A(net207),
    .B(_0642_),
    .X(_1116_));
 sky130_fd_sc_hd__inv_2 _4295_ (.A(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__nor2_4 _4296_ (.A(_0914_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__a22oi_1 _4297_ (.A1(net41),
    .A2(_1115_),
    .B1(_1118_),
    .B2(\as2650.r123_2[2][0] ),
    .Y(_1119_));
 sky130_fd_sc_hd__o21ai_1 _4298_ (.A1(_0652_),
    .A2(_1116_),
    .B1(_1119_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ba_4 _4299_ (.A1(_1085_),
    .A2(_1089_),
    .B1_N(_1087_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _4300_ (.A(net256),
    .B(net188),
    .Y(_1121_));
 sky130_fd_sc_hd__nand2_2 _4301_ (.A(net256),
    .B(net178),
    .Y(_1122_));
 sky130_fd_sc_hd__xor2_2 _4302_ (.A(_1091_),
    .B(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__and3_2 _4303_ (.A(net252),
    .B(net180),
    .C(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a21oi_2 _4304_ (.A1(net252),
    .A2(net180),
    .B1(_1123_),
    .Y(_1125_));
 sky130_fd_sc_hd__nor2_4 _4305_ (.A(_1124_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__a31o_2 _4306_ (.A1(net256),
    .A2(net180),
    .A3(_1094_),
    .B1(_1092_),
    .X(_1127_));
 sky130_fd_sc_hd__and2_1 _4307_ (.A(_1126_),
    .B(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__xnor2_4 _4308_ (.A(_1126_),
    .B(_1127_),
    .Y(_1129_));
 sky130_fd_sc_hd__nand2_2 _4309_ (.A(net244),
    .B(net184),
    .Y(_1130_));
 sky130_fd_sc_hd__xor2_1 _4310_ (.A(_1086_),
    .B(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__and3_1 _4311_ (.A(net240),
    .B(net186),
    .C(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__a21oi_1 _4312_ (.A1(net240),
    .A2(net186),
    .B1(_1131_),
    .Y(_1133_));
 sky130_fd_sc_hd__or2_4 _4313_ (.A(_1132_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_1 _4314_ (.A(_1129_),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__xor2_4 _4315_ (.A(_1129_),
    .B(_1134_),
    .X(_1136_));
 sky130_fd_sc_hd__o21a_2 _4316_ (.A1(_1090_),
    .A2(_1099_),
    .B1(_1098_),
    .X(_1137_));
 sky130_fd_sc_hd__and2b_1 _4317_ (.A_N(_1137_),
    .B(_1136_),
    .X(_1138_));
 sky130_fd_sc_hd__xnor2_4 _4318_ (.A(_1136_),
    .B(_1137_),
    .Y(_1139_));
 sky130_fd_sc_hd__and2b_1 _4319_ (.A_N(_1120_),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__xnor2_4 _4320_ (.A(_1120_),
    .B(_1139_),
    .Y(_1141_));
 sky130_fd_sc_hd__nor2_2 _4321_ (.A(_1102_),
    .B(_1104_),
    .Y(_1142_));
 sky130_fd_sc_hd__and2b_1 _4322_ (.A_N(_1142_),
    .B(_1141_),
    .X(_1143_));
 sky130_fd_sc_hd__xnor2_2 _4323_ (.A(_1141_),
    .B(_1142_),
    .Y(_1144_));
 sky130_fd_sc_hd__and2_1 _4324_ (.A(_1082_),
    .B(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__xnor2_2 _4325_ (.A(_1082_),
    .B(_1144_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4326_ (.A(_1106_),
    .B(_1108_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2b_2 _4327_ (.A_N(_1146_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__xor2_1 _4328_ (.A(_1146_),
    .B(_1147_),
    .X(_1149_));
 sky130_fd_sc_hd__a21o_2 _4329_ (.A1(_1111_),
    .A2(_1113_),
    .B1(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__nand3_1 _4330_ (.A(_1111_),
    .B(_1113_),
    .C(_1149_),
    .Y(_1151_));
 sky130_fd_sc_hd__and2_1 _4331_ (.A(_1150_),
    .B(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a22oi_1 _4332_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1118_),
    .B1(_1152_),
    .B2(net41),
    .Y(_1153_));
 sky130_fd_sc_hd__o21ai_1 _4333_ (.A1(_0670_),
    .A2(_1116_),
    .B1(_1153_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_2 _4334_ (.A(net252),
    .B(net178),
    .Y(_1154_));
 sky130_fd_sc_hd__xor2_1 _4335_ (.A(_1121_),
    .B(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__and3_1 _4336_ (.A(net249),
    .B(net180),
    .C(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a21oi_1 _4337_ (.A1(net249),
    .A2(net181),
    .B1(_1155_),
    .Y(_1157_));
 sky130_fd_sc_hd__nor2_1 _4338_ (.A(_1156_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__o21bai_2 _4339_ (.A1(_1091_),
    .A2(_1122_),
    .B1_N(_1124_),
    .Y(_1159_));
 sky130_fd_sc_hd__xnor2_1 _4340_ (.A(_1158_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__a22o_1 _4341_ (.A1(net240),
    .A2(net184),
    .B1(net182),
    .B2(net244),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_4 _4342_ (.A(net240),
    .B(net182),
    .Y(_1162_));
 sky130_fd_sc_hd__nor2_1 _4343_ (.A(_1130_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__o21ai_2 _4344_ (.A1(_1130_),
    .A2(_1162_),
    .B1(_1161_),
    .Y(_1164_));
 sky130_fd_sc_hd__xor2_1 _4345_ (.A(_1160_),
    .B(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__o21a_1 _4346_ (.A1(_1128_),
    .A2(_1135_),
    .B1(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__nor3_1 _4347_ (.A(_1128_),
    .B(_1135_),
    .C(_1165_),
    .Y(_1167_));
 sky130_fd_sc_hd__nor2_1 _4348_ (.A(_1166_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__o21ba_2 _4349_ (.A1(_1086_),
    .A2(_1130_),
    .B1_N(_1132_),
    .X(_1169_));
 sky130_fd_sc_hd__xnor2_2 _4350_ (.A(_1168_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__nor2_1 _4351_ (.A(_1138_),
    .B(_1140_),
    .Y(_1171_));
 sky130_fd_sc_hd__and2b_2 _4352_ (.A_N(_1171_),
    .B(_1170_),
    .X(_1172_));
 sky130_fd_sc_hd__xnor2_1 _4353_ (.A(_1170_),
    .B(_1171_),
    .Y(_1173_));
 sky130_fd_sc_hd__o21a_2 _4354_ (.A1(_1143_),
    .A2(_1145_),
    .B1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__nor3_1 _4355_ (.A(_1143_),
    .B(_1145_),
    .C(_1173_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_2 _4356_ (.A(_1174_),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__a21oi_4 _4357_ (.A1(_1148_),
    .A2(_1150_),
    .B1(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__and3_1 _4358_ (.A(_1148_),
    .B(_1150_),
    .C(_1176_),
    .X(_1178_));
 sky130_fd_sc_hd__nor2_1 _4359_ (.A(_1177_),
    .B(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__a22oi_1 _4360_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_1118_),
    .B1(_1179_),
    .B2(net41),
    .Y(_1180_));
 sky130_fd_sc_hd__o21ai_1 _4361_ (.A1(_0681_),
    .A2(_1116_),
    .B1(_1180_),
    .Y(_0108_));
 sky130_fd_sc_hd__nand2_4 _4362_ (.A(net249),
    .B(net188),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_2 _4363_ (.A(_1154_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__a22o_1 _4364_ (.A1(net252),
    .A2(net188),
    .B1(net178),
    .B2(net249),
    .X(_1183_));
 sky130_fd_sc_hd__o21a_1 _4365_ (.A1(_1154_),
    .A2(_1181_),
    .B1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__and3_2 _4366_ (.A(net244),
    .B(net180),
    .C(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__a21oi_2 _4367_ (.A1(net244),
    .A2(net180),
    .B1(_1184_),
    .Y(_1186_));
 sky130_fd_sc_hd__or2_4 _4368_ (.A(_1185_),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__o21ba_4 _4369_ (.A1(_1121_),
    .A2(_1154_),
    .B1_N(_1156_),
    .X(_1188_));
 sky130_fd_sc_hd__xnor2_4 _4370_ (.A(_1187_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__xnor2_2 _4371_ (.A(_1162_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__o2bb2a_1 _4372_ (.A1_N(_1158_),
    .A2_N(_1159_),
    .B1(_1160_),
    .B2(_1164_),
    .X(_1191_));
 sky130_fd_sc_hd__xor2_1 _4373_ (.A(_1190_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _4374_ (.A(_1163_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__or2_1 _4375_ (.A(_1163_),
    .B(_1192_),
    .X(_1194_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__o21ba_1 _4377_ (.A1(_1167_),
    .A2(_1169_),
    .B1_N(_1166_),
    .X(_1196_));
 sky130_fd_sc_hd__or2_1 _4378_ (.A(_1195_),
    .B(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__nand2_1 _4379_ (.A(_1195_),
    .B(_1196_),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nor2_1 _4382_ (.A(_1172_),
    .B(_1174_),
    .Y(_1201_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(_1201_),
    .A1(_1172_),
    .S(_1177_),
    .X(_1202_));
 sky130_fd_sc_hd__xnor2_1 _4384_ (.A(_1200_),
    .B(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__a22oi_1 _4385_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_1118_),
    .B1(_1203_),
    .B2(net41),
    .Y(_1204_));
 sky130_fd_sc_hd__o21ai_1 _4386_ (.A1(_0692_),
    .A2(_1116_),
    .B1(_1204_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_2 _4387_ (.A(net244),
    .B(net178),
    .Y(_1205_));
 sky130_fd_sc_hd__xor2_1 _4388_ (.A(_1181_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__and3_1 _4389_ (.A(net240),
    .B(net180),
    .C(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__a21oi_1 _4390_ (.A1(net240),
    .A2(net180),
    .B1(_1206_),
    .Y(_1208_));
 sky130_fd_sc_hd__nor2_2 _4391_ (.A(_1207_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__o21ai_4 _4392_ (.A1(_1182_),
    .A2(_1185_),
    .B1(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__or3_1 _4393_ (.A(_1182_),
    .B(_1185_),
    .C(_1209_),
    .X(_1211_));
 sky130_fd_sc_hd__nand2_2 _4394_ (.A(_1210_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__o32a_4 _4395_ (.A1(_1185_),
    .A2(_1186_),
    .A3(_1188_),
    .B1(_1189_),
    .B2(_1162_),
    .X(_1213_));
 sky130_fd_sc_hd__xor2_2 _4396_ (.A(_1212_),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__o21a_1 _4397_ (.A1(_1190_),
    .A2(_1191_),
    .B1(_1193_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2b_1 _4398_ (.A_N(_1215_),
    .B(_1214_),
    .Y(_1216_));
 sky130_fd_sc_hd__xor2_1 _4399_ (.A(_1214_),
    .B(_1215_),
    .X(_1217_));
 sky130_fd_sc_hd__nor2_1 _4400_ (.A(_1197_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__and2_1 _4401_ (.A(_1197_),
    .B(_1217_),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_1 _4402_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__o31ai_2 _4403_ (.A1(_1172_),
    .A2(_1174_),
    .A3(_1177_),
    .B1(_1200_),
    .Y(_1221_));
 sky130_fd_sc_hd__o311a_1 _4404_ (.A1(_1172_),
    .A2(_1174_),
    .A3(_1177_),
    .B1(_1200_),
    .C1(_1220_),
    .X(_1222_));
 sky130_fd_sc_hd__xnor2_1 _4405_ (.A(_1220_),
    .B(_1221_),
    .Y(_1223_));
 sky130_fd_sc_hd__a22oi_1 _4406_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1118_),
    .B1(_1223_),
    .B2(net41),
    .Y(_1224_));
 sky130_fd_sc_hd__o21ai_1 _4407_ (.A1(_0703_),
    .A2(_1116_),
    .B1(_1224_),
    .Y(_0110_));
 sky130_fd_sc_hd__o21bai_4 _4408_ (.A1(_1181_),
    .A2(_1205_),
    .B1_N(_1207_),
    .Y(_1225_));
 sky130_fd_sc_hd__a22oi_4 _4409_ (.A1(net244),
    .A2(net188),
    .B1(net178),
    .B2(net240),
    .Y(_1226_));
 sky130_fd_sc_hd__and4_1 _4410_ (.A(net240),
    .B(net244),
    .C(net188),
    .D(net178),
    .X(_1227_));
 sky130_fd_sc_hd__nor2_4 _4411_ (.A(_1226_),
    .B(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(_1225_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__xnor2_4 _4413_ (.A(_1225_),
    .B(_1228_),
    .Y(_1230_));
 sky130_fd_sc_hd__o21ai_2 _4414_ (.A1(_1212_),
    .A2(_1213_),
    .B1(_1210_),
    .Y(_1231_));
 sky130_fd_sc_hd__xnor2_2 _4415_ (.A(_1230_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2b_1 _4416_ (.A_N(_1216_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__xnor2_1 _4417_ (.A(_1216_),
    .B(_1232_),
    .Y(_1234_));
 sky130_fd_sc_hd__o21ai_2 _4418_ (.A1(_1218_),
    .A2(_1222_),
    .B1(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__or3_1 _4419_ (.A(_1218_),
    .B(_1222_),
    .C(_1234_),
    .X(_1236_));
 sky130_fd_sc_hd__and2_1 _4420_ (.A(_1235_),
    .B(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__a22oi_1 _4421_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_1118_),
    .B1(_1237_),
    .B2(net41),
    .Y(_1238_));
 sky130_fd_sc_hd__o21ai_1 _4422_ (.A1(_0714_),
    .A2(_1116_),
    .B1(_1238_),
    .Y(_0111_));
 sky130_fd_sc_hd__a2bb2o_1 _4423_ (.A1_N(_0724_),
    .A2_N(_1116_),
    .B1(_1118_),
    .B2(\as2650.r123_2[2][6] ),
    .X(_1239_));
 sky130_fd_sc_hd__or3_4 _4424_ (.A(_1212_),
    .B(_1213_),
    .C(_1230_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(net240),
    .B(net188),
    .Y(_1241_));
 sky130_fd_sc_hd__and3_2 _4426_ (.A(net240),
    .B(net188),
    .C(_1205_),
    .X(_1242_));
 sky130_fd_sc_hd__o21ai_4 _4427_ (.A1(_1210_),
    .A2(_1230_),
    .B1(_1229_),
    .Y(_1243_));
 sky130_fd_sc_hd__xnor2_4 _4428_ (.A(_1242_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__xnor2_1 _4429_ (.A(_1240_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__a21o_1 _4430_ (.A1(_1233_),
    .A2(_1235_),
    .B1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__nand3_1 _4431_ (.A(_1233_),
    .B(_1235_),
    .C(_1245_),
    .Y(_1247_));
 sky130_fd_sc_hd__and2_1 _4432_ (.A(_1246_),
    .B(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__a21o_1 _4433_ (.A1(net41),
    .A2(_1248_),
    .B1(_1239_),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _4434_ (.A1(_0735_),
    .A2(_1117_),
    .B1(_1118_),
    .B2(\as2650.r123_2[2][7] ),
    .X(_1249_));
 sky130_fd_sc_hd__a21oi_2 _4435_ (.A1(net244),
    .A2(net178),
    .B1(_1243_),
    .Y(_1250_));
 sky130_fd_sc_hd__o221ai_4 _4436_ (.A1(_1240_),
    .A2(_1244_),
    .B1(_1250_),
    .B2(_1241_),
    .C1(_1246_),
    .Y(_1251_));
 sky130_fd_sc_hd__a21o_1 _4437_ (.A1(net41),
    .A2(_1251_),
    .B1(_1249_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(net288),
    .A1(\as2650.stack[4][0] ),
    .S(_0784_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(net265),
    .A1(_1252_),
    .S(_0781_),
    .X(_0114_));
 sky130_fd_sc_hd__or2_1 _4440_ (.A(\as2650.stack[4][1] ),
    .B(_0783_),
    .X(_1253_));
 sky130_fd_sc_hd__o21a_1 _4441_ (.A1(net285),
    .A2(_0784_),
    .B1(_0781_),
    .X(_1254_));
 sky130_fd_sc_hd__a22o_1 _4442_ (.A1(net261),
    .A2(_0780_),
    .B1(_1253_),
    .B2(_1254_),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _4443_ (.A(\as2650.stack[4][2] ),
    .B(_0783_),
    .X(_1255_));
 sky130_fd_sc_hd__a21oi_1 _4444_ (.A1(_2634_),
    .A2(_0783_),
    .B1(_0780_),
    .Y(_1256_));
 sky130_fd_sc_hd__a22o_1 _4445_ (.A1(net257),
    .A2(_0780_),
    .B1(_1255_),
    .B2(_1256_),
    .X(_0116_));
 sky130_fd_sc_hd__or2_1 _4446_ (.A(\as2650.stack[4][3] ),
    .B(_0783_),
    .X(_1257_));
 sky130_fd_sc_hd__a21oi_1 _4447_ (.A1(_2633_),
    .A2(_0783_),
    .B1(_0780_),
    .Y(_1258_));
 sky130_fd_sc_hd__a22o_1 _4448_ (.A1(net254),
    .A2(_0780_),
    .B1(_1257_),
    .B2(_1258_),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _4449_ (.A(\as2650.stack[4][4] ),
    .B(_0783_),
    .X(_1259_));
 sky130_fd_sc_hd__a21oi_1 _4450_ (.A1(_2632_),
    .A2(_0783_),
    .B1(_0780_),
    .Y(_1260_));
 sky130_fd_sc_hd__a22o_1 _4451_ (.A1(net251),
    .A2(_0780_),
    .B1(_1259_),
    .B2(_1260_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_1 _4452_ (.A(\as2650.stack[4][5] ),
    .B(_0783_),
    .X(_1261_));
 sky130_fd_sc_hd__o21a_1 _4453_ (.A1(net280),
    .A2(_0784_),
    .B1(_0781_),
    .X(_1262_));
 sky130_fd_sc_hd__a22o_1 _4454_ (.A1(net247),
    .A2(_0780_),
    .B1(_1261_),
    .B2(_1262_),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _4455_ (.A(\as2650.stack[4][6] ),
    .B(_0783_),
    .X(_1263_));
 sky130_fd_sc_hd__o21a_1 _4456_ (.A1(net277),
    .A2(_0784_),
    .B1(_0781_),
    .X(_1264_));
 sky130_fd_sc_hd__a22o_1 _4457_ (.A1(net243),
    .A2(_0780_),
    .B1(_1263_),
    .B2(_1264_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _4458_ (.A(\as2650.stack[4][7] ),
    .B(_0783_),
    .X(_1265_));
 sky130_fd_sc_hd__o21a_1 _4459_ (.A1(net275),
    .A2(_0784_),
    .B1(_0781_),
    .X(_1266_));
 sky130_fd_sc_hd__a22o_1 _4460_ (.A1(net239),
    .A2(_0780_),
    .B1(_1265_),
    .B2(_1266_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4461_ (.A0(net286),
    .A1(\as2650.stack[2][0] ),
    .S(_0907_),
    .X(_1267_));
 sky130_fd_sc_hd__or3_4 _4462_ (.A(net206),
    .B(_0591_),
    .C(_0897_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(net265),
    .A1(_1267_),
    .S(_0898_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(net284),
    .A1(\as2650.stack[2][1] ),
    .S(_0907_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(net261),
    .A1(_1269_),
    .S(_0898_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(\as2650.pc[2] ),
    .A1(\as2650.stack[2][2] ),
    .S(_0907_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(net257),
    .A1(_1270_),
    .S(_1268_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(net283),
    .A1(\as2650.stack[2][3] ),
    .S(_0907_),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(net254),
    .A1(_1271_),
    .S(_1268_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(net281),
    .A1(\as2650.stack[2][4] ),
    .S(_0907_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(net251),
    .A1(_1272_),
    .S(_0898_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(net280),
    .A1(\as2650.stack[2][5] ),
    .S(_0907_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(net247),
    .A1(_1273_),
    .S(_0898_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(net277),
    .A1(\as2650.stack[2][6] ),
    .S(_0907_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(net243),
    .A1(_1274_),
    .S(_0898_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(net275),
    .A1(\as2650.stack[2][7] ),
    .S(_0907_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(net239),
    .A1(_1275_),
    .S(_1268_),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _4478_ (.A(\as2650.stack[1][0] ),
    .B(_1071_),
    .X(_1276_));
 sky130_fd_sc_hd__a21oi_1 _4479_ (.A1(_2635_),
    .A2(net48),
    .B1(_0908_),
    .Y(_1277_));
 sky130_fd_sc_hd__a22o_1 _4480_ (.A1(net265),
    .A2(_0908_),
    .B1(_1276_),
    .B2(_1277_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_1 _4481_ (.A(\as2650.stack[1][1] ),
    .B(net48),
    .X(_1278_));
 sky130_fd_sc_hd__o21a_1 _4482_ (.A1(net284),
    .A2(_1072_),
    .B1(_0909_),
    .X(_1279_));
 sky130_fd_sc_hd__a22o_1 _4483_ (.A1(net261),
    .A2(net51),
    .B1(_1278_),
    .B2(_1279_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _4484_ (.A(\as2650.stack[1][2] ),
    .B(net48),
    .X(_1280_));
 sky130_fd_sc_hd__a21oi_1 _4485_ (.A1(_2634_),
    .A2(net48),
    .B1(net51),
    .Y(_1281_));
 sky130_fd_sc_hd__a22o_1 _4486_ (.A1(net257),
    .A2(net51),
    .B1(_1280_),
    .B2(_1281_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _4487_ (.A(\as2650.stack[1][3] ),
    .B(net48),
    .X(_1282_));
 sky130_fd_sc_hd__a21oi_1 _4488_ (.A1(_2633_),
    .A2(net48),
    .B1(net51),
    .Y(_1283_));
 sky130_fd_sc_hd__a22o_1 _4489_ (.A1(net254),
    .A2(net51),
    .B1(_1282_),
    .B2(_1283_),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _4490_ (.A(\as2650.stack[1][4] ),
    .B(_1071_),
    .X(_1284_));
 sky130_fd_sc_hd__a21oi_1 _4491_ (.A1(_2632_),
    .A2(net48),
    .B1(net51),
    .Y(_1285_));
 sky130_fd_sc_hd__a22o_1 _4492_ (.A1(net251),
    .A2(net51),
    .B1(_1284_),
    .B2(_1285_),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _4493_ (.A(\as2650.stack[1][5] ),
    .B(net48),
    .X(_1286_));
 sky130_fd_sc_hd__o21a_1 _4494_ (.A1(net279),
    .A2(_1072_),
    .B1(_0909_),
    .X(_1287_));
 sky130_fd_sc_hd__a22o_1 _4495_ (.A1(net247),
    .A2(net51),
    .B1(_1286_),
    .B2(_1287_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _4496_ (.A(\as2650.stack[1][6] ),
    .B(net48),
    .X(_1288_));
 sky130_fd_sc_hd__o21a_1 _4497_ (.A1(net278),
    .A2(_1072_),
    .B1(_0909_),
    .X(_1289_));
 sky130_fd_sc_hd__a22o_1 _4498_ (.A1(net243),
    .A2(net51),
    .B1(_1288_),
    .B2(_1289_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _4499_ (.A(\as2650.stack[1][7] ),
    .B(net48),
    .X(_1290_));
 sky130_fd_sc_hd__o21a_1 _4500_ (.A1(net275),
    .A2(_1072_),
    .B1(_0909_),
    .X(_1291_));
 sky130_fd_sc_hd__a22o_1 _4501_ (.A1(net239),
    .A2(net51),
    .B1(_1290_),
    .B2(_1291_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(net286),
    .A1(\as2650.stack[3][0] ),
    .S(_0900_),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(net265),
    .A1(_1292_),
    .S(_0786_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(net284),
    .A1(\as2650.stack[3][1] ),
    .S(_0900_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(net261),
    .A1(_1293_),
    .S(_0786_),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _4506_ (.A(\as2650.stack[3][2] ),
    .B(_0899_),
    .X(_1294_));
 sky130_fd_sc_hd__a21oi_1 _4507_ (.A1(_2634_),
    .A2(_0899_),
    .B1(_0785_),
    .Y(_1295_));
 sky130_fd_sc_hd__a22o_1 _4508_ (.A1(net257),
    .A2(_0785_),
    .B1(_1294_),
    .B2(_1295_),
    .X(_0148_));
 sky130_fd_sc_hd__or2_1 _4509_ (.A(\as2650.stack[3][3] ),
    .B(_0899_),
    .X(_1296_));
 sky130_fd_sc_hd__a21oi_1 _4510_ (.A1(_2633_),
    .A2(_0899_),
    .B1(_0785_),
    .Y(_1297_));
 sky130_fd_sc_hd__a22o_1 _4511_ (.A1(net254),
    .A2(_0785_),
    .B1(_1296_),
    .B2(_1297_),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _4512_ (.A(\as2650.stack[3][4] ),
    .B(_0899_),
    .X(_1298_));
 sky130_fd_sc_hd__a21oi_1 _4513_ (.A1(_2632_),
    .A2(_0899_),
    .B1(_0785_),
    .Y(_1299_));
 sky130_fd_sc_hd__a22o_1 _4514_ (.A1(net251),
    .A2(_0785_),
    .B1(_1298_),
    .B2(_1299_),
    .X(_0150_));
 sky130_fd_sc_hd__or2_1 _4515_ (.A(\as2650.stack[3][5] ),
    .B(_0899_),
    .X(_1300_));
 sky130_fd_sc_hd__o21a_1 _4516_ (.A1(net279),
    .A2(_0900_),
    .B1(_0786_),
    .X(_1301_));
 sky130_fd_sc_hd__a22o_1 _4517_ (.A1(net247),
    .A2(_0785_),
    .B1(_1300_),
    .B2(_1301_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(net277),
    .A1(\as2650.stack[3][6] ),
    .S(_0900_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(net243),
    .A1(_1302_),
    .S(_0786_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(net275),
    .A1(\as2650.stack[3][7] ),
    .S(_0900_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(net239),
    .A1(_1303_),
    .S(_0786_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _4522_ (.A(net318),
    .B(\lfsr[1] ),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _4523_ (.A(net324),
    .B(\lfsr[2] ),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _4524_ (.A(net318),
    .B(\lfsr[3] ),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _4525_ (.A(net324),
    .B(\lfsr[4] ),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _4526_ (.A(net318),
    .B(\as2650.sense ),
    .X(_0158_));
 sky130_fd_sc_hd__or2_1 _4527_ (.A(net324),
    .B(\lfsr[6] ),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _4528_ (.A(net318),
    .B(\lfsr[7] ),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _4529_ (.A(net324),
    .B(\lfsr[8] ),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _4530_ (.A(net318),
    .B(\lfsr[9] ),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _4531_ (.A(net325),
    .B(\lfsr[10] ),
    .X(_0163_));
 sky130_fd_sc_hd__a21oi_1 _4532_ (.A1(\lfsr[0] ),
    .A2(\lfsr[11] ),
    .B1(net324),
    .Y(_1304_));
 sky130_fd_sc_hd__o21a_1 _4533_ (.A1(\lfsr[0] ),
    .A2(\lfsr[11] ),
    .B1(_1304_),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _4534_ (.A(net324),
    .B(\lfsr[12] ),
    .X(_0165_));
 sky130_fd_sc_hd__a21oi_1 _4535_ (.A1(\lfsr[0] ),
    .A2(\lfsr[13] ),
    .B1(net324),
    .Y(_1305_));
 sky130_fd_sc_hd__o21a_1 _4536_ (.A1(\lfsr[0] ),
    .A2(\lfsr[13] ),
    .B1(_1305_),
    .X(_0166_));
 sky130_fd_sc_hd__a21oi_1 _4537_ (.A1(_2663_),
    .A2(\lfsr[14] ),
    .B1(net324),
    .Y(_1306_));
 sky130_fd_sc_hd__o21ai_1 _4538_ (.A1(_2663_),
    .A2(\lfsr[14] ),
    .B1(_1306_),
    .Y(_0167_));
 sky130_fd_sc_hd__and2_1 _4539_ (.A(net318),
    .B(\lfsr[15] ),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _4540_ (.A(net324),
    .B(\lfsr[0] ),
    .X(_0169_));
 sky130_fd_sc_hd__or2_1 _4541_ (.A(\as2650.stack[0][0] ),
    .B(net47),
    .X(_1307_));
 sky130_fd_sc_hd__a21oi_1 _4542_ (.A1(_2635_),
    .A2(net47),
    .B1(net50),
    .Y(_1308_));
 sky130_fd_sc_hd__a22o_1 _4543_ (.A1(net265),
    .A2(net50),
    .B1(_1307_),
    .B2(_1308_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _4544_ (.A(\as2650.stack[0][1] ),
    .B(net47),
    .X(_1309_));
 sky130_fd_sc_hd__o21a_1 _4545_ (.A1(net284),
    .A2(_1078_),
    .B1(_1074_),
    .X(_1310_));
 sky130_fd_sc_hd__a22o_1 _4546_ (.A1(net261),
    .A2(net50),
    .B1(_1309_),
    .B2(_1310_),
    .X(_0171_));
 sky130_fd_sc_hd__or2_1 _4547_ (.A(\as2650.stack[0][2] ),
    .B(net47),
    .X(_1311_));
 sky130_fd_sc_hd__a21oi_1 _4548_ (.A1(_2634_),
    .A2(net47),
    .B1(net50),
    .Y(_1312_));
 sky130_fd_sc_hd__a22o_1 _4549_ (.A1(net257),
    .A2(net50),
    .B1(_1311_),
    .B2(_1312_),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _4550_ (.A(\as2650.stack[0][3] ),
    .B(_1077_),
    .X(_1313_));
 sky130_fd_sc_hd__a21oi_1 _4551_ (.A1(_2633_),
    .A2(net47),
    .B1(_1073_),
    .Y(_1314_));
 sky130_fd_sc_hd__a22o_1 _4552_ (.A1(net254),
    .A2(_1073_),
    .B1(_1313_),
    .B2(_1314_),
    .X(_0173_));
 sky130_fd_sc_hd__or2_1 _4553_ (.A(\as2650.stack[0][4] ),
    .B(_1077_),
    .X(_1315_));
 sky130_fd_sc_hd__a21oi_1 _4554_ (.A1(_2632_),
    .A2(net47),
    .B1(net50),
    .Y(_1316_));
 sky130_fd_sc_hd__a22o_1 _4555_ (.A1(net251),
    .A2(net50),
    .B1(_1315_),
    .B2(_1316_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _4556_ (.A(\as2650.stack[0][5] ),
    .B(net47),
    .X(_1317_));
 sky130_fd_sc_hd__o21a_1 _4557_ (.A1(net279),
    .A2(_1078_),
    .B1(_1074_),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _4558_ (.A1(net247),
    .A2(net50),
    .B1(_1317_),
    .B2(_1318_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _4559_ (.A(\as2650.stack[0][6] ),
    .B(net47),
    .X(_1319_));
 sky130_fd_sc_hd__o21a_1 _4560_ (.A1(net278),
    .A2(_1078_),
    .B1(_1074_),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_1 _4561_ (.A1(net243),
    .A2(net50),
    .B1(_1319_),
    .B2(_1320_),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _4562_ (.A(\as2650.stack[0][7] ),
    .B(net47),
    .X(_1321_));
 sky130_fd_sc_hd__o21a_1 _4563_ (.A1(net275),
    .A2(_1078_),
    .B1(_1074_),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_1 _4564_ (.A1(net239),
    .A2(net50),
    .B1(_1321_),
    .B2(_1322_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_2 _4565_ (.A(net154),
    .B(net81),
    .Y(_1323_));
 sky130_fd_sc_hd__and3b_1 _4566_ (.A_N(_2734_),
    .B(_2795_),
    .C(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_2 _4567_ (.A(net294),
    .B(net173),
    .Y(_1325_));
 sky130_fd_sc_hd__and3_1 _4568_ (.A(_2688_),
    .B(_2765_),
    .C(_0761_),
    .X(_1326_));
 sky130_fd_sc_hd__or3b_1 _4569_ (.A(net163),
    .B(_1326_),
    .C_N(_1325_),
    .X(_1327_));
 sky130_fd_sc_hd__o32a_1 _4570_ (.A1(net148),
    .A2(_2698_),
    .A3(_0837_),
    .B1(_0836_),
    .B2(net87),
    .X(_1328_));
 sky130_fd_sc_hd__a21oi_1 _4571_ (.A1(net171),
    .A2(_0746_),
    .B1(net59),
    .Y(_1329_));
 sky130_fd_sc_hd__and3b_1 _4572_ (.A_N(_1327_),
    .B(_1328_),
    .C(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__o211a_2 _4573_ (.A1(_2686_),
    .A2(_0834_),
    .B1(_1324_),
    .C1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__a22o_1 _4574_ (.A1(net230),
    .A2(net161),
    .B1(_2729_),
    .B2(net217),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(net26),
    .A1(_1332_),
    .S(_1331_),
    .X(_1333_));
 sky130_fd_sc_hd__and2_1 _4576_ (.A(net317),
    .B(_1333_),
    .X(_0178_));
 sky130_fd_sc_hd__or4_1 _4577_ (.A(net236),
    .B(net132),
    .C(_2790_),
    .D(_0843_),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_1 _4578_ (.A0(net298),
    .A1(net28),
    .S(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__and2_1 _4579_ (.A(net316),
    .B(_1335_),
    .X(_0179_));
 sky130_fd_sc_hd__or3_1 _4580_ (.A(_2668_),
    .B(net154),
    .C(_0837_),
    .X(_1336_));
 sky130_fd_sc_hd__o221a_2 _4581_ (.A1(_2726_),
    .A2(net103),
    .B1(_0837_),
    .B2(net159),
    .C1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a21oi_1 _4582_ (.A1(net141),
    .A2(net126),
    .B1(_2794_),
    .Y(_1338_));
 sky130_fd_sc_hd__o221a_2 _4583_ (.A1(_0747_),
    .A2(_0760_),
    .B1(_1338_),
    .B2(_2731_),
    .C1(_1337_),
    .X(_1339_));
 sky130_fd_sc_hd__a21boi_1 _4584_ (.A1(_0842_),
    .A2(_1339_),
    .B1_N(net27),
    .Y(_1340_));
 sky130_fd_sc_hd__a311o_1 _4585_ (.A1(_2703_),
    .A2(_0842_),
    .A3(_1339_),
    .B1(_1340_),
    .C1(net322),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_4 _4586_ (.A(net132),
    .B(_0814_),
    .Y(_1341_));
 sky130_fd_sc_hd__or4_4 _4587_ (.A(net95),
    .B(_2794_),
    .C(_0747_),
    .D(net70),
    .X(_1342_));
 sky130_fd_sc_hd__or2_4 _4588_ (.A(net229),
    .B(_2726_),
    .X(_1343_));
 sky130_fd_sc_hd__inv_2 _4589_ (.A(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__or4b_4 _4590_ (.A(net87),
    .B(net198),
    .C(_0823_),
    .D_N(_0826_),
    .X(_1345_));
 sky130_fd_sc_hd__o22ai_2 _4591_ (.A1(_2726_),
    .A2(_1342_),
    .B1(_1343_),
    .B2(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__or2_1 _4592_ (.A(_2722_),
    .B(_2782_),
    .X(_1347_));
 sky130_fd_sc_hd__xnor2_2 _4593_ (.A(net291),
    .B(net293),
    .Y(_1348_));
 sky130_fd_sc_hd__nor2_1 _4594_ (.A(_2805_),
    .B(_0743_),
    .Y(_1349_));
 sky130_fd_sc_hd__a31o_2 _4595_ (.A1(net233),
    .A2(_2672_),
    .A3(_0742_),
    .B1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__and4_2 _4596_ (.A(net172),
    .B(_2728_),
    .C(net129),
    .D(_2826_),
    .X(_1351_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_1350_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__o41a_1 _4598_ (.A1(net96),
    .A2(_2727_),
    .A3(_2739_),
    .A4(_1347_),
    .B1(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__a21o_1 _4599_ (.A1(net73),
    .A2(net125),
    .B1(net88),
    .X(_1354_));
 sky130_fd_sc_hd__nor2_1 _4600_ (.A(net212),
    .B(_2731_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_4 _4601_ (.A(net229),
    .B(net129),
    .Y(_1356_));
 sky130_fd_sc_hd__a21oi_2 _4602_ (.A1(_2669_),
    .A2(_2696_),
    .B1(net294),
    .Y(_1357_));
 sky130_fd_sc_hd__inv_2 _4603_ (.A(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__or4_1 _4604_ (.A(net87),
    .B(_2789_),
    .C(net125),
    .D(net163),
    .X(_1359_));
 sky130_fd_sc_hd__and4_1 _4605_ (.A(_2733_),
    .B(_1323_),
    .C(_1354_),
    .D(_1357_),
    .X(_1360_));
 sky130_fd_sc_hd__o31a_2 _4606_ (.A1(net305),
    .A2(net88),
    .A3(_0752_),
    .B1(_0587_),
    .X(_1361_));
 sky130_fd_sc_hd__o21a_1 _4607_ (.A1(_0817_),
    .A2(_0823_),
    .B1(net96),
    .X(_1362_));
 sky130_fd_sc_hd__and3_1 _4608_ (.A(net305),
    .B(net95),
    .C(_0751_),
    .X(_1363_));
 sky130_fd_sc_hd__a21oi_2 _4609_ (.A1(net95),
    .A2(_0755_),
    .B1(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__o21a_1 _4610_ (.A1(_2726_),
    .A2(_2776_),
    .B1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__o21a_1 _4611_ (.A1(net128),
    .A2(_0760_),
    .B1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nor3_1 _4612_ (.A(net210),
    .B(_2706_),
    .C(_2726_),
    .Y(_1367_));
 sky130_fd_sc_hd__o221a_1 _4613_ (.A1(_2790_),
    .A2(_0760_),
    .B1(net103),
    .B2(_2726_),
    .C1(_2730_),
    .X(_1368_));
 sky130_fd_sc_hd__or2_4 _4614_ (.A(_2815_),
    .B(_2865_),
    .X(_1369_));
 sky130_fd_sc_hd__nor3_1 _4615_ (.A(_0758_),
    .B(_0817_),
    .C(_0823_),
    .Y(_1370_));
 sky130_fd_sc_hd__o2111a_1 _4616_ (.A1(net87),
    .A2(_1370_),
    .B1(_1369_),
    .C1(_1368_),
    .D1(_0587_),
    .X(_1371_));
 sky130_fd_sc_hd__nand3_1 _4617_ (.A(_1353_),
    .B(_1366_),
    .C(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__or4b_4 _4618_ (.A(_1346_),
    .B(_1367_),
    .C(_1372_),
    .D_N(_1360_),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_1 _4619_ (.A(_2947_),
    .B(_0344_),
    .Y(_1374_));
 sky130_fd_sc_hd__and4_1 _4620_ (.A(_2881_),
    .B(_3000_),
    .C(_0506_),
    .D(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__and4b_4 _4621_ (.A_N(_0402_),
    .B(_0455_),
    .C(_0540_),
    .D(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__and3_2 _4622_ (.A(net232),
    .B(net298),
    .C(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_4 _4623_ (.A(_1351_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_8 _4624_ (.A(_0829_),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__nor2_1 _4625_ (.A(_1373_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a21oi_2 _4626_ (.A1(_2819_),
    .A2(_2906_),
    .B1(_2651_),
    .Y(_1381_));
 sky130_fd_sc_hd__a31o_1 _4627_ (.A1(_2651_),
    .A2(_2819_),
    .A3(_2906_),
    .B1(net83),
    .X(_1382_));
 sky130_fd_sc_hd__and3_1 _4628_ (.A(net347),
    .B(net196),
    .C(_2912_),
    .X(_1383_));
 sky130_fd_sc_hd__a21oi_1 _4629_ (.A1(net196),
    .A2(_2912_),
    .B1(net347),
    .Y(_1384_));
 sky130_fd_sc_hd__o21ai_2 _4630_ (.A1(_1383_),
    .A2(_1384_),
    .B1(_2718_),
    .Y(_1385_));
 sky130_fd_sc_hd__o21ai_4 _4631_ (.A1(_1381_),
    .A2(_1382_),
    .B1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_2 _4632_ (.A(net286),
    .B(net349),
    .Y(_1387_));
 sky130_fd_sc_hd__or2_1 _4633_ (.A(net286),
    .B(net349),
    .X(_1388_));
 sky130_fd_sc_hd__and2_2 _4634_ (.A(_1387_),
    .B(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__a221o_1 _4635_ (.A1(net36),
    .A2(net131),
    .B1(net79),
    .B2(_1389_),
    .C1(net80),
    .X(_1390_));
 sky130_fd_sc_hd__a21oi_1 _4636_ (.A1(_2720_),
    .A2(_1386_),
    .B1(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(net36),
    .A1(_1389_),
    .S(net327),
    .X(_1392_));
 sky130_fd_sc_hd__nor2_4 _4638_ (.A(net215),
    .B(net137),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_8 _4639_ (.A(net238),
    .B(net132),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _4640_ (.A(_2744_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__and2_4 _4641_ (.A(net301),
    .B(net160),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_4 _4642_ (.A(net303),
    .B(net160),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_1 _4643_ (.A(net132),
    .B(net63),
    .Y(_1398_));
 sky130_fd_sc_hd__nor2_4 _4644_ (.A(_1394_),
    .B(_1396_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _4645_ (.A(net64),
    .B(net63),
    .Y(_1400_));
 sky130_fd_sc_hd__nor2_4 _4646_ (.A(net160),
    .B(net146),
    .Y(_1401_));
 sky130_fd_sc_hd__nand2_1 _4647_ (.A(net36),
    .B(_0574_),
    .Y(_1402_));
 sky130_fd_sc_hd__nor2_8 _4648_ (.A(_2648_),
    .B(net149),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_8 _4649_ (.A(net309),
    .B(net153),
    .Y(_1404_));
 sky130_fd_sc_hd__o221a_1 _4650_ (.A1(net36),
    .A2(net148),
    .B1(_1404_),
    .B2(_2651_),
    .C1(_1401_),
    .X(_1405_));
 sky130_fd_sc_hd__o2bb2a_1 _4651_ (.A1_N(_1402_),
    .A2_N(_1405_),
    .B1(_2744_),
    .B2(_1392_),
    .X(_1406_));
 sky130_fd_sc_hd__o221a_1 _4652_ (.A1(net286),
    .A2(_1399_),
    .B1(_1406_),
    .B2(_1394_),
    .C1(net229),
    .X(_1407_));
 sky130_fd_sc_hd__o21a_1 _4653_ (.A1(_1391_),
    .A2(_1407_),
    .B1(net129),
    .X(_1408_));
 sky130_fd_sc_hd__nor2_1 _4654_ (.A(_2731_),
    .B(net59),
    .Y(_1409_));
 sky130_fd_sc_hd__o21ai_1 _4655_ (.A1(_2635_),
    .A2(net52),
    .B1(net40),
    .Y(_1410_));
 sky130_fd_sc_hd__o221a_1 _4656_ (.A1(net36),
    .A2(net40),
    .B1(_1408_),
    .B2(_1410_),
    .C1(net316),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _4657_ (.A(net346),
    .B(_2962_),
    .X(_1411_));
 sky130_fd_sc_hd__xnor2_4 _4658_ (.A(_2652_),
    .B(_2962_),
    .Y(_1412_));
 sky130_fd_sc_hd__and2_2 _4659_ (.A(net347),
    .B(_2906_),
    .X(_1413_));
 sky130_fd_sc_hd__xor2_1 _4660_ (.A(_1412_),
    .B(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _4661_ (.A0(net2),
    .A1(_1414_),
    .S(_2819_),
    .X(_1415_));
 sky130_fd_sc_hd__and2_1 _4662_ (.A(net345),
    .B(_2965_),
    .X(_1416_));
 sky130_fd_sc_hd__or2_1 _4663_ (.A(net345),
    .B(_2965_),
    .X(_1417_));
 sky130_fd_sc_hd__nand2b_1 _4664_ (.A_N(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__and2_1 _4665_ (.A(net348),
    .B(_2912_),
    .X(_1419_));
 sky130_fd_sc_hd__xnor2_1 _4666_ (.A(_1418_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(net345),
    .A1(_1420_),
    .S(net196),
    .X(_1421_));
 sky130_fd_sc_hd__a22o_2 _4668_ (.A1(net86),
    .A2(_1415_),
    .B1(_1421_),
    .B2(_2718_),
    .X(_1422_));
 sky130_fd_sc_hd__xor2_1 _4669_ (.A(net37),
    .B(net36),
    .X(_1423_));
 sky130_fd_sc_hd__and2_1 _4670_ (.A(net284),
    .B(net345),
    .X(_1424_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(net284),
    .B(net345),
    .Y(_1425_));
 sky130_fd_sc_hd__nor2_1 _4672_ (.A(net284),
    .B(net345),
    .Y(_1426_));
 sky130_fd_sc_hd__nor2_2 _4673_ (.A(_1424_),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_1388_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__or2_1 _4675_ (.A(_1388_),
    .B(_1427_),
    .X(_1429_));
 sky130_fd_sc_hd__and3_1 _4676_ (.A(net78),
    .B(_1428_),
    .C(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__a221o_1 _4677_ (.A1(_2720_),
    .A2(_1422_),
    .B1(_1423_),
    .B2(net131),
    .C1(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__xnor2_2 _4678_ (.A(_1387_),
    .B(_1427_),
    .Y(_1432_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(net37),
    .A1(_1432_),
    .S(net327),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(net37),
    .A1(net345),
    .S(net309),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(_1423_),
    .A1(_1434_),
    .S(net148),
    .X(_1435_));
 sky130_fd_sc_hd__a22o_1 _4682_ (.A1(_2743_),
    .A2(_1433_),
    .B1(_1435_),
    .B2(_1401_),
    .X(_1436_));
 sky130_fd_sc_hd__a221o_1 _4683_ (.A1(net284),
    .A2(_1400_),
    .B1(_1436_),
    .B2(net64),
    .C1(net212),
    .X(_1437_));
 sky130_fd_sc_hd__o21ai_1 _4684_ (.A1(net80),
    .A2(_1431_),
    .B1(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__a2bb2o_1 _4685_ (.A1_N(net284),
    .A2_N(net52),
    .B1(_1438_),
    .B2(net129),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(net38),
    .B(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__o211a_1 _4687_ (.A1(net37),
    .A2(net39),
    .B1(_1440_),
    .C1(net314),
    .X(_0182_));
 sky130_fd_sc_hd__a21o_1 _4688_ (.A1(_1417_),
    .A2(_1419_),
    .B1(_1416_),
    .X(_1441_));
 sky130_fd_sc_hd__or2_2 _4689_ (.A(net342),
    .B(_0316_),
    .X(_1442_));
 sky130_fd_sc_hd__nand2_1 _4690_ (.A(net342),
    .B(_0316_),
    .Y(_1443_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_1442_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_1 _4692_ (.A(_1441_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21o_1 _4693_ (.A1(_1441_),
    .A2(_1444_),
    .B1(_2784_),
    .X(_1446_));
 sky130_fd_sc_hd__o22a_1 _4694_ (.A1(net342),
    .A2(net196),
    .B1(_1445_),
    .B2(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__a21o_1 _4695_ (.A1(_1412_),
    .A2(_1413_),
    .B1(_1411_),
    .X(_1448_));
 sky130_fd_sc_hd__or2_4 _4696_ (.A(net344),
    .B(_0312_),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _4697_ (.A(net344),
    .B(_0312_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_1449_),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__xnor2_1 _4699_ (.A(_1448_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(net344),
    .A1(_1452_),
    .S(_2819_),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_4 _4701_ (.A1(_2718_),
    .A2(_1447_),
    .B1(_1453_),
    .B2(net86),
    .X(_1454_));
 sky130_fd_sc_hd__and3_1 _4702_ (.A(net12),
    .B(net37),
    .C(net36),
    .X(_1455_));
 sky130_fd_sc_hd__a21oi_1 _4703_ (.A1(net37),
    .A2(net36),
    .B1(net12),
    .Y(_1456_));
 sky130_fd_sc_hd__or2_1 _4704_ (.A(_1455_),
    .B(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_2715_),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand2_2 _4706_ (.A(\as2650.pc[2] ),
    .B(net342),
    .Y(_1459_));
 sky130_fd_sc_hd__or2_1 _4707_ (.A(\as2650.pc[2] ),
    .B(net342),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_2 _4708_ (.A(_1459_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__a21o_1 _4709_ (.A1(_1425_),
    .A2(_1428_),
    .B1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nand3_1 _4710_ (.A(_1425_),
    .B(_1428_),
    .C(_1461_),
    .Y(_1463_));
 sky130_fd_sc_hd__a32o_1 _4711_ (.A1(net78),
    .A2(_1462_),
    .A3(_1463_),
    .B1(_1454_),
    .B2(_2720_),
    .X(_1464_));
 sky130_fd_sc_hd__o21a_1 _4712_ (.A1(_1387_),
    .A2(_1426_),
    .B1(_1425_),
    .X(_1465_));
 sky130_fd_sc_hd__xnor2_2 _4713_ (.A(_1461_),
    .B(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(net326),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__o211a_1 _4715_ (.A1(net12),
    .A2(net327),
    .B1(_2743_),
    .C1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__nand2_1 _4716_ (.A(net149),
    .B(_1457_),
    .Y(_1469_));
 sky130_fd_sc_hd__o22a_1 _4717_ (.A1(net12),
    .A2(_0575_),
    .B1(_1404_),
    .B2(net342),
    .X(_1470_));
 sky130_fd_sc_hd__a31o_1 _4718_ (.A1(_1401_),
    .A2(_1469_),
    .A3(_1470_),
    .B1(_1468_),
    .X(_1471_));
 sky130_fd_sc_hd__a221o_1 _4719_ (.A1(\as2650.pc[2] ),
    .A2(_1400_),
    .B1(_1471_),
    .B2(net64),
    .C1(net212),
    .X(_1472_));
 sky130_fd_sc_hd__o31a_1 _4720_ (.A1(net80),
    .A2(_1458_),
    .A3(_1464_),
    .B1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__or2_1 _4721_ (.A(net12),
    .B(net39),
    .X(_1474_));
 sky130_fd_sc_hd__o22a_1 _4722_ (.A1(\as2650.pc[2] ),
    .A2(net52),
    .B1(_1473_),
    .B2(net130),
    .X(_1475_));
 sky130_fd_sc_hd__o311a_1 _4723_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1475_),
    .B1(_1474_),
    .C1(net313),
    .X(_0183_));
 sky130_fd_sc_hd__nor2_1 _4724_ (.A(net340),
    .B(_0362_),
    .Y(_1476_));
 sky130_fd_sc_hd__or2_2 _4725_ (.A(net340),
    .B(_0362_),
    .X(_1477_));
 sky130_fd_sc_hd__and2_2 _4726_ (.A(net340),
    .B(_0362_),
    .X(_1478_));
 sky130_fd_sc_hd__nor2_1 _4727_ (.A(_1476_),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__a221o_4 _4728_ (.A1(net344),
    .A2(_0312_),
    .B1(_1412_),
    .B2(_1413_),
    .C1(_1411_),
    .X(_1480_));
 sky130_fd_sc_hd__a21oi_1 _4729_ (.A1(_1449_),
    .A2(_1480_),
    .B1(_1479_),
    .Y(_1481_));
 sky130_fd_sc_hd__a31o_1 _4730_ (.A1(_1449_),
    .A2(_1479_),
    .A3(_1480_),
    .B1(_2820_),
    .X(_1482_));
 sky130_fd_sc_hd__a2bb2o_1 _4731_ (.A1_N(_1481_),
    .A2_N(_1482_),
    .B1(net340),
    .B2(_2820_),
    .X(_1483_));
 sky130_fd_sc_hd__nor2_1 _4732_ (.A(net340),
    .B(_0364_),
    .Y(_1484_));
 sky130_fd_sc_hd__or2_1 _4733_ (.A(net341),
    .B(_0364_),
    .X(_1485_));
 sky130_fd_sc_hd__and2_1 _4734_ (.A(net340),
    .B(_0364_),
    .X(_1486_));
 sky130_fd_sc_hd__nor2_1 _4735_ (.A(_1484_),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__a221o_1 _4736_ (.A1(net343),
    .A2(_0316_),
    .B1(_1417_),
    .B2(_1419_),
    .C1(_1416_),
    .X(_1488_));
 sky130_fd_sc_hd__a21oi_1 _4737_ (.A1(_1442_),
    .A2(_1488_),
    .B1(_1487_),
    .Y(_1489_));
 sky130_fd_sc_hd__a31o_1 _4738_ (.A1(_1442_),
    .A2(_1487_),
    .A3(_1488_),
    .B1(_2784_),
    .X(_1490_));
 sky130_fd_sc_hd__o22a_1 _4739_ (.A1(_2654_),
    .A2(net196),
    .B1(_1489_),
    .B2(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a2bb2o_4 _4740_ (.A1_N(net83),
    .A2_N(_1483_),
    .B1(_1491_),
    .B2(_2718_),
    .X(_1492_));
 sky130_fd_sc_hd__and2_1 _4741_ (.A(net13),
    .B(_1455_),
    .X(_1493_));
 sky130_fd_sc_hd__nor2_1 _4742_ (.A(net13),
    .B(_1455_),
    .Y(_1494_));
 sky130_fd_sc_hd__or2_1 _4743_ (.A(_1493_),
    .B(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2_8 _4744_ (.A(\as2650.cycle[7] ),
    .B(net131),
    .Y(_1496_));
 sky130_fd_sc_hd__inv_2 _4745_ (.A(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__a221o_1 _4746_ (.A1(net131),
    .A2(_1495_),
    .B1(_1496_),
    .B2(_1492_),
    .C1(net78),
    .X(_1498_));
 sky130_fd_sc_hd__or2_4 _4747_ (.A(net283),
    .B(net341),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_4 _4748_ (.A(net283),
    .B(net341),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_4 _4749_ (.A(_1499_),
    .B(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__nand2_1 _4750_ (.A(_1459_),
    .B(_1462_),
    .Y(_1502_));
 sky130_fd_sc_hd__a31o_1 _4751_ (.A1(_1499_),
    .A2(_1500_),
    .A3(_1502_),
    .B1(_2737_),
    .X(_1503_));
 sky130_fd_sc_hd__a31o_1 _4752_ (.A1(_1459_),
    .A2(_1462_),
    .A3(_1501_),
    .B1(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__nand3_1 _4753_ (.A(net81),
    .B(_1498_),
    .C(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__o21a_2 _4754_ (.A1(_1461_),
    .A2(_1465_),
    .B1(_1459_),
    .X(_1506_));
 sky130_fd_sc_hd__xor2_4 _4755_ (.A(_1501_),
    .B(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(net13),
    .A1(_1507_),
    .S(net327),
    .X(_1508_));
 sky130_fd_sc_hd__o21ai_1 _4757_ (.A1(net148),
    .A2(_1495_),
    .B1(_1401_),
    .Y(_1509_));
 sky130_fd_sc_hd__a22o_1 _4758_ (.A1(net13),
    .A2(_0574_),
    .B1(_1403_),
    .B2(net341),
    .X(_1510_));
 sky130_fd_sc_hd__or2_1 _4759_ (.A(_1509_),
    .B(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__o21a_1 _4760_ (.A1(_2744_),
    .A2(_1508_),
    .B1(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__o2bb2a_1 _4761_ (.A1_N(_2633_),
    .A2_N(_1398_),
    .B1(_1512_),
    .B2(net137),
    .X(_1513_));
 sky130_fd_sc_hd__o221a_1 _4762_ (.A1(\as2650.pc[3] ),
    .A2(_2794_),
    .B1(_1513_),
    .B2(net210),
    .C1(_1505_),
    .X(_1514_));
 sky130_fd_sc_hd__o22a_1 _4763_ (.A1(net283),
    .A2(net52),
    .B1(_1514_),
    .B2(net130),
    .X(_1515_));
 sky130_fd_sc_hd__or2_1 _4764_ (.A(net13),
    .B(net40),
    .X(_1516_));
 sky130_fd_sc_hd__o311a_1 _4765_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1515_),
    .B1(_1516_),
    .C1(net313),
    .X(_0184_));
 sky130_fd_sc_hd__and2_1 _4766_ (.A(net338),
    .B(_0416_),
    .X(_1517_));
 sky130_fd_sc_hd__xnor2_2 _4767_ (.A(_2655_),
    .B(_0416_),
    .Y(_1518_));
 sky130_fd_sc_hd__a31o_2 _4768_ (.A1(_1442_),
    .A2(_1485_),
    .A3(_1488_),
    .B1(_1486_),
    .X(_1519_));
 sky130_fd_sc_hd__xnor2_1 _4769_ (.A(_1518_),
    .B(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_2655_),
    .A1(_1520_),
    .S(net196),
    .X(_1521_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(net339),
    .B(_0413_),
    .Y(_1522_));
 sky130_fd_sc_hd__xnor2_2 _4772_ (.A(net339),
    .B(_0413_),
    .Y(_1523_));
 sky130_fd_sc_hd__a31oi_4 _4773_ (.A1(_1449_),
    .A2(_1477_),
    .A3(_1480_),
    .B1(_1478_),
    .Y(_1524_));
 sky130_fd_sc_hd__xor2_1 _4774_ (.A(_1523_),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _4775_ (.A0(net339),
    .A1(_1525_),
    .S(_2819_),
    .X(_1526_));
 sky130_fd_sc_hd__a2bb2o_2 _4776_ (.A1_N(_2719_),
    .A2_N(_1521_),
    .B1(_1526_),
    .B2(net85),
    .X(_1527_));
 sky130_fd_sc_hd__xnor2_1 _4777_ (.A(net14),
    .B(_1493_),
    .Y(_1528_));
 sky130_fd_sc_hd__o21a_1 _4778_ (.A1(_2715_),
    .A2(_1528_),
    .B1(net81),
    .X(_1529_));
 sky130_fd_sc_hd__nand2_2 _4779_ (.A(net281),
    .B(net338),
    .Y(_1530_));
 sky130_fd_sc_hd__or2_1 _4780_ (.A(net281),
    .B(net338),
    .X(_1531_));
 sky130_fd_sc_hd__nand2_2 _4781_ (.A(_1530_),
    .B(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_2 _4782_ (.A(_1499_),
    .B(_1502_),
    .Y(_1533_));
 sky130_fd_sc_hd__a21oi_4 _4783_ (.A1(_1500_),
    .A2(_1533_),
    .B1(_1532_),
    .Y(_1534_));
 sky130_fd_sc_hd__a31o_1 _4784_ (.A1(_1500_),
    .A2(_1532_),
    .A3(_1533_),
    .B1(_2737_),
    .X(_1535_));
 sky130_fd_sc_hd__o21ai_2 _4785_ (.A1(_1534_),
    .A2(_1535_),
    .B1(_1529_),
    .Y(_1536_));
 sky130_fd_sc_hd__a21o_1 _4786_ (.A1(_2720_),
    .A2(_1527_),
    .B1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__o2bb2a_1 _4787_ (.A1_N(net147),
    .A2_N(_1528_),
    .B1(_0575_),
    .B2(net14),
    .X(_1538_));
 sky130_fd_sc_hd__o211a_1 _4788_ (.A1(net338),
    .A2(_1404_),
    .B1(_1538_),
    .C1(_1401_),
    .X(_1539_));
 sky130_fd_sc_hd__a21o_1 _4789_ (.A1(_2633_),
    .A2(_2654_),
    .B1(_1506_),
    .X(_1540_));
 sky130_fd_sc_hd__a21o_1 _4790_ (.A1(_1500_),
    .A2(_1540_),
    .B1(_1532_),
    .X(_1541_));
 sky130_fd_sc_hd__nand3_1 _4791_ (.A(_1500_),
    .B(_1532_),
    .C(_1540_),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_1541_),
    .B(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(net326),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__or2_1 _4794_ (.A(net14),
    .B(net327),
    .X(_1545_));
 sky130_fd_sc_hd__a31o_1 _4795_ (.A1(_2743_),
    .A2(_1544_),
    .A3(_1545_),
    .B1(_1539_),
    .X(_1546_));
 sky130_fd_sc_hd__a221o_1 _4796_ (.A1(net281),
    .A2(_1398_),
    .B1(_1546_),
    .B2(net132),
    .C1(net210),
    .X(_1547_));
 sky130_fd_sc_hd__o211a_1 _4797_ (.A1(net281),
    .A2(_2794_),
    .B1(_1537_),
    .C1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__o22a_1 _4798_ (.A1(net281),
    .A2(net53),
    .B1(_1548_),
    .B2(net130),
    .X(_1549_));
 sky130_fd_sc_hd__or2_1 _4799_ (.A(net14),
    .B(net40),
    .X(_1550_));
 sky130_fd_sc_hd__o311a_1 _4800_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1549_),
    .B1(_1550_),
    .C1(net316),
    .X(_0185_));
 sky130_fd_sc_hd__a21oi_1 _4801_ (.A1(_1518_),
    .A2(_1519_),
    .B1(_1517_),
    .Y(_1551_));
 sky130_fd_sc_hd__or2_2 _4802_ (.A(net336),
    .B(_0452_),
    .X(_1552_));
 sky130_fd_sc_hd__nand2_1 _4803_ (.A(net336),
    .B(_0452_),
    .Y(_1553_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_1552_),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__xnor2_1 _4805_ (.A(_1551_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(_2657_),
    .A1(_1555_),
    .S(net196),
    .X(_1556_));
 sky130_fd_sc_hd__and2_1 _4807_ (.A(net6),
    .B(_0469_),
    .X(_1557_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(net6),
    .B(_0469_),
    .X(_1558_));
 sky130_fd_sc_hd__and2b_1 _4809_ (.A_N(_1557_),
    .B(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__o21ai_2 _4810_ (.A1(_1523_),
    .A2(_1524_),
    .B1(_1522_),
    .Y(_1560_));
 sky130_fd_sc_hd__xnor2_1 _4811_ (.A(_1559_),
    .B(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(_2657_),
    .A1(_1561_),
    .S(_2819_),
    .X(_1562_));
 sky130_fd_sc_hd__a22o_2 _4813_ (.A1(_2718_),
    .A2(_1556_),
    .B1(_1562_),
    .B2(net86),
    .X(_1563_));
 sky130_fd_sc_hd__and3_1 _4814_ (.A(net15),
    .B(net14),
    .C(_1493_),
    .X(_1564_));
 sky130_fd_sc_hd__a21oi_1 _4815_ (.A1(net14),
    .A2(_1493_),
    .B1(net15),
    .Y(_1565_));
 sky130_fd_sc_hd__or2_1 _4816_ (.A(_1564_),
    .B(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__a221o_1 _4817_ (.A1(_1496_),
    .A2(_1563_),
    .B1(_1566_),
    .B2(net131),
    .C1(net78),
    .X(_1567_));
 sky130_fd_sc_hd__nand2_2 _4818_ (.A(net279),
    .B(net337),
    .Y(_1568_));
 sky130_fd_sc_hd__or2_4 _4819_ (.A(net279),
    .B(net337),
    .X(_1569_));
 sky130_fd_sc_hd__nand2_4 _4820_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__a21o_1 _4821_ (.A1(net281),
    .A2(net338),
    .B1(_1534_),
    .X(_1571_));
 sky130_fd_sc_hd__xor2_2 _4822_ (.A(_1570_),
    .B(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__o211a_1 _4823_ (.A1(_2737_),
    .A2(_1572_),
    .B1(_1567_),
    .C1(net81),
    .X(_1573_));
 sky130_fd_sc_hd__nor2_1 _4824_ (.A(net153),
    .B(_1566_),
    .Y(_1574_));
 sky130_fd_sc_hd__a221o_1 _4825_ (.A1(net15),
    .A2(_0574_),
    .B1(_1403_),
    .B2(net337),
    .C1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__nand2_4 _4826_ (.A(net141),
    .B(_0579_),
    .Y(_1576_));
 sky130_fd_sc_hd__o22a_1 _4827_ (.A1(net279),
    .A2(_1399_),
    .B1(_1575_),
    .B2(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_2 _4828_ (.A(_1530_),
    .B(_1541_),
    .Y(_1578_));
 sky130_fd_sc_hd__xnor2_2 _4829_ (.A(_1570_),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__and2_1 _4830_ (.A(net15),
    .B(net311),
    .X(_1580_));
 sky130_fd_sc_hd__a2111o_1 _4831_ (.A1(net326),
    .A2(_1579_),
    .B1(_1580_),
    .C1(_2744_),
    .D1(_1394_),
    .X(_1581_));
 sky130_fd_sc_hd__a21oi_1 _4832_ (.A1(_1577_),
    .A2(_1581_),
    .B1(net65),
    .Y(_1582_));
 sky130_fd_sc_hd__a2bb2o_1 _4833_ (.A1_N(net279),
    .A2_N(net52),
    .B1(_1573_),
    .B2(net129),
    .X(_1583_));
 sky130_fd_sc_hd__o21ai_1 _4834_ (.A1(_1582_),
    .A2(_1583_),
    .B1(net39),
    .Y(_1584_));
 sky130_fd_sc_hd__o211a_1 _4835_ (.A1(net15),
    .A2(net38),
    .B1(_1584_),
    .C1(net314),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _4836_ (.A(net334),
    .B(_0518_),
    .X(_1585_));
 sky130_fd_sc_hd__or2_2 _4837_ (.A(net334),
    .B(_0518_),
    .X(_1586_));
 sky130_fd_sc_hd__nand2b_2 _4838_ (.A_N(_1585_),
    .B(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__a221o_2 _4839_ (.A1(net336),
    .A2(_0452_),
    .B1(_1518_),
    .B2(_1519_),
    .C1(_1517_),
    .X(_1588_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(_1552_),
    .B(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__xor2_2 _4841_ (.A(_1587_),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__nand2_1 _4842_ (.A(_2658_),
    .B(_2784_),
    .Y(_1591_));
 sky130_fd_sc_hd__o211a_1 _4843_ (.A1(_2784_),
    .A2(_1590_),
    .B1(_1591_),
    .C1(_2718_),
    .X(_1592_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(net335),
    .B(_0515_),
    .Y(_1593_));
 sky130_fd_sc_hd__inv_2 _4845_ (.A(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__or2_2 _4846_ (.A(net335),
    .B(_0515_),
    .X(_1595_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_1593_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__a21o_2 _4848_ (.A1(_1558_),
    .A2(_1560_),
    .B1(_1557_),
    .X(_1597_));
 sky130_fd_sc_hd__xnor2_1 _4849_ (.A(_1596_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_2658_),
    .B(_2820_),
    .Y(_1599_));
 sky130_fd_sc_hd__o211a_1 _4851_ (.A1(_2820_),
    .A2(_1598_),
    .B1(_1599_),
    .C1(net86),
    .X(_1600_));
 sky130_fd_sc_hd__o21a_2 _4852_ (.A1(_1592_),
    .A2(_1600_),
    .B1(_2720_),
    .X(_1601_));
 sky130_fd_sc_hd__and2_2 _4853_ (.A(net16),
    .B(_1564_),
    .X(_1602_));
 sky130_fd_sc_hd__nor2_1 _4854_ (.A(net16),
    .B(_1564_),
    .Y(_1603_));
 sky130_fd_sc_hd__or2_1 _4855_ (.A(_1602_),
    .B(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__o21ai_1 _4856_ (.A1(_2715_),
    .A2(_1604_),
    .B1(net81),
    .Y(_1605_));
 sky130_fd_sc_hd__and2_4 _4857_ (.A(net278),
    .B(net332),
    .X(_1606_));
 sky130_fd_sc_hd__nor2_4 _4858_ (.A(net278),
    .B(net332),
    .Y(_1607_));
 sky130_fd_sc_hd__nor2_8 _4859_ (.A(_1606_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_1530_),
    .B(_1568_),
    .Y(_1609_));
 sky130_fd_sc_hd__o21a_2 _4861_ (.A1(_1534_),
    .A2(_1609_),
    .B1(_1569_),
    .X(_1610_));
 sky130_fd_sc_hd__xor2_2 _4862_ (.A(_1608_),
    .B(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__a211o_1 _4863_ (.A1(net78),
    .A2(_1611_),
    .B1(_1605_),
    .C1(_1601_),
    .X(_1612_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(net149),
    .B(_1604_),
    .Y(_1613_));
 sky130_fd_sc_hd__o221a_1 _4865_ (.A1(net16),
    .A2(_0575_),
    .B1(_1404_),
    .B2(net333),
    .C1(_1401_),
    .X(_1614_));
 sky130_fd_sc_hd__a21bo_4 _4866_ (.A1(_1569_),
    .A2(_1578_),
    .B1_N(_1568_),
    .X(_1615_));
 sky130_fd_sc_hd__xor2_2 _4867_ (.A(_1608_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(net16),
    .A1(_1616_),
    .S(net326),
    .X(_1617_));
 sky130_fd_sc_hd__a22o_1 _4869_ (.A1(_1613_),
    .A2(_1614_),
    .B1(_1617_),
    .B2(_2743_),
    .X(_1618_));
 sky130_fd_sc_hd__a221o_1 _4870_ (.A1(net278),
    .A2(_1400_),
    .B1(_1618_),
    .B2(net64),
    .C1(net212),
    .X(_1619_));
 sky130_fd_sc_hd__a21oi_1 _4871_ (.A1(_1612_),
    .A2(_1619_),
    .B1(net130),
    .Y(_1620_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(net278),
    .B(net52),
    .Y(_1621_));
 sky130_fd_sc_hd__o21ai_1 _4873_ (.A1(_1620_),
    .A2(_1621_),
    .B1(net38),
    .Y(_1622_));
 sky130_fd_sc_hd__o211a_1 _4874_ (.A1(net16),
    .A2(net38),
    .B1(_1622_),
    .C1(net314),
    .X(_0187_));
 sky130_fd_sc_hd__a31o_1 _4875_ (.A1(_1552_),
    .A2(_1586_),
    .A3(_1588_),
    .B1(_1585_),
    .X(_1623_));
 sky130_fd_sc_hd__and2_1 _4876_ (.A(net329),
    .B(_0552_),
    .X(_1624_));
 sky130_fd_sc_hd__or2_2 _4877_ (.A(net329),
    .B(_0552_),
    .X(_1625_));
 sky130_fd_sc_hd__and2b_1 _4878_ (.A_N(_1624_),
    .B(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_1623_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__o21a_1 _4880_ (.A1(_1623_),
    .A2(_1626_),
    .B1(net196),
    .X(_1628_));
 sky130_fd_sc_hd__o2bb2a_1 _4881_ (.A1_N(_1627_),
    .A2_N(_1628_),
    .B1(_2650_),
    .B2(net196),
    .X(_1629_));
 sky130_fd_sc_hd__a21oi_1 _4882_ (.A1(_1595_),
    .A2(_1597_),
    .B1(_1594_),
    .Y(_1630_));
 sky130_fd_sc_hd__xnor2_1 _4883_ (.A(net329),
    .B(_0550_),
    .Y(_1631_));
 sky130_fd_sc_hd__a21oi_1 _4884_ (.A1(_1630_),
    .A2(_1631_),
    .B1(_2820_),
    .Y(_1632_));
 sky130_fd_sc_hd__o21ai_1 _4885_ (.A1(_1630_),
    .A2(_1631_),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_1 _4886_ (.A(net329),
    .B(_2820_),
    .Y(_1634_));
 sky130_fd_sc_hd__a32o_2 _4887_ (.A1(net86),
    .A2(_1633_),
    .A3(_1634_),
    .B1(_2718_),
    .B2(_1629_),
    .X(_1635_));
 sky130_fd_sc_hd__xnor2_1 _4888_ (.A(net17),
    .B(_1602_),
    .Y(_1636_));
 sky130_fd_sc_hd__a221o_1 _4889_ (.A1(_1496_),
    .A2(_1635_),
    .B1(_1636_),
    .B2(_2714_),
    .C1(net79),
    .X(_1637_));
 sky130_fd_sc_hd__and2_2 _4890_ (.A(net275),
    .B(net332),
    .X(_1638_));
 sky130_fd_sc_hd__nor2_2 _4891_ (.A(net275),
    .B(net332),
    .Y(_1639_));
 sky130_fd_sc_hd__nor2_8 _4892_ (.A(_1638_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__a21o_2 _4893_ (.A1(_1608_),
    .A2(_1610_),
    .B1(_1606_),
    .X(_1641_));
 sky130_fd_sc_hd__xnor2_4 _4894_ (.A(_1640_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__o211ai_1 _4895_ (.A1(_2737_),
    .A2(_1642_),
    .B1(_1637_),
    .C1(net81),
    .Y(_1643_));
 sky130_fd_sc_hd__nor2_1 _4896_ (.A(net153),
    .B(_1636_),
    .Y(_1644_));
 sky130_fd_sc_hd__a221o_1 _4897_ (.A1(net17),
    .A2(_0574_),
    .B1(_1403_),
    .B2(net328),
    .C1(_1576_),
    .X(_1645_));
 sky130_fd_sc_hd__o22a_1 _4898_ (.A1(net276),
    .A2(_1399_),
    .B1(_1644_),
    .B2(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__a21oi_4 _4899_ (.A1(_1608_),
    .A2(_1615_),
    .B1(_1606_),
    .Y(_1647_));
 sky130_fd_sc_hd__xnor2_4 _4900_ (.A(_1640_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__a211o_1 _4901_ (.A1(net327),
    .A2(_1648_),
    .B1(_2744_),
    .C1(net137),
    .X(_1649_));
 sky130_fd_sc_hd__a211o_1 _4902_ (.A1(net17),
    .A2(net312),
    .B1(net210),
    .C1(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__o211a_1 _4903_ (.A1(net212),
    .A2(_1646_),
    .B1(_1650_),
    .C1(_1643_),
    .X(_1651_));
 sky130_fd_sc_hd__o22a_1 _4904_ (.A1(net276),
    .A2(net53),
    .B1(_1651_),
    .B2(net130),
    .X(_1652_));
 sky130_fd_sc_hd__or2_1 _4905_ (.A(net17),
    .B(net40),
    .X(_1653_));
 sky130_fd_sc_hd__o311a_1 _4906_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1652_),
    .B1(_1653_),
    .C1(net316),
    .X(_0188_));
 sky130_fd_sc_hd__a221oi_4 _4907_ (.A1(net329),
    .A2(_0550_),
    .B1(_1595_),
    .B2(_1597_),
    .C1(_1594_),
    .Y(_1654_));
 sky130_fd_sc_hd__o21ai_4 _4908_ (.A1(net329),
    .A2(_0550_),
    .B1(_2819_),
    .Y(_1655_));
 sky130_fd_sc_hd__or2_1 _4909_ (.A(_1654_),
    .B(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__xnor2_1 _4910_ (.A(net310),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__a311o_4 _4911_ (.A1(_1552_),
    .A2(_1586_),
    .A3(_1588_),
    .B1(_1624_),
    .C1(_1585_),
    .X(_1658_));
 sky130_fd_sc_hd__and2_1 _4912_ (.A(net197),
    .B(_1625_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_1 _4913_ (.A(_1658_),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__xnor2_1 _4914_ (.A(net310),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__o22a_1 _4915_ (.A1(net84),
    .A2(_1657_),
    .B1(_1661_),
    .B2(_2719_),
    .X(_1662_));
 sky130_fd_sc_hd__and3_1 _4916_ (.A(net18),
    .B(net17),
    .C(_1602_),
    .X(_1663_));
 sky130_fd_sc_hd__a21oi_1 _4917_ (.A1(net17),
    .A2(_1602_),
    .B1(net18),
    .Y(_1664_));
 sky130_fd_sc_hd__nor2_1 _4918_ (.A(_1663_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__o221a_1 _4919_ (.A1(_1497_),
    .A2(_1662_),
    .B1(_1665_),
    .B2(_2715_),
    .C1(_2737_),
    .X(_1666_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(net274),
    .B(net332),
    .Y(_1667_));
 sky130_fd_sc_hd__or2_1 _4921_ (.A(net274),
    .B(net332),
    .X(_1668_));
 sky130_fd_sc_hd__and2_2 _4922_ (.A(_1667_),
    .B(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__a41o_1 _4923_ (.A1(_1569_),
    .A2(_1608_),
    .A3(_1609_),
    .A4(_1640_),
    .B1(_1606_),
    .X(_1670_));
 sky130_fd_sc_hd__or2_1 _4924_ (.A(_1638_),
    .B(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__or4b_2 _4925_ (.A(_1570_),
    .B(_1606_),
    .C(_1607_),
    .D_N(_1640_),
    .X(_1672_));
 sky130_fd_sc_hd__inv_2 _4926_ (.A(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__a21o_1 _4927_ (.A1(_1534_),
    .A2(_1673_),
    .B1(_1671_),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_1669_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__or2_1 _4929_ (.A(_1669_),
    .B(_1674_),
    .X(_1676_));
 sky130_fd_sc_hd__and3_1 _4930_ (.A(net78),
    .B(_1675_),
    .C(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__or4_1 _4931_ (.A(net80),
    .B(net130),
    .C(_1666_),
    .D(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__o21ba_1 _4932_ (.A1(_1541_),
    .A2(_1672_),
    .B1_N(_1671_),
    .X(_1679_));
 sky130_fd_sc_hd__nand2b_1 _4933_ (.A_N(_1679_),
    .B(_1669_),
    .Y(_1680_));
 sky130_fd_sc_hd__xor2_2 _4934_ (.A(_1669_),
    .B(_1679_),
    .X(_1681_));
 sky130_fd_sc_hd__o21ai_1 _4935_ (.A1(net18),
    .A2(net326),
    .B1(_1395_),
    .Y(_1682_));
 sky130_fd_sc_hd__a21o_1 _4936_ (.A1(net326),
    .A2(_1681_),
    .B1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__o22a_1 _4937_ (.A1(net18),
    .A2(_0575_),
    .B1(_1404_),
    .B2(net310),
    .X(_1684_));
 sky130_fd_sc_hd__o21ai_1 _4938_ (.A1(net148),
    .A2(_1665_),
    .B1(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__o221a_1 _4939_ (.A1(_2631_),
    .A2(_1399_),
    .B1(_1576_),
    .B2(_1685_),
    .C1(net69),
    .X(_1686_));
 sky130_fd_sc_hd__o2bb2a_1 _4940_ (.A1_N(_1683_),
    .A2_N(_1686_),
    .B1(net274),
    .B2(net52),
    .X(_1687_));
 sky130_fd_sc_hd__a21bo_1 _4941_ (.A1(_1678_),
    .A2(_1687_),
    .B1_N(net38),
    .X(_1688_));
 sky130_fd_sc_hd__o211a_1 _4942_ (.A1(net18),
    .A2(net38),
    .B1(_1688_),
    .C1(net314),
    .X(_0189_));
 sky130_fd_sc_hd__nor2_1 _4943_ (.A(_2660_),
    .B(_2661_),
    .Y(_1689_));
 sky130_fd_sc_hd__o31a_2 _4944_ (.A1(_2660_),
    .A2(_2661_),
    .A3(_1660_),
    .B1(_2718_),
    .X(_1690_));
 sky130_fd_sc_hd__or3b_4 _4945_ (.A(_1654_),
    .B(_1655_),
    .C_N(_1689_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(net85),
    .B(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__a21oi_2 _4947_ (.A1(net85),
    .A2(_1691_),
    .B1(_1690_),
    .Y(_1693_));
 sky130_fd_sc_hd__a31o_1 _4948_ (.A1(net310),
    .A2(_1658_),
    .A3(_1659_),
    .B1(\as2650.addr_buff[1] ),
    .X(_1694_));
 sky130_fd_sc_hd__o21a_1 _4949_ (.A1(_2660_),
    .A2(_1656_),
    .B1(_2661_),
    .X(_1695_));
 sky130_fd_sc_hd__a2bb2o_1 _4950_ (.A1_N(_1695_),
    .A2_N(_1692_),
    .B1(_1690_),
    .B2(_1694_),
    .X(_1696_));
 sky130_fd_sc_hd__and2_2 _4951_ (.A(net19),
    .B(_1663_),
    .X(_1697_));
 sky130_fd_sc_hd__nor2_1 _4952_ (.A(net19),
    .B(_1663_),
    .Y(_1698_));
 sky130_fd_sc_hd__or2_1 _4953_ (.A(_1697_),
    .B(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__a2bb2o_1 _4954_ (.A1_N(_2715_),
    .A2_N(_1699_),
    .B1(_1696_),
    .B2(_1496_),
    .X(_1700_));
 sky130_fd_sc_hd__xnor2_4 _4955_ (.A(net273),
    .B(net332),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _4956_ (.A(_1667_),
    .B(_1675_),
    .Y(_1702_));
 sky130_fd_sc_hd__xnor2_2 _4957_ (.A(_1701_),
    .B(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__mux2_1 _4958_ (.A0(_1700_),
    .A1(_1703_),
    .S(net79),
    .X(_1704_));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(net153),
    .B(_1699_),
    .Y(_1705_));
 sky130_fd_sc_hd__a221o_1 _4960_ (.A1(net19),
    .A2(_0574_),
    .B1(_1403_),
    .B2(\as2650.addr_buff[1] ),
    .C1(_1576_),
    .X(_1706_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(\as2650.addr_buff[1] ),
    .B(net155),
    .Y(_1707_));
 sky130_fd_sc_hd__o22a_1 _4962_ (.A1(net273),
    .A2(_1399_),
    .B1(_1705_),
    .B2(_1706_),
    .X(_1708_));
 sky130_fd_sc_hd__or2_1 _4963_ (.A(net212),
    .B(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _4964_ (.A(_1667_),
    .B(_1680_),
    .Y(_1710_));
 sky130_fd_sc_hd__xnor2_1 _4965_ (.A(_1701_),
    .B(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__a211o_1 _4966_ (.A1(net326),
    .A2(_1711_),
    .B1(_2744_),
    .C1(net137),
    .X(_1712_));
 sky130_fd_sc_hd__a211o_1 _4967_ (.A1(net19),
    .A2(net312),
    .B1(net210),
    .C1(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__o211a_1 _4968_ (.A1(net80),
    .A2(_1704_),
    .B1(_1709_),
    .C1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o22a_1 _4969_ (.A1(net273),
    .A2(net53),
    .B1(_1714_),
    .B2(net130),
    .X(_1715_));
 sky130_fd_sc_hd__or2_1 _4970_ (.A(net19),
    .B(net40),
    .X(_1716_));
 sky130_fd_sc_hd__o311a_1 _4971_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1715_),
    .B1(_1716_),
    .C1(net316),
    .X(_0190_));
 sky130_fd_sc_hd__nand3_2 _4972_ (.A(_2718_),
    .B(_1658_),
    .C(_1659_),
    .Y(_1717_));
 sky130_fd_sc_hd__o31ai_4 _4973_ (.A1(net84),
    .A2(_1654_),
    .A3(_1655_),
    .B1(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__and3_2 _4974_ (.A(net310),
    .B(\as2650.addr_buff[1] ),
    .C(\as2650.addr_buff[2] ),
    .X(_1719_));
 sky130_fd_sc_hd__a2bb2o_1 _4975_ (.A1_N(\as2650.addr_buff[2] ),
    .A2_N(_1693_),
    .B1(_1718_),
    .B2(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__xnor2_1 _4976_ (.A(net20),
    .B(_1697_),
    .Y(_1721_));
 sky130_fd_sc_hd__a221o_1 _4977_ (.A1(_1496_),
    .A2(_1720_),
    .B1(_1721_),
    .B2(net131),
    .C1(net78),
    .X(_1722_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(net271),
    .B(net332),
    .Y(_1723_));
 sky130_fd_sc_hd__or2_1 _4979_ (.A(net271),
    .B(net332),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_2 _4980_ (.A(_1723_),
    .B(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__inv_2 _4981_ (.A(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__o21ai_2 _4982_ (.A1(net273),
    .A2(net274),
    .B1(net332),
    .Y(_1727_));
 sky130_fd_sc_hd__or2_2 _4983_ (.A(_1675_),
    .B(_1701_),
    .X(_1728_));
 sky130_fd_sc_hd__a21oi_1 _4984_ (.A1(_1727_),
    .A2(_1728_),
    .B1(_1725_),
    .Y(_1729_));
 sky130_fd_sc_hd__a31o_1 _4985_ (.A1(_1725_),
    .A2(_1727_),
    .A3(_1728_),
    .B1(_2737_),
    .X(_1730_));
 sky130_fd_sc_hd__o2111a_1 _4986_ (.A1(_1729_),
    .A2(_1730_),
    .B1(net81),
    .C1(net129),
    .D1(_1722_),
    .X(_1731_));
 sky130_fd_sc_hd__or2_1 _4987_ (.A(_1680_),
    .B(_1701_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_1727_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__xnor2_1 _4989_ (.A(_1726_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(net326),
    .B(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__o211a_1 _4991_ (.A1(net20),
    .A2(net326),
    .B1(_1395_),
    .C1(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__nand2_1 _4992_ (.A(net149),
    .B(_1721_),
    .Y(_1737_));
 sky130_fd_sc_hd__o221a_1 _4993_ (.A1(net20),
    .A2(_0575_),
    .B1(_1404_),
    .B2(\as2650.addr_buff[2] ),
    .C1(net141),
    .X(_1738_));
 sky130_fd_sc_hd__a22o_1 _4994_ (.A1(net271),
    .A2(_1396_),
    .B1(_1737_),
    .B2(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__a221o_1 _4995_ (.A1(net271),
    .A2(_1394_),
    .B1(_1739_),
    .B2(_0579_),
    .C1(net65),
    .X(_1740_));
 sky130_fd_sc_hd__o22ai_1 _4996_ (.A1(net271),
    .A2(net52),
    .B1(_1736_),
    .B2(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__o21ai_1 _4997_ (.A1(_1731_),
    .A2(_1741_),
    .B1(net39),
    .Y(_1742_));
 sky130_fd_sc_hd__o211a_1 _4998_ (.A1(net20),
    .A2(net38),
    .B1(_1742_),
    .C1(net314),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _4999_ (.A(\as2650.addr_buff[2] ),
    .B(_2716_),
    .Y(_1743_));
 sky130_fd_sc_hd__a2111o_1 _5000_ (.A1(net85),
    .A2(_1691_),
    .B1(_1743_),
    .C1(_1690_),
    .D1(\as2650.addr_buff[3] ),
    .X(_1744_));
 sky130_fd_sc_hd__a21bo_1 _5001_ (.A1(_1718_),
    .A2(_1719_),
    .B1_N(\as2650.addr_buff[3] ),
    .X(_1745_));
 sky130_fd_sc_hd__and3_1 _5002_ (.A(net21),
    .B(net20),
    .C(_1697_),
    .X(_1746_));
 sky130_fd_sc_hd__a21oi_1 _5003_ (.A1(net20),
    .A2(_1697_),
    .B1(net21),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _5004_ (.A(_1746_),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a32o_1 _5005_ (.A1(_1496_),
    .A2(_1744_),
    .A3(_1745_),
    .B1(_1748_),
    .B2(net131),
    .X(_1749_));
 sky130_fd_sc_hd__xor2_1 _5006_ (.A(net270),
    .B(net333),
    .X(_1750_));
 sky130_fd_sc_hd__clkinv_2 _5007_ (.A(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__a21oi_1 _5008_ (.A1(net271),
    .A2(net333),
    .B1(_1729_),
    .Y(_1752_));
 sky130_fd_sc_hd__xnor2_1 _5009_ (.A(_1751_),
    .B(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__mux2_1 _5010_ (.A0(_1749_),
    .A1(_1753_),
    .S(net78),
    .X(_1754_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(net153),
    .B(_1748_),
    .Y(_1755_));
 sky130_fd_sc_hd__a221o_1 _5012_ (.A1(net21),
    .A2(_0574_),
    .B1(_1403_),
    .B2(\as2650.addr_buff[3] ),
    .C1(net143),
    .X(_1756_));
 sky130_fd_sc_hd__o22a_1 _5013_ (.A1(net270),
    .A2(net63),
    .B1(_1755_),
    .B2(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__a21bo_1 _5014_ (.A1(_1726_),
    .A2(_1733_),
    .B1_N(_1723_),
    .X(_1758_));
 sky130_fd_sc_hd__xnor2_1 _5015_ (.A(_1751_),
    .B(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__mux2_1 _5016_ (.A0(net21),
    .A1(_1759_),
    .S(net327),
    .X(_1760_));
 sky130_fd_sc_hd__o32a_1 _5017_ (.A1(net137),
    .A2(_2744_),
    .A3(_1760_),
    .B1(_1757_),
    .B2(net146),
    .X(_1761_));
 sky130_fd_sc_hd__o22a_1 _5018_ (.A1(net270),
    .A2(net64),
    .B1(_1761_),
    .B2(net215),
    .X(_1762_));
 sky130_fd_sc_hd__a2bb2o_1 _5019_ (.A1_N(net212),
    .A2_N(_1762_),
    .B1(_1754_),
    .B2(net81),
    .X(_1763_));
 sky130_fd_sc_hd__a2bb2o_1 _5020_ (.A1_N(net270),
    .A2_N(net52),
    .B1(_1763_),
    .B2(net129),
    .X(_1764_));
 sky130_fd_sc_hd__nand2_1 _5021_ (.A(net38),
    .B(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__o211a_1 _5022_ (.A1(net21),
    .A2(net38),
    .B1(_1765_),
    .C1(net314),
    .X(_0192_));
 sky130_fd_sc_hd__a31o_1 _5023_ (.A1(\as2650.addr_buff[3] ),
    .A2(_1718_),
    .A3(_1719_),
    .B1(_2662_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(\as2650.addr_buff[2] ),
    .B(\as2650.addr_buff[3] ),
    .Y(_1767_));
 sky130_fd_sc_hd__inv_2 _5025_ (.A(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__o211ai_2 _5026_ (.A1(_2716_),
    .A2(_1768_),
    .B1(_1693_),
    .C1(_2662_),
    .Y(_1769_));
 sky130_fd_sc_hd__xnor2_1 _5027_ (.A(net23),
    .B(_1746_),
    .Y(_1770_));
 sky130_fd_sc_hd__a32o_1 _5028_ (.A1(_1496_),
    .A2(_1766_),
    .A3(_1769_),
    .B1(_1770_),
    .B2(net131),
    .X(_1771_));
 sky130_fd_sc_hd__xor2_4 _5029_ (.A(net269),
    .B(net333),
    .X(_1772_));
 sky130_fd_sc_hd__o41a_1 _5030_ (.A1(net270),
    .A2(net271),
    .A3(net273),
    .A4(net274),
    .B1(net333),
    .X(_1773_));
 sky130_fd_sc_hd__inv_2 _5031_ (.A(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__o31a_1 _5032_ (.A1(_1725_),
    .A2(_1728_),
    .A3(_1751_),
    .B1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__xnor2_1 _5033_ (.A(_1772_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(net78),
    .B(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__o21ai_1 _5035_ (.A1(net78),
    .A2(_1771_),
    .B1(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nor2_1 _5036_ (.A(net153),
    .B(_1770_),
    .Y(_1779_));
 sky130_fd_sc_hd__a221o_1 _5037_ (.A1(net23),
    .A2(_0574_),
    .B1(_1403_),
    .B2(\as2650.addr_buff[4] ),
    .C1(net143),
    .X(_1780_));
 sky130_fd_sc_hd__o22a_1 _5038_ (.A1(net269),
    .A2(net63),
    .B1(_1779_),
    .B2(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__o31a_1 _5039_ (.A1(_1725_),
    .A2(_1732_),
    .A3(_1751_),
    .B1(_1774_),
    .X(_1782_));
 sky130_fd_sc_hd__xnor2_2 _5040_ (.A(_1772_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(net23),
    .A1(_1783_),
    .S(net327),
    .X(_1784_));
 sky130_fd_sc_hd__o32a_1 _5042_ (.A1(net92),
    .A2(_2744_),
    .A3(_1784_),
    .B1(_1781_),
    .B2(net146),
    .X(_1785_));
 sky130_fd_sc_hd__o22a_1 _5043_ (.A1(net269),
    .A2(net64),
    .B1(_1785_),
    .B2(net215),
    .X(_1786_));
 sky130_fd_sc_hd__o22a_1 _5044_ (.A1(net80),
    .A2(_1778_),
    .B1(_1786_),
    .B2(net212),
    .X(_1787_));
 sky130_fd_sc_hd__o22a_1 _5045_ (.A1(net269),
    .A2(net52),
    .B1(_1787_),
    .B2(net130),
    .X(_1788_));
 sky130_fd_sc_hd__or2_1 _5046_ (.A(net23),
    .B(net38),
    .X(_1789_));
 sky130_fd_sc_hd__o311a_1 _5047_ (.A1(_1373_),
    .A2(_1379_),
    .A3(_1788_),
    .B1(_1789_),
    .C1(net314),
    .X(_0193_));
 sky130_fd_sc_hd__and3b_1 _5048_ (.A_N(_1346_),
    .B(_1365_),
    .C(_0587_),
    .X(_1790_));
 sky130_fd_sc_hd__nor2_1 _5049_ (.A(_2717_),
    .B(net80),
    .Y(_1791_));
 sky130_fd_sc_hd__and3_1 _5050_ (.A(net328),
    .B(net79),
    .C(_2738_),
    .X(_1792_));
 sky130_fd_sc_hd__or4_1 _5051_ (.A(\as2650.cycle[7] ),
    .B(_2708_),
    .C(_2713_),
    .D(net80),
    .X(_1793_));
 sky130_fd_sc_hd__or2_1 _5052_ (.A(_1791_),
    .B(_1792_),
    .X(_1794_));
 sky130_fd_sc_hd__nor2_1 _5053_ (.A(net229),
    .B(net84),
    .Y(_1795_));
 sky130_fd_sc_hd__nand2_2 _5054_ (.A(net309),
    .B(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__o31a_1 _5055_ (.A1(net328),
    .A2(net158),
    .A3(net145),
    .B1(_2728_),
    .X(_1797_));
 sky130_fd_sc_hd__o2111a_1 _5056_ (.A1(net229),
    .A2(_1496_),
    .B1(_1796_),
    .C1(_1797_),
    .D1(_1337_),
    .X(_1798_));
 sky130_fd_sc_hd__nand2_2 _5057_ (.A(net235),
    .B(_2677_),
    .Y(_1799_));
 sky130_fd_sc_hd__or4_1 _5058_ (.A(net94),
    .B(_2727_),
    .C(net65),
    .D(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__and4b_1 _5059_ (.A_N(_1794_),
    .B(_1798_),
    .C(_1800_),
    .D(_1369_),
    .X(_1801_));
 sky130_fd_sc_hd__o2bb2a_1 _5060_ (.A1_N(net213),
    .A2_N(_2688_),
    .B1(net128),
    .B2(_0760_),
    .X(_1802_));
 sky130_fd_sc_hd__o211a_1 _5061_ (.A1(net87),
    .A2(_1370_),
    .B1(_1802_),
    .C1(_0829_),
    .X(_1803_));
 sky130_fd_sc_hd__and4_1 _5062_ (.A(_1353_),
    .B(_1360_),
    .C(_1801_),
    .D(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__and3_2 _5063_ (.A(_1378_),
    .B(_1790_),
    .C(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__a211o_1 _5064_ (.A1(net10),
    .A2(_2764_),
    .B1(_0573_),
    .C1(net96),
    .X(_1806_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(net213),
    .B(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__o21ai_1 _5066_ (.A1(net87),
    .A2(_0836_),
    .B1(net171),
    .Y(_1808_));
 sky130_fd_sc_hd__a31o_1 _5067_ (.A1(net24),
    .A2(net87),
    .A3(net126),
    .B1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__a31o_1 _5068_ (.A1(net24),
    .A2(net101),
    .A3(net133),
    .B1(net210),
    .X(_1810_));
 sky130_fd_sc_hd__and4_1 _5069_ (.A(net129),
    .B(_1807_),
    .C(_1809_),
    .D(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(net24),
    .A1(_1811_),
    .S(_1805_),
    .X(_1812_));
 sky130_fd_sc_hd__and2_1 _5071_ (.A(net316),
    .B(_1812_),
    .X(_0194_));
 sky130_fd_sc_hd__and3_1 _5072_ (.A(net328),
    .B(_2741_),
    .C(_0579_),
    .X(_1813_));
 sky130_fd_sc_hd__a31o_1 _5073_ (.A1(net172),
    .A2(_1393_),
    .A3(_1396_),
    .B1(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__inv_2 _5074_ (.A(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__and3_1 _5075_ (.A(net173),
    .B(_2669_),
    .C(net145),
    .X(_1816_));
 sky130_fd_sc_hd__o21a_1 _5076_ (.A1(_2682_),
    .A2(_2703_),
    .B1(net101),
    .X(_1817_));
 sky130_fd_sc_hd__and3b_1 _5077_ (.A_N(_2683_),
    .B(_1816_),
    .C(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__a311o_1 _5078_ (.A1(net293),
    .A2(_2680_),
    .A3(_2683_),
    .B1(_2845_),
    .C1(_1358_),
    .X(_1819_));
 sky130_fd_sc_hd__or3b_2 _5079_ (.A(_1819_),
    .B(_1818_),
    .C_N(_1369_),
    .X(_1820_));
 sky130_fd_sc_hd__or3b_1 _5080_ (.A(_1362_),
    .B(_1820_),
    .C_N(_1361_),
    .X(_1821_));
 sky130_fd_sc_hd__o221a_1 _5081_ (.A1(net89),
    .A2(net125),
    .B1(_1397_),
    .B2(net172),
    .C1(_1337_),
    .X(_1822_));
 sky130_fd_sc_hd__o211a_1 _5082_ (.A1(_1343_),
    .A2(_1345_),
    .B1(_1352_),
    .C1(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_1366_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__a211o_2 _5084_ (.A1(net229),
    .A2(_1814_),
    .B1(_1821_),
    .C1(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__nor2_1 _5085_ (.A(_1379_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__a311o_1 _5086_ (.A1(net25),
    .A2(net158),
    .A3(_0836_),
    .B1(net136),
    .C1(net235),
    .X(_1827_));
 sky130_fd_sc_hd__a21o_1 _5087_ (.A1(net97),
    .A2(_0576_),
    .B1(_1403_),
    .X(_1828_));
 sky130_fd_sc_hd__a32o_1 _5088_ (.A1(net25),
    .A2(_1401_),
    .A3(_1828_),
    .B1(net328),
    .B2(net146),
    .X(_1829_));
 sky130_fd_sc_hd__o21ai_1 _5089_ (.A1(_1394_),
    .A2(_1829_),
    .B1(_1827_),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _5090_ (.A(net229),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__a31o_1 _5091_ (.A1(net25),
    .A2(net158),
    .A3(_0576_),
    .B1(net80),
    .X(_1832_));
 sky130_fd_sc_hd__a31o_1 _5092_ (.A1(_2728_),
    .A2(_1831_),
    .A3(_1832_),
    .B1(net130),
    .X(_1833_));
 sky130_fd_sc_hd__or3_1 _5093_ (.A(_1379_),
    .B(_1825_),
    .C(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__o211a_1 _5094_ (.A1(net25),
    .A2(_1826_),
    .B1(_1834_),
    .C1(net316),
    .X(_0195_));
 sky130_fd_sc_hd__or3_1 _5095_ (.A(_2726_),
    .B(net59),
    .C(_1795_),
    .X(_1835_));
 sky130_fd_sc_hd__or3_1 _5096_ (.A(net96),
    .B(_2721_),
    .C(_2727_),
    .X(_1836_));
 sky130_fd_sc_hd__or3b_4 _5097_ (.A(net294),
    .B(_1836_),
    .C_N(_1835_),
    .X(_1837_));
 sky130_fd_sc_hd__a21oi_1 _5098_ (.A1(\as2650.addr_buff[5] ),
    .A2(_2732_),
    .B1(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__a211oi_1 _5099_ (.A1(_2640_),
    .A2(_1837_),
    .B1(_1838_),
    .C1(net322),
    .Y(_0196_));
 sky130_fd_sc_hd__a21oi_1 _5100_ (.A1(\as2650.addr_buff[6] ),
    .A2(_2732_),
    .B1(_1837_),
    .Y(_1839_));
 sky130_fd_sc_hd__a211oi_1 _5101_ (.A1(_2639_),
    .A2(_1837_),
    .B1(_1839_),
    .C1(net322),
    .Y(_0197_));
 sky130_fd_sc_hd__a31o_1 _5102_ (.A1(net140),
    .A2(net202),
    .A3(_0807_),
    .B1(_2779_),
    .X(_1840_));
 sky130_fd_sc_hd__a21o_1 _5103_ (.A1(net158),
    .A2(_0827_),
    .B1(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__nor2_1 _5104_ (.A(_2766_),
    .B(_1345_),
    .Y(_1842_));
 sky130_fd_sc_hd__or3_4 _5105_ (.A(_0825_),
    .B(_1841_),
    .C(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(net268),
    .A1(net348),
    .S(net134),
    .X(_1844_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(_1844_),
    .A1(\as2650.holding_reg[0] ),
    .S(_1843_),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_2 _5108_ (.A(_2652_),
    .B(net135),
    .Y(_1845_));
 sky130_fd_sc_hd__or2_1 _5109_ (.A(net264),
    .B(net134),
    .X(_1846_));
 sky130_fd_sc_hd__and2_1 _5110_ (.A(_1845_),
    .B(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(_1847_),
    .A1(\as2650.holding_reg[1] ),
    .S(_1843_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5112_ (.A0(net260),
    .A1(net344),
    .S(net134),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(_1848_),
    .A1(\as2650.holding_reg[2] ),
    .S(_1843_),
    .X(_0200_));
 sky130_fd_sc_hd__nor2_1 _5114_ (.A(net340),
    .B(net140),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(\as2650.r0[3] ),
    .B(net136),
    .Y(_1850_));
 sky130_fd_sc_hd__o21a_1 _5116_ (.A1(_2654_),
    .A2(net95),
    .B1(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__inv_2 _5117_ (.A(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(_1852_),
    .A1(\as2650.holding_reg[3] ),
    .S(_1843_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _5119_ (.A(net339),
    .B(net138),
    .Y(_1853_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(\as2650.r0[4] ),
    .B(net138),
    .Y(_1854_));
 sky130_fd_sc_hd__o21a_1 _5121_ (.A1(_2655_),
    .A2(net95),
    .B1(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__inv_2 _5122_ (.A(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(_1856_),
    .A1(\as2650.holding_reg[4] ),
    .S(_1843_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_2 _5124_ (.A0(net250),
    .A1(net337),
    .S(net134),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _5125_ (.A0(_1857_),
    .A1(\as2650.holding_reg[5] ),
    .S(_1843_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(net246),
    .A1(net335),
    .S(net133),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(_1858_),
    .A1(\as2650.holding_reg[6] ),
    .S(_1843_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5128_ (.A0(net242),
    .A1(net328),
    .S(net133),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(_1859_),
    .A1(\as2650.holding_reg[7] ),
    .S(_1843_),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _5130_ (.A1(net218),
    .A2(_0844_),
    .B1(net323),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_2638_),
    .B(net142),
    .Y(_1860_));
 sky130_fd_sc_hd__or2_4 _5132_ (.A(_1350_),
    .B(_1377_),
    .X(_1861_));
 sky130_fd_sc_hd__or2_4 _5133_ (.A(net89),
    .B(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__o211a_1 _5134_ (.A1(_2683_),
    .A2(_1860_),
    .B1(_1862_),
    .C1(_2677_),
    .X(_1863_));
 sky130_fd_sc_hd__a211o_1 _5135_ (.A1(net217),
    .A2(_2682_),
    .B1(_1403_),
    .C1(net97),
    .X(_1864_));
 sky130_fd_sc_hd__and3b_1 _5136_ (.A_N(_1863_),
    .B(_1864_),
    .C(net235),
    .X(_1865_));
 sky130_fd_sc_hd__or4_1 _5137_ (.A(net293),
    .B(net163),
    .C(net70),
    .D(_0753_),
    .X(_1866_));
 sky130_fd_sc_hd__or2_2 _5138_ (.A(_2937_),
    .B(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__a2bb2o_1 _5139_ (.A1_N(net147),
    .A2_N(_0836_),
    .B1(_1860_),
    .B2(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__o211ai_2 _5140_ (.A1(net142),
    .A2(_0743_),
    .B1(_0737_),
    .C1(_2638_),
    .Y(_1869_));
 sky130_fd_sc_hd__a21oi_2 _5141_ (.A1(_1868_),
    .A2(_1869_),
    .B1(net235),
    .Y(_1870_));
 sky130_fd_sc_hd__o32ai_4 _5142_ (.A1(_2726_),
    .A2(_1865_),
    .A3(_1870_),
    .B1(net145),
    .B2(_2638_),
    .Y(_1871_));
 sky130_fd_sc_hd__nor2_1 _5143_ (.A(_2710_),
    .B(_2764_),
    .Y(_1872_));
 sky130_fd_sc_hd__a21o_1 _5144_ (.A1(net309),
    .A2(net85),
    .B1(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__a21oi_1 _5145_ (.A1(net312),
    .A2(_2764_),
    .B1(_2737_),
    .Y(_1874_));
 sky130_fd_sc_hd__a211o_1 _5146_ (.A1(net293),
    .A2(_2710_),
    .B1(_1873_),
    .C1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__or4_1 _5147_ (.A(net148),
    .B(net136),
    .C(_1326_),
    .D(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(net96),
    .B(_0761_),
    .Y(_1877_));
 sky130_fd_sc_hd__a32o_1 _5149_ (.A1(_1344_),
    .A2(_1876_),
    .A3(_1877_),
    .B1(_1871_),
    .B2(net230),
    .X(_1878_));
 sky130_fd_sc_hd__o22a_1 _5150_ (.A1(net218),
    .A2(net217),
    .B1(_0843_),
    .B2(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__nor2_1 _5151_ (.A(net322),
    .B(_1879_),
    .Y(_0207_));
 sky130_fd_sc_hd__o21ai_1 _5152_ (.A1(net101),
    .A2(_0573_),
    .B1(net235),
    .Y(_1880_));
 sky130_fd_sc_hd__a211oi_1 _5153_ (.A1(net142),
    .A2(_1880_),
    .B1(_1817_),
    .C1(_2696_),
    .Y(_1881_));
 sky130_fd_sc_hd__a211oi_1 _5154_ (.A1(_0744_),
    .A2(_0830_),
    .B1(net213),
    .C1(_2726_),
    .Y(_1882_));
 sky130_fd_sc_hd__o221a_1 _5155_ (.A1(_2815_),
    .A2(_1867_),
    .B1(_1881_),
    .B2(_1348_),
    .C1(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__o21a_1 _5156_ (.A1(_1799_),
    .A2(_1862_),
    .B1(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__o21a_1 _5157_ (.A1(_1348_),
    .A2(_1873_),
    .B1(_2737_),
    .X(_1885_));
 sky130_fd_sc_hd__or4_1 _5158_ (.A(net136),
    .B(_0573_),
    .C(_1874_),
    .D(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__a311o_1 _5159_ (.A1(_1344_),
    .A2(_1877_),
    .A3(_1886_),
    .B1(net130),
    .C1(net295),
    .X(_1887_));
 sky130_fd_sc_hd__o2bb2a_1 _5160_ (.A1_N(net295),
    .A2_N(net292),
    .B1(_1884_),
    .B2(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__nor2_1 _5161_ (.A(net322),
    .B(_1888_),
    .Y(_0208_));
 sky130_fd_sc_hd__and3_2 _5162_ (.A(\as2650.cycle[2] ),
    .B(net291),
    .C(net293),
    .X(_1889_));
 sky130_fd_sc_hd__a21oi_2 _5163_ (.A1(net291),
    .A2(\as2650.cycle[0] ),
    .B1(net290),
    .Y(_1890_));
 sky130_fd_sc_hd__nor3_1 _5164_ (.A(net154),
    .B(_1889_),
    .C(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__or4_2 _5165_ (.A(net198),
    .B(_2765_),
    .C(_0807_),
    .D(_0827_),
    .X(_1892_));
 sky130_fd_sc_hd__nand2b_1 _5166_ (.A_N(_1891_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__a211o_1 _5167_ (.A1(net161),
    .A2(net71),
    .B1(_1889_),
    .C1(_1890_),
    .X(_1894_));
 sky130_fd_sc_hd__a31o_1 _5168_ (.A1(net297),
    .A2(_2694_),
    .A3(_2789_),
    .B1(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__nand3b_1 _5169_ (.A_N(_0836_),
    .B(_1894_),
    .C(_2694_),
    .Y(_1896_));
 sky130_fd_sc_hd__o2111ai_2 _5170_ (.A1(_2667_),
    .A2(_0738_),
    .B1(_1895_),
    .C1(_1896_),
    .D1(net216),
    .Y(_1897_));
 sky130_fd_sc_hd__o311a_1 _5171_ (.A1(net98),
    .A2(_2682_),
    .A3(_2703_),
    .B1(net77),
    .C1(_1891_),
    .X(_1898_));
 sky130_fd_sc_hd__nor2_1 _5172_ (.A(net98),
    .B(_1404_),
    .Y(_1899_));
 sky130_fd_sc_hd__o21ai_1 _5173_ (.A1(_2689_),
    .A2(net145),
    .B1(net235),
    .Y(_1900_));
 sky130_fd_sc_hd__o31a_1 _5174_ (.A1(_1898_),
    .A2(_1899_),
    .A3(_1900_),
    .B1(net69),
    .X(_1901_));
 sky130_fd_sc_hd__a221o_1 _5175_ (.A1(_2738_),
    .A2(_1893_),
    .B1(_1897_),
    .B2(_1901_),
    .C1(net295),
    .X(_1902_));
 sky130_fd_sc_hd__o211a_1 _5176_ (.A1(net218),
    .A2(net290),
    .B1(net316),
    .C1(_1902_),
    .X(_0209_));
 sky130_fd_sc_hd__o21ai_2 _5177_ (.A1(_2676_),
    .A2(_0576_),
    .B1(_2742_),
    .Y(_1903_));
 sky130_fd_sc_hd__nor2_1 _5178_ (.A(net289),
    .B(_1889_),
    .Y(_1904_));
 sky130_fd_sc_hd__and2_1 _5179_ (.A(net289),
    .B(_1889_),
    .X(_1905_));
 sky130_fd_sc_hd__or2_1 _5180_ (.A(_1904_),
    .B(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__a211oi_1 _5181_ (.A1(net235),
    .A2(_1903_),
    .B1(_1906_),
    .C1(net213),
    .Y(_1907_));
 sky130_fd_sc_hd__o211a_1 _5182_ (.A1(_2764_),
    .A2(_2783_),
    .B1(_1906_),
    .C1(net84),
    .X(_1908_));
 sky130_fd_sc_hd__o21a_1 _5183_ (.A1(net309),
    .A2(_2764_),
    .B1(net85),
    .X(_1909_));
 sky130_fd_sc_hd__o22a_1 _5184_ (.A1(_2737_),
    .A2(_2764_),
    .B1(_1908_),
    .B2(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__a2111o_1 _5185_ (.A1(net8),
    .A2(net79),
    .B1(_0573_),
    .C1(_1326_),
    .D1(net230),
    .X(_1911_));
 sky130_fd_sc_hd__nor2_1 _5186_ (.A(_1910_),
    .B(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__a32o_1 _5187_ (.A1(_2667_),
    .A2(net172),
    .A3(_1403_),
    .B1(_2741_),
    .B2(net8),
    .X(_1913_));
 sky130_fd_sc_hd__a211o_1 _5188_ (.A1(net173),
    .A2(_1913_),
    .B1(_1912_),
    .C1(net295),
    .X(_1914_));
 sky130_fd_sc_hd__o221a_1 _5189_ (.A1(net218),
    .A2(net289),
    .B1(_1907_),
    .B2(_1914_),
    .C1(net316),
    .X(_0210_));
 sky130_fd_sc_hd__a21oi_1 _5190_ (.A1(net218),
    .A2(_1905_),
    .B1(\as2650.cycle[4] ),
    .Y(_1915_));
 sky130_fd_sc_hd__and3_1 _5191_ (.A(net218),
    .B(\as2650.cycle[4] ),
    .C(_1905_),
    .X(_1916_));
 sky130_fd_sc_hd__nor3_1 _5192_ (.A(net322),
    .B(_1915_),
    .C(_1916_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _5193_ (.A1(\as2650.cycle[5] ),
    .A2(_1916_),
    .B1(net322),
    .Y(_1917_));
 sky130_fd_sc_hd__o21a_1 _5194_ (.A1(\as2650.cycle[5] ),
    .A2(_1916_),
    .B1(_1917_),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _5195_ (.A(\as2650.cycle[5] ),
    .B(\as2650.cycle[4] ),
    .C(_1905_),
    .X(_1918_));
 sky130_fd_sc_hd__and2_1 _5196_ (.A(\as2650.cycle[6] ),
    .B(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__or2_1 _5197_ (.A(\as2650.cycle[6] ),
    .B(_1918_),
    .X(_1920_));
 sky130_fd_sc_hd__a31o_1 _5198_ (.A1(_2737_),
    .A2(_2781_),
    .A3(_2783_),
    .B1(_2739_),
    .X(_1921_));
 sky130_fd_sc_hd__and3b_1 _5199_ (.A_N(_1919_),
    .B(_1920_),
    .C(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__a311o_1 _5200_ (.A1(net301),
    .A2(_2738_),
    .A3(_2826_),
    .B1(_1792_),
    .C1(net294),
    .X(_1923_));
 sky130_fd_sc_hd__o221a_1 _5201_ (.A1(net218),
    .A2(\as2650.cycle[6] ),
    .B1(_1922_),
    .B2(_1923_),
    .C1(net316),
    .X(_0213_));
 sky130_fd_sc_hd__xnor2_1 _5202_ (.A(\as2650.cycle[7] ),
    .B(_1919_),
    .Y(_1924_));
 sky130_fd_sc_hd__or4b_1 _5203_ (.A(net59),
    .B(_1924_),
    .C(_1795_),
    .D_N(_2740_),
    .X(_1925_));
 sky130_fd_sc_hd__a21oi_1 _5204_ (.A1(net235),
    .A2(net59),
    .B1(net294),
    .Y(_1926_));
 sky130_fd_sc_hd__a221oi_2 _5205_ (.A1(net294),
    .A2(_2637_),
    .B1(_1925_),
    .B2(_1926_),
    .C1(net322),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_0832_),
    .B(_0841_),
    .Y(_1927_));
 sky130_fd_sc_hd__mux2_1 _5207_ (.A0(\as2650.psu[7] ),
    .A1(_0775_),
    .S(net331),
    .X(_1928_));
 sky130_fd_sc_hd__o22a_1 _5208_ (.A1(net239),
    .A2(_0832_),
    .B1(_1927_),
    .B2(\as2650.sense ),
    .X(_1929_));
 sky130_fd_sc_hd__o21a_1 _5209_ (.A1(_0841_),
    .A2(_1928_),
    .B1(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__or2_1 _5210_ (.A(\as2650.psu[7] ),
    .B(_2636_),
    .X(_1931_));
 sky130_fd_sc_hd__o211a_1 _5211_ (.A1(net296),
    .A2(_1930_),
    .B1(_1931_),
    .C1(net320),
    .X(_0215_));
 sky130_fd_sc_hd__o221a_1 _5212_ (.A1(net349),
    .A2(net149),
    .B1(_2692_),
    .B2(net310),
    .C1(net159),
    .X(_1932_));
 sky130_fd_sc_hd__mux2_2 _5213_ (.A0(net286),
    .A1(_1389_),
    .S(net312),
    .X(_1933_));
 sky130_fd_sc_hd__inv_2 _5214_ (.A(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__nand2_1 _5215_ (.A(net286),
    .B(net301),
    .Y(_1935_));
 sky130_fd_sc_hd__o211a_1 _5216_ (.A1(net301),
    .A2(_1933_),
    .B1(_1935_),
    .C1(net160),
    .X(_1936_));
 sky130_fd_sc_hd__nor2_1 _5217_ (.A(_1932_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__or2_2 _5218_ (.A(net286),
    .B(net301),
    .X(_1938_));
 sky130_fd_sc_hd__and2_1 _5219_ (.A(_1935_),
    .B(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(net287),
    .A1(_1939_),
    .S(_1376_),
    .X(_1940_));
 sky130_fd_sc_hd__nor2_1 _5221_ (.A(_2635_),
    .B(_1350_),
    .Y(_1941_));
 sky130_fd_sc_hd__a221o_1 _5222_ (.A1(net232),
    .A2(net298),
    .B1(_1350_),
    .B2(_1939_),
    .C1(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__o211a_1 _5223_ (.A1(_2769_),
    .A2(_1940_),
    .B1(_1942_),
    .C1(net137),
    .X(_1943_));
 sky130_fd_sc_hd__a211o_1 _5224_ (.A1(net132),
    .A2(_1937_),
    .B1(_1943_),
    .C1(net100),
    .X(_1944_));
 sky130_fd_sc_hd__a21oi_1 _5225_ (.A1(net155),
    .A2(_2873_),
    .B1(net347),
    .Y(_1945_));
 sky130_fd_sc_hd__and3_1 _5226_ (.A(net347),
    .B(net155),
    .C(_2873_),
    .X(_1946_));
 sky130_fd_sc_hd__nor2_4 _5227_ (.A(net97),
    .B(net143),
    .Y(_1947_));
 sky130_fd_sc_hd__o21a_1 _5228_ (.A1(_1945_),
    .A2(_1946_),
    .B1(net141),
    .X(_1948_));
 sky130_fd_sc_hd__a211o_1 _5229_ (.A1(net288),
    .A2(net143),
    .B1(_1948_),
    .C1(net97),
    .X(_1949_));
 sky130_fd_sc_hd__o221a_1 _5230_ (.A1(net287),
    .A2(_2827_),
    .B1(_1394_),
    .B2(_1934_),
    .C1(_0580_),
    .X(_1950_));
 sky130_fd_sc_hd__a31o_1 _5231_ (.A1(net145),
    .A2(_1944_),
    .A3(_1949_),
    .B1(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__o22a_1 _5232_ (.A1(\as2650.stack[3][0] ),
    .A2(net193),
    .B1(net189),
    .B2(\as2650.stack[2][0] ),
    .X(_1952_));
 sky130_fd_sc_hd__o221a_2 _5233_ (.A1(\as2650.stack[0][0] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][0] ),
    .C1(_2859_),
    .X(_1953_));
 sky130_fd_sc_hd__mux4_2 _5234_ (.A0(\as2650.stack[7][0] ),
    .A1(\as2650.stack[4][0] ),
    .A2(\as2650.stack[5][0] ),
    .A3(\as2650.stack[6][0] ),
    .S0(net224),
    .S1(net225),
    .X(_1954_));
 sky130_fd_sc_hd__a22oi_4 _5235_ (.A1(_1952_),
    .A2(_1953_),
    .B1(_1954_),
    .B2(net122),
    .Y(_1955_));
 sky130_fd_sc_hd__inv_2 _5236_ (.A(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__o221a_1 _5237_ (.A1(net287),
    .A2(_0815_),
    .B1(net103),
    .B2(_1955_),
    .C1(_1951_),
    .X(_1957_));
 sky130_fd_sc_hd__or3_1 _5238_ (.A(net101),
    .B(_2686_),
    .C(net154),
    .X(_1958_));
 sky130_fd_sc_hd__or4_1 _5239_ (.A(net210),
    .B(_2668_),
    .C(net146),
    .D(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__o311a_1 _5240_ (.A1(_2637_),
    .A2(\as2650.cycle[6] ),
    .A3(net229),
    .B1(_2728_),
    .C1(_2733_),
    .X(_1960_));
 sky130_fd_sc_hd__and3_1 _5241_ (.A(net95),
    .B(_0761_),
    .C(_1349_),
    .X(_1961_));
 sky130_fd_sc_hd__inv_2 _5242_ (.A(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a21o_1 _5243_ (.A1(_0576_),
    .A2(_1836_),
    .B1(_2739_),
    .X(_1963_));
 sky130_fd_sc_hd__and3_1 _5244_ (.A(net172),
    .B(_2688_),
    .C(net64),
    .X(_1964_));
 sky130_fd_sc_hd__a31o_1 _5245_ (.A1(net238),
    .A2(net172),
    .A3(_1403_),
    .B1(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__a21oi_1 _5246_ (.A1(net173),
    .A2(_1965_),
    .B1(_1820_),
    .Y(_1966_));
 sky130_fd_sc_hd__a211o_1 _5247_ (.A1(net136),
    .A2(_2790_),
    .B1(_0746_),
    .C1(_0760_),
    .X(_1967_));
 sky130_fd_sc_hd__and4_1 _5248_ (.A(_1359_),
    .B(_1959_),
    .C(_1962_),
    .D(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__and4b_1 _5249_ (.A_N(_1899_),
    .B(_1960_),
    .C(_1968_),
    .D(_1803_),
    .X(_1969_));
 sky130_fd_sc_hd__and4_4 _5250_ (.A(_1790_),
    .B(_1963_),
    .C(_1966_),
    .D(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__clkinv_4 _5251_ (.A(net45),
    .Y(_1971_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(net287),
    .A1(_1957_),
    .S(net68),
    .X(_1972_));
 sky130_fd_sc_hd__o21ai_1 _5253_ (.A1(net287),
    .A2(net46),
    .B1(net317),
    .Y(_1973_));
 sky130_fd_sc_hd__a21oi_1 _5254_ (.A1(net46),
    .A2(_1972_),
    .B1(_1973_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_2 _5255_ (.A(net285),
    .B(net286),
    .Y(_1974_));
 sky130_fd_sc_hd__or2_1 _5256_ (.A(net285),
    .B(net287),
    .X(_1975_));
 sky130_fd_sc_hd__nand2_2 _5257_ (.A(_1974_),
    .B(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__nor2_1 _5258_ (.A(net293),
    .B(net99),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5259_ (.A(net285),
    .B(_1938_),
    .Y(_1978_));
 sky130_fd_sc_hd__o21ai_1 _5260_ (.A1(net303),
    .A2(_1975_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__nand2_2 _5261_ (.A(net345),
    .B(net150),
    .Y(_1980_));
 sky130_fd_sc_hd__and2_2 _5262_ (.A(net345),
    .B(_2885_),
    .X(_1981_));
 sky130_fd_sc_hd__xnor2_4 _5263_ (.A(net345),
    .B(_2885_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand2_2 _5264_ (.A(net348),
    .B(_2873_),
    .Y(_1983_));
 sky130_fd_sc_hd__nor2_4 _5265_ (.A(_1982_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__a21o_1 _5266_ (.A1(_1982_),
    .A2(_1983_),
    .B1(net150),
    .X(_1985_));
 sky130_fd_sc_hd__o211ai_4 _5267_ (.A1(_1984_),
    .A2(_1985_),
    .B1(_2680_),
    .C1(_1980_),
    .Y(_1986_));
 sky130_fd_sc_hd__mux2_2 _5268_ (.A0(net284),
    .A1(_1432_),
    .S(net312),
    .X(_1987_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(net346),
    .A1(\as2650.addr_buff[1] ),
    .S(net147),
    .X(_1988_));
 sky130_fd_sc_hd__a2bb2o_1 _5270_ (.A1_N(net63),
    .A2_N(_1976_),
    .B1(_1988_),
    .B2(net157),
    .X(_1989_));
 sky130_fd_sc_hd__a211o_1 _5271_ (.A1(_2741_),
    .A2(_1987_),
    .B1(_1989_),
    .C1(net99),
    .X(_1990_));
 sky130_fd_sc_hd__a21oi_1 _5272_ (.A1(_1986_),
    .A2(_1990_),
    .B1(net93),
    .Y(_1991_));
 sky130_fd_sc_hd__o21a_2 _5273_ (.A1(net293),
    .A2(_1861_),
    .B1(net97),
    .X(_1992_));
 sky130_fd_sc_hd__inv_2 _5274_ (.A(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__a32o_1 _5275_ (.A1(_1861_),
    .A2(_1977_),
    .A3(_1979_),
    .B1(_1993_),
    .B2(_1976_),
    .X(_1994_));
 sky130_fd_sc_hd__a211o_1 _5276_ (.A1(net143),
    .A2(_1994_),
    .B1(_1991_),
    .C1(net72),
    .X(_1995_));
 sky130_fd_sc_hd__and3_1 _5277_ (.A(net227),
    .B(\as2650.stack[3][1] ),
    .C(net195),
    .X(_1996_));
 sky130_fd_sc_hd__o22a_1 _5278_ (.A1(\as2650.stack[0][1] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][1] ),
    .X(_1997_));
 sky130_fd_sc_hd__o221a_2 _5279_ (.A1(\as2650.stack[2][1] ),
    .A2(net189),
    .B1(_1996_),
    .B2(_2849_),
    .C1(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__o22a_1 _5280_ (.A1(\as2650.stack[7][1] ),
    .A2(net193),
    .B1(net190),
    .B2(\as2650.stack[6][1] ),
    .X(_1999_));
 sky130_fd_sc_hd__o22a_1 _5281_ (.A1(\as2650.stack[4][1] ),
    .A2(net170),
    .B1(net166),
    .B2(\as2650.stack[5][1] ),
    .X(_2000_));
 sky130_fd_sc_hd__a31o_4 _5282_ (.A1(net122),
    .A2(_1999_),
    .A3(_2000_),
    .B1(_1998_),
    .X(_2001_));
 sky130_fd_sc_hd__inv_2 _5283_ (.A(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nor2_1 _5284_ (.A(net93),
    .B(_1987_),
    .Y(_2003_));
 sky130_fd_sc_hd__a211o_1 _5285_ (.A1(net93),
    .A2(_1976_),
    .B1(_2003_),
    .C1(net144),
    .X(_2004_));
 sky130_fd_sc_hd__o221a_1 _5286_ (.A1(_0815_),
    .A2(_1976_),
    .B1(_2002_),
    .B2(net102),
    .C1(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__a21oi_1 _5287_ (.A1(_1995_),
    .A2(_2005_),
    .B1(net65),
    .Y(_2006_));
 sky130_fd_sc_hd__o21ai_1 _5288_ (.A1(net67),
    .A2(_1976_),
    .B1(_1970_),
    .Y(_2007_));
 sky130_fd_sc_hd__o221a_1 _5289_ (.A1(net285),
    .A2(net45),
    .B1(_2006_),
    .B2(_2007_),
    .C1(net319),
    .X(_0217_));
 sky130_fd_sc_hd__nand2_4 _5290_ (.A(net93),
    .B(_1861_),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2_4 _5291_ (.A(net99),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__and3_1 _5292_ (.A(\as2650.pc[2] ),
    .B(net285),
    .C(_1938_),
    .X(_2010_));
 sky130_fd_sc_hd__a21oi_1 _5293_ (.A1(net285),
    .A2(_1938_),
    .B1(\as2650.pc[2] ),
    .Y(_2011_));
 sky130_fd_sc_hd__o21ai_1 _5294_ (.A1(_2010_),
    .A2(_2011_),
    .B1(_2009_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand2_4 _5295_ (.A(net343),
    .B(_2948_),
    .Y(_2013_));
 sky130_fd_sc_hd__or2_2 _5296_ (.A(net343),
    .B(_2948_),
    .X(_2014_));
 sky130_fd_sc_hd__o211ai_4 _5297_ (.A1(_1981_),
    .A2(_1984_),
    .B1(_2013_),
    .C1(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__a211o_1 _5298_ (.A1(_2013_),
    .A2(_2014_),
    .B1(_1981_),
    .C1(_1984_),
    .X(_2016_));
 sky130_fd_sc_hd__a21oi_2 _5299_ (.A1(_2015_),
    .A2(_2016_),
    .B1(net150),
    .Y(_2017_));
 sky130_fd_sc_hd__a21oi_2 _5300_ (.A1(_2653_),
    .A2(net147),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__mux2_2 _5301_ (.A0(_2634_),
    .A1(_1466_),
    .S(net311),
    .X(_2019_));
 sky130_fd_sc_hd__nor2_1 _5302_ (.A(net77),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net342),
    .A1(\as2650.addr_buff[2] ),
    .S(net147),
    .X(_2021_));
 sky130_fd_sc_hd__nor2_1 _5304_ (.A(_2634_),
    .B(_1974_),
    .Y(_2022_));
 sky130_fd_sc_hd__and2_1 _5305_ (.A(_2634_),
    .B(_1974_),
    .X(_2023_));
 sky130_fd_sc_hd__nor2_2 _5306_ (.A(_2022_),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__a221o_1 _5307_ (.A1(net157),
    .A2(_2021_),
    .B1(_2024_),
    .B2(_1396_),
    .C1(net100),
    .X(_2025_));
 sky130_fd_sc_hd__o22a_1 _5308_ (.A1(_2681_),
    .A2(_2018_),
    .B1(_2020_),
    .B2(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__o21a_1 _5309_ (.A1(net92),
    .A2(_2026_),
    .B1(net144),
    .X(_2027_));
 sky130_fd_sc_hd__nor2_4 _5310_ (.A(net141),
    .B(_1992_),
    .Y(_2028_));
 sky130_fd_sc_hd__or2_4 _5311_ (.A(net141),
    .B(_1992_),
    .X(_2029_));
 sky130_fd_sc_hd__or2_1 _5312_ (.A(_2024_),
    .B(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__o21ai_1 _5313_ (.A1(_2827_),
    .A2(_2024_),
    .B1(net72),
    .Y(_2031_));
 sky130_fd_sc_hd__a21oi_1 _5314_ (.A1(_1393_),
    .A2(_2019_),
    .B1(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__a31o_1 _5315_ (.A1(_2012_),
    .A2(_2027_),
    .A3(_2030_),
    .B1(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__and3_1 _5316_ (.A(net227),
    .B(\as2650.stack[3][2] ),
    .C(net195),
    .X(_2034_));
 sky130_fd_sc_hd__o22a_1 _5317_ (.A1(\as2650.stack[0][2] ),
    .A2(net168),
    .B1(net167),
    .B2(\as2650.stack[1][2] ),
    .X(_2035_));
 sky130_fd_sc_hd__o221a_1 _5318_ (.A1(\as2650.stack[2][2] ),
    .A2(net189),
    .B1(_2034_),
    .B2(_2849_),
    .C1(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__o22a_1 _5319_ (.A1(\as2650.stack[5][2] ),
    .A2(net167),
    .B1(net190),
    .B2(\as2650.stack[6][2] ),
    .X(_2037_));
 sky130_fd_sc_hd__o22a_1 _5320_ (.A1(\as2650.stack[7][2] ),
    .A2(net193),
    .B1(_2852_),
    .B2(\as2650.stack[4][2] ),
    .X(_2038_));
 sky130_fd_sc_hd__a31o_4 _5321_ (.A1(net122),
    .A2(_2037_),
    .A3(_2038_),
    .B1(_2036_),
    .X(_2039_));
 sky130_fd_sc_hd__o221a_1 _5322_ (.A1(net104),
    .A2(_2024_),
    .B1(_2039_),
    .B2(net102),
    .C1(net67),
    .X(_2040_));
 sky130_fd_sc_hd__a221o_1 _5323_ (.A1(net66),
    .A2(_2024_),
    .B1(_2033_),
    .B2(_2040_),
    .C1(_1971_),
    .X(_2041_));
 sky130_fd_sc_hd__o211a_1 _5324_ (.A1(\as2650.pc[2] ),
    .A2(net46),
    .B1(_2041_),
    .C1(net315),
    .X(_0218_));
 sky130_fd_sc_hd__and2_2 _5325_ (.A(net283),
    .B(_2010_),
    .X(_2042_));
 sky130_fd_sc_hd__nor2_1 _5326_ (.A(\as2650.pc[3] ),
    .B(_2010_),
    .Y(_2043_));
 sky130_fd_sc_hd__or3_1 _5327_ (.A(_2008_),
    .B(_2042_),
    .C(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(\as2650.pc[3] ),
    .A1(_1507_),
    .S(net312),
    .X(_2045_));
 sky130_fd_sc_hd__inv_2 _5329_ (.A(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _5330_ (.A(\as2650.addr_buff[3] ),
    .B(net149),
    .Y(_2047_));
 sky130_fd_sc_hd__o211a_1 _5331_ (.A1(_2654_),
    .A2(net149),
    .B1(_2047_),
    .C1(net157),
    .X(_2048_));
 sky130_fd_sc_hd__and2_4 _5332_ (.A(net283),
    .B(_2022_),
    .X(_2049_));
 sky130_fd_sc_hd__nor2_1 _5333_ (.A(net283),
    .B(_2022_),
    .Y(_2050_));
 sky130_fd_sc_hd__or2_4 _5334_ (.A(_2049_),
    .B(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__a211o_1 _5335_ (.A1(_1396_),
    .A2(_2051_),
    .B1(_2048_),
    .C1(net94),
    .X(_2052_));
 sky130_fd_sc_hd__a21o_1 _5336_ (.A1(_2741_),
    .A2(_2046_),
    .B1(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__o211a_1 _5337_ (.A1(_1862_),
    .A2(_2051_),
    .B1(_2053_),
    .C1(net172),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _5338_ (.A(_2044_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__o221a_1 _5339_ (.A1(_1394_),
    .A2(_2046_),
    .B1(_2051_),
    .B2(_2827_),
    .C1(net72),
    .X(_2056_));
 sky130_fd_sc_hd__and2_2 _5340_ (.A(net341),
    .B(_0303_),
    .X(_2057_));
 sky130_fd_sc_hd__nor2_2 _5341_ (.A(net341),
    .B(_0303_),
    .Y(_2058_));
 sky130_fd_sc_hd__o211a_1 _5342_ (.A1(_2057_),
    .A2(_2058_),
    .B1(_2013_),
    .C1(_2015_),
    .X(_2059_));
 sky130_fd_sc_hd__a211oi_4 _5343_ (.A1(_2013_),
    .A2(_2015_),
    .B1(_2057_),
    .C1(_2058_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(net341),
    .B(net150),
    .Y(_2061_));
 sky130_fd_sc_hd__o311a_2 _5345_ (.A1(net150),
    .A2(_2059_),
    .A3(_2060_),
    .B1(_2061_),
    .C1(_1947_),
    .X(_2062_));
 sky130_fd_sc_hd__a31o_1 _5346_ (.A1(net99),
    .A2(net143),
    .A3(_2051_),
    .B1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__or3b_2 _5347_ (.A(_2063_),
    .B(_2056_),
    .C_N(_2055_),
    .X(_2064_));
 sky130_fd_sc_hd__o22a_1 _5348_ (.A1(\as2650.stack[7][3] ),
    .A2(net193),
    .B1(net190),
    .B2(\as2650.stack[6][3] ),
    .X(_2065_));
 sky130_fd_sc_hd__o221a_1 _5349_ (.A1(\as2650.stack[4][3] ),
    .A2(net168),
    .B1(net167),
    .B2(\as2650.stack[5][3] ),
    .C1(net122),
    .X(_2066_));
 sky130_fd_sc_hd__o22a_1 _5350_ (.A1(\as2650.stack[3][3] ),
    .A2(net193),
    .B1(net189),
    .B2(\as2650.stack[2][3] ),
    .X(_2067_));
 sky130_fd_sc_hd__o221a_2 _5351_ (.A1(\as2650.stack[0][3] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][3] ),
    .C1(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__a22o_4 _5352_ (.A1(_2065_),
    .A2(_2066_),
    .B1(_2068_),
    .B2(_2859_),
    .X(_2069_));
 sky130_fd_sc_hd__inv_2 _5353_ (.A(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__nor2_1 _5354_ (.A(net67),
    .B(_2051_),
    .Y(_2071_));
 sky130_fd_sc_hd__o221a_1 _5355_ (.A1(net104),
    .A2(_2051_),
    .B1(_2070_),
    .B2(net102),
    .C1(_2064_),
    .X(_2072_));
 sky130_fd_sc_hd__o21ai_1 _5356_ (.A1(net65),
    .A2(_2072_),
    .B1(net46),
    .Y(_2073_));
 sky130_fd_sc_hd__o221a_1 _5357_ (.A1(net283),
    .A2(net46),
    .B1(_2071_),
    .B2(_2073_),
    .C1(net315),
    .X(_0219_));
 sky130_fd_sc_hd__xnor2_4 _5358_ (.A(net281),
    .B(_2049_),
    .Y(_2074_));
 sky130_fd_sc_hd__mux2_2 _5359_ (.A0(_2632_),
    .A1(_1543_),
    .S(net311),
    .X(_2075_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(net338),
    .A1(\as2650.addr_buff[4] ),
    .S(net147),
    .X(_2076_));
 sky130_fd_sc_hd__inv_2 _5361_ (.A(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__o221a_1 _5362_ (.A1(_1397_),
    .A2(_2074_),
    .B1(_2077_),
    .B2(net160),
    .C1(net97),
    .X(_2078_));
 sky130_fd_sc_hd__o21a_1 _5363_ (.A1(net77),
    .A2(_2075_),
    .B1(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(net338),
    .B(net152),
    .Y(_2080_));
 sky130_fd_sc_hd__and2_1 _5365_ (.A(net338),
    .B(_0347_),
    .X(_2081_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(net338),
    .B(_0347_),
    .Y(_2082_));
 sky130_fd_sc_hd__or2_1 _5367_ (.A(net338),
    .B(_0347_),
    .X(_2083_));
 sky130_fd_sc_hd__a211o_1 _5368_ (.A1(_2082_),
    .A2(_2083_),
    .B1(_2057_),
    .C1(_2060_),
    .X(_2084_));
 sky130_fd_sc_hd__o211a_1 _5369_ (.A1(_2057_),
    .A2(_2060_),
    .B1(_2082_),
    .C1(_2083_),
    .X(_2085_));
 sky130_fd_sc_hd__or3b_2 _5370_ (.A(_2085_),
    .B(net150),
    .C_N(_2084_),
    .X(_2086_));
 sky130_fd_sc_hd__a31o_1 _5371_ (.A1(_2680_),
    .A2(_2080_),
    .A3(_2086_),
    .B1(_2079_),
    .X(_2087_));
 sky130_fd_sc_hd__o221a_1 _5372_ (.A1(_2827_),
    .A2(_2074_),
    .B1(_2075_),
    .B2(_1394_),
    .C1(net72),
    .X(_2088_));
 sky130_fd_sc_hd__a21o_1 _5373_ (.A1(_2702_),
    .A2(_2087_),
    .B1(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__xnor2_1 _5374_ (.A(net282),
    .B(_2042_),
    .Y(_2090_));
 sky130_fd_sc_hd__a31o_1 _5375_ (.A1(net144),
    .A2(_2009_),
    .A3(_2090_),
    .B1(_2089_),
    .X(_2091_));
 sky130_fd_sc_hd__a22o_1 _5376_ (.A1(_2028_),
    .A2(_2074_),
    .B1(_2091_),
    .B2(net67),
    .X(_2092_));
 sky130_fd_sc_hd__mux4_2 _5377_ (.A0(\as2650.stack[7][4] ),
    .A1(\as2650.stack[4][4] ),
    .A2(\as2650.stack[5][4] ),
    .A3(\as2650.stack[6][4] ),
    .S0(net224),
    .S1(net225),
    .X(_2093_));
 sky130_fd_sc_hd__o22a_2 _5378_ (.A1(\as2650.stack[3][4] ),
    .A2(net193),
    .B1(net189),
    .B2(\as2650.stack[2][4] ),
    .X(_2094_));
 sky130_fd_sc_hd__o221a_2 _5379_ (.A1(\as2650.stack[0][4] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][4] ),
    .C1(_2859_),
    .X(_2095_));
 sky130_fd_sc_hd__a22oi_4 _5380_ (.A1(net122),
    .A2(_2093_),
    .B1(_2094_),
    .B2(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__o21a_1 _5381_ (.A1(net102),
    .A2(_2096_),
    .B1(_2092_),
    .X(_2097_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(net66),
    .A2(_2074_),
    .B1(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__o21ai_1 _5383_ (.A1(net104),
    .A2(_2074_),
    .B1(net45),
    .Y(_2099_));
 sky130_fd_sc_hd__o221a_1 _5384_ (.A1(net282),
    .A2(net45),
    .B1(_2098_),
    .B2(_2099_),
    .C1(net315),
    .X(_0220_));
 sky130_fd_sc_hd__and3_2 _5385_ (.A(net279),
    .B(net282),
    .C(_2042_),
    .X(_2100_));
 sky130_fd_sc_hd__a21oi_1 _5386_ (.A1(net282),
    .A2(_2042_),
    .B1(net280),
    .Y(_2101_));
 sky130_fd_sc_hd__and3_2 _5387_ (.A(net280),
    .B(net282),
    .C(_2049_),
    .X(_2102_));
 sky130_fd_sc_hd__a21oi_2 _5388_ (.A1(net282),
    .A2(_2049_),
    .B1(net280),
    .Y(_2103_));
 sky130_fd_sc_hd__nor2_4 _5389_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__nand2_2 _5390_ (.A(net336),
    .B(_0394_),
    .Y(_2105_));
 sky130_fd_sc_hd__inv_2 _5391_ (.A(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__or2_1 _5392_ (.A(net336),
    .B(_0394_),
    .X(_2107_));
 sky130_fd_sc_hd__o211a_1 _5393_ (.A1(_2081_),
    .A2(_2085_),
    .B1(_2105_),
    .C1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__a211oi_1 _5394_ (.A1(_2105_),
    .A2(_2107_),
    .B1(_2081_),
    .C1(_2085_),
    .Y(_2109_));
 sky130_fd_sc_hd__o21ai_1 _5395_ (.A1(_2108_),
    .A2(_2109_),
    .B1(net155),
    .Y(_2110_));
 sky130_fd_sc_hd__o211a_1 _5396_ (.A1(net336),
    .A2(net155),
    .B1(_1947_),
    .C1(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(net279),
    .A1(_1579_),
    .S(net311),
    .X(_2112_));
 sky130_fd_sc_hd__a221o_1 _5398_ (.A1(net337),
    .A2(net153),
    .B1(net147),
    .B2(\as2650.addr_buff[5] ),
    .C1(net160),
    .X(_2113_));
 sky130_fd_sc_hd__o211a_1 _5399_ (.A1(net63),
    .A2(_2104_),
    .B1(_2113_),
    .C1(net89),
    .X(_2114_));
 sky130_fd_sc_hd__o21ai_1 _5400_ (.A1(net77),
    .A2(_2112_),
    .B1(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__o31a_1 _5401_ (.A1(_2008_),
    .A2(_2100_),
    .A3(_2101_),
    .B1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__a2bb2o_1 _5402_ (.A1_N(net99),
    .A2_N(_2116_),
    .B1(_2104_),
    .B2(_2028_),
    .X(_2117_));
 sky130_fd_sc_hd__or3_1 _5403_ (.A(net146),
    .B(_2111_),
    .C(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__a221o_1 _5404_ (.A1(_2826_),
    .A2(_2104_),
    .B1(_2112_),
    .B2(net64),
    .C1(_0579_),
    .X(_2119_));
 sky130_fd_sc_hd__and3_1 _5405_ (.A(net227),
    .B(\as2650.stack[3][5] ),
    .C(net195),
    .X(_2120_));
 sky130_fd_sc_hd__o22a_1 _5406_ (.A1(\as2650.stack[0][5] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][5] ),
    .X(_2121_));
 sky130_fd_sc_hd__o221a_1 _5407_ (.A1(\as2650.stack[2][5] ),
    .A2(net189),
    .B1(_2120_),
    .B2(_2849_),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__mux4_2 _5408_ (.A0(\as2650.stack[7][5] ),
    .A1(\as2650.stack[4][5] ),
    .A2(\as2650.stack[5][5] ),
    .A3(\as2650.stack[6][5] ),
    .S0(net224),
    .S1(net225),
    .X(_2123_));
 sky130_fd_sc_hd__a21o_2 _5409_ (.A1(net122),
    .A2(_2123_),
    .B1(_2122_),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _5410_ (.A1(_0814_),
    .A2(_2104_),
    .B1(_2124_),
    .B2(_0830_),
    .X(_2125_));
 sky130_fd_sc_hd__a21oi_1 _5411_ (.A1(_2118_),
    .A2(_2119_),
    .B1(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__nor2_1 _5412_ (.A(net66),
    .B(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__a211o_1 _5413_ (.A1(net65),
    .A2(_2104_),
    .B1(_2127_),
    .C1(_1971_),
    .X(_2128_));
 sky130_fd_sc_hd__o211a_1 _5414_ (.A1(net279),
    .A2(net46),
    .B1(_2128_),
    .C1(net315),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(net277),
    .B(_2100_),
    .Y(_2129_));
 sky130_fd_sc_hd__or2_1 _5416_ (.A(net277),
    .B(_2100_),
    .X(_2130_));
 sky130_fd_sc_hd__a211o_1 _5417_ (.A1(_2129_),
    .A2(_2130_),
    .B1(net99),
    .C1(_2008_),
    .X(_2131_));
 sky130_fd_sc_hd__mux2_4 _5418_ (.A0(net278),
    .A1(_1616_),
    .S(net311),
    .X(_2132_));
 sky130_fd_sc_hd__and2_4 _5419_ (.A(net277),
    .B(_2102_),
    .X(_2133_));
 sky130_fd_sc_hd__nor2_1 _5420_ (.A(\as2650.pc[6] ),
    .B(_2102_),
    .Y(_2134_));
 sky130_fd_sc_hd__nor2_2 _5421_ (.A(_2133_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(\as2650.addr_buff[6] ),
    .A1(net334),
    .S(_2692_),
    .X(_2136_));
 sky130_fd_sc_hd__a221o_1 _5423_ (.A1(_1396_),
    .A2(_2135_),
    .B1(_2136_),
    .B2(net157),
    .C1(net99),
    .X(_2137_));
 sky130_fd_sc_hd__a21oi_1 _5424_ (.A1(_2741_),
    .A2(_2132_),
    .B1(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(net334),
    .B(net150),
    .Y(_2139_));
 sky130_fd_sc_hd__and2_1 _5426_ (.A(net334),
    .B(_0458_),
    .X(_2140_));
 sky130_fd_sc_hd__inv_2 _5427_ (.A(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__or2_1 _5428_ (.A(net334),
    .B(_0458_),
    .X(_2142_));
 sky130_fd_sc_hd__a211oi_1 _5429_ (.A1(_2141_),
    .A2(_2142_),
    .B1(_2106_),
    .C1(_2108_),
    .Y(_2143_));
 sky130_fd_sc_hd__o211a_1 _5430_ (.A1(_2106_),
    .A2(_2108_),
    .B1(_2141_),
    .C1(_2142_),
    .X(_2144_));
 sky130_fd_sc_hd__o311a_1 _5431_ (.A1(_2693_),
    .A2(_2143_),
    .A3(_2144_),
    .B1(_2139_),
    .C1(_2680_),
    .X(_2145_));
 sky130_fd_sc_hd__o21ai_1 _5432_ (.A1(_2138_),
    .A2(_2145_),
    .B1(net90),
    .Y(_2146_));
 sky130_fd_sc_hd__o211a_1 _5433_ (.A1(_2029_),
    .A2(_2135_),
    .B1(_2131_),
    .C1(net144),
    .X(_2147_));
 sky130_fd_sc_hd__o221a_1 _5434_ (.A1(_1394_),
    .A2(_2132_),
    .B1(_2135_),
    .B2(_2827_),
    .C1(net72),
    .X(_2148_));
 sky130_fd_sc_hd__a21o_1 _5435_ (.A1(_2146_),
    .A2(_2147_),
    .B1(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__and3_1 _5436_ (.A(net227),
    .B(\as2650.stack[3][6] ),
    .C(net195),
    .X(_2150_));
 sky130_fd_sc_hd__o22a_1 _5437_ (.A1(\as2650.stack[0][6] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][6] ),
    .X(_2151_));
 sky130_fd_sc_hd__o221a_2 _5438_ (.A1(\as2650.stack[2][6] ),
    .A2(net189),
    .B1(_2150_),
    .B2(_2849_),
    .C1(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__o22a_1 _5439_ (.A1(\as2650.stack[7][6] ),
    .A2(net194),
    .B1(net191),
    .B2(\as2650.stack[6][6] ),
    .X(_2153_));
 sky130_fd_sc_hd__o22a_1 _5440_ (.A1(\as2650.stack[4][6] ),
    .A2(net170),
    .B1(net166),
    .B2(\as2650.stack[5][6] ),
    .X(_2154_));
 sky130_fd_sc_hd__a31o_4 _5441_ (.A1(net122),
    .A2(_2153_),
    .A3(_2154_),
    .B1(_2152_),
    .X(_2155_));
 sky130_fd_sc_hd__or2_1 _5442_ (.A(net102),
    .B(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__o211a_1 _5443_ (.A1(net104),
    .A2(_2135_),
    .B1(_2156_),
    .C1(net68),
    .X(_2157_));
 sky130_fd_sc_hd__a221o_1 _5444_ (.A1(net65),
    .A2(_2135_),
    .B1(_2149_),
    .B2(_2157_),
    .C1(_1971_),
    .X(_2158_));
 sky130_fd_sc_hd__o211a_1 _5445_ (.A1(net278),
    .A2(net45),
    .B1(_2158_),
    .C1(net319),
    .X(_0222_));
 sky130_fd_sc_hd__and3_2 _5446_ (.A(net276),
    .B(net277),
    .C(_2100_),
    .X(_2159_));
 sky130_fd_sc_hd__a21oi_1 _5447_ (.A1(net278),
    .A2(_2100_),
    .B1(net276),
    .Y(_2160_));
 sky130_fd_sc_hd__xnor2_4 _5448_ (.A(net276),
    .B(_2133_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(net330),
    .B(_2891_),
    .Y(_2162_));
 sky130_fd_sc_hd__or2_1 _5450_ (.A(net330),
    .B(_2891_),
    .X(_2163_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_2162_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__nor2_1 _5452_ (.A(_2140_),
    .B(_2144_),
    .Y(_2165_));
 sky130_fd_sc_hd__xnor2_1 _5453_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__nor2_1 _5454_ (.A(net329),
    .B(net155),
    .Y(_2167_));
 sky130_fd_sc_hd__mux2_2 _5455_ (.A0(net276),
    .A1(_1648_),
    .S(net311),
    .X(_2168_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(\as2650.addr_buff[7] ),
    .A1(net329),
    .S(_2692_),
    .X(_2169_));
 sky130_fd_sc_hd__o2bb2a_1 _5457_ (.A1_N(_1396_),
    .A2_N(_2161_),
    .B1(_2169_),
    .B2(net160),
    .X(_2170_));
 sky130_fd_sc_hd__o211ai_1 _5458_ (.A1(net77),
    .A2(_2168_),
    .B1(_2170_),
    .C1(net89),
    .Y(_2171_));
 sky130_fd_sc_hd__o31a_1 _5459_ (.A1(_2008_),
    .A2(_2159_),
    .A3(_2160_),
    .B1(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__a21bo_1 _5460_ (.A1(net155),
    .A2(_2166_),
    .B1_N(_1947_),
    .X(_2173_));
 sky130_fd_sc_hd__o221a_1 _5461_ (.A1(net99),
    .A2(_2172_),
    .B1(_2173_),
    .B2(_2167_),
    .C1(net144),
    .X(_2174_));
 sky130_fd_sc_hd__o21a_1 _5462_ (.A1(_2029_),
    .A2(_2161_),
    .B1(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__nand2_1 _5463_ (.A(net64),
    .B(_2168_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_1 _5464_ (.A(_2827_),
    .B(_2161_),
    .X(_2177_));
 sky130_fd_sc_hd__a31o_1 _5465_ (.A1(net72),
    .A2(_2176_),
    .A3(_2177_),
    .B1(_2175_),
    .X(_2178_));
 sky130_fd_sc_hd__o22a_1 _5466_ (.A1(\as2650.stack[7][7] ),
    .A2(net193),
    .B1(net190),
    .B2(\as2650.stack[6][7] ),
    .X(_2179_));
 sky130_fd_sc_hd__o221a_1 _5467_ (.A1(\as2650.stack[4][7] ),
    .A2(net170),
    .B1(net166),
    .B2(\as2650.stack[5][7] ),
    .C1(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__o22a_1 _5468_ (.A1(\as2650.stack[0][7] ),
    .A2(net168),
    .B1(net164),
    .B2(\as2650.stack[1][7] ),
    .X(_2181_));
 sky130_fd_sc_hd__o221a_1 _5469_ (.A1(\as2650.stack[3][7] ),
    .A2(net193),
    .B1(net189),
    .B2(\as2650.stack[2][7] ),
    .C1(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_4 _5470_ (.A0(_2180_),
    .A1(_2182_),
    .S(_2859_),
    .X(_2183_));
 sky130_fd_sc_hd__o2bb2a_1 _5471_ (.A1_N(_0830_),
    .A2_N(_2183_),
    .B1(_2161_),
    .B2(net104),
    .X(_2184_));
 sky130_fd_sc_hd__a21o_1 _5472_ (.A1(_2178_),
    .A2(_2184_),
    .B1(net65),
    .X(_2185_));
 sky130_fd_sc_hd__o211ai_1 _5473_ (.A1(net68),
    .A2(_2161_),
    .B1(_2185_),
    .C1(net45),
    .Y(_2186_));
 sky130_fd_sc_hd__o211a_1 _5474_ (.A1(net275),
    .A2(net45),
    .B1(_2186_),
    .C1(net319),
    .X(_0223_));
 sky130_fd_sc_hd__o21a_2 _5475_ (.A1(_2164_),
    .A2(_2165_),
    .B1(_2162_),
    .X(_2187_));
 sky130_fd_sc_hd__nor2_2 _5476_ (.A(net152),
    .B(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__a21oi_1 _5477_ (.A1(net310),
    .A2(_2188_),
    .B1(_2681_),
    .Y(_2189_));
 sky130_fd_sc_hd__o21ai_1 _5478_ (.A1(net310),
    .A2(_2188_),
    .B1(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__mux2_2 _5479_ (.A0(_2631_),
    .A1(_1681_),
    .S(net311),
    .X(_2191_));
 sky130_fd_sc_hd__and3_2 _5480_ (.A(net274),
    .B(net276),
    .C(_2133_),
    .X(_2192_));
 sky130_fd_sc_hd__a21oi_2 _5481_ (.A1(net276),
    .A2(_2133_),
    .B1(\as2650.pc[8] ),
    .Y(_2193_));
 sky130_fd_sc_hd__nor2_4 _5482_ (.A(_2192_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(net349),
    .A1(\as2650.addr_buff[0] ),
    .S(net148),
    .X(_2195_));
 sky130_fd_sc_hd__o221a_1 _5484_ (.A1(net63),
    .A2(_2194_),
    .B1(_2195_),
    .B2(net160),
    .C1(net97),
    .X(_2196_));
 sky130_fd_sc_hd__a21bo_1 _5485_ (.A1(_2741_),
    .A2(_2191_),
    .B1_N(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__a21oi_1 _5486_ (.A1(_2190_),
    .A2(_2197_),
    .B1(net92),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(\as2650.pc[8] ),
    .B(_2159_),
    .Y(_2199_));
 sky130_fd_sc_hd__or2_1 _5488_ (.A(net274),
    .B(_2159_),
    .X(_2200_));
 sky130_fd_sc_hd__a31o_1 _5489_ (.A1(_2009_),
    .A2(_2199_),
    .A3(_2200_),
    .B1(net72),
    .X(_2201_));
 sky130_fd_sc_hd__a211o_1 _5490_ (.A1(_2028_),
    .A2(_2194_),
    .B1(_2198_),
    .C1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__nor2_1 _5491_ (.A(net92),
    .B(_2191_),
    .Y(_2203_));
 sky130_fd_sc_hd__a211o_1 _5492_ (.A1(net92),
    .A2(_2194_),
    .B1(_2203_),
    .C1(net144),
    .X(_2204_));
 sky130_fd_sc_hd__o22a_1 _5493_ (.A1(_2863_),
    .A2(net102),
    .B1(_2194_),
    .B2(net104),
    .X(_2205_));
 sky130_fd_sc_hd__and3_1 _5494_ (.A(net69),
    .B(_2204_),
    .C(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__a221o_1 _5495_ (.A1(net65),
    .A2(_2194_),
    .B1(_2202_),
    .B2(_2206_),
    .C1(_1971_),
    .X(_2207_));
 sky130_fd_sc_hd__o211a_1 _5496_ (.A1(net274),
    .A2(net46),
    .B1(_2207_),
    .C1(net315),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_2 _5497_ (.A0(net273),
    .A1(_1711_),
    .S(net311),
    .X(_2208_));
 sky130_fd_sc_hd__nor2_1 _5498_ (.A(net77),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__and2_4 _5499_ (.A(net273),
    .B(_2192_),
    .X(_2210_));
 sky130_fd_sc_hd__nor2_1 _5500_ (.A(\as2650.pc[9] ),
    .B(_2192_),
    .Y(_2211_));
 sky130_fd_sc_hd__or2_4 _5501_ (.A(_2210_),
    .B(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__a32o_1 _5502_ (.A1(net159),
    .A2(_1707_),
    .A3(_1980_),
    .B1(_2212_),
    .B2(_1396_),
    .X(_2213_));
 sky130_fd_sc_hd__or3_1 _5503_ (.A(net139),
    .B(_2209_),
    .C(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__and3_2 _5504_ (.A(net273),
    .B(\as2650.pc[8] ),
    .C(_2159_),
    .X(_2215_));
 sky130_fd_sc_hd__a21oi_1 _5505_ (.A1(\as2650.pc[8] ),
    .A2(_2159_),
    .B1(net273),
    .Y(_2216_));
 sky130_fd_sc_hd__o31a_1 _5506_ (.A1(_2008_),
    .A2(_2215_),
    .A3(_2216_),
    .B1(_2214_),
    .X(_2217_));
 sky130_fd_sc_hd__or2_1 _5507_ (.A(net99),
    .B(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__a21oi_1 _5508_ (.A1(\as2650.addr_buff[0] ),
    .A2(_2188_),
    .B1(\as2650.addr_buff[1] ),
    .Y(_2219_));
 sky130_fd_sc_hd__and3b_1 _5509_ (.A_N(_2187_),
    .B(_1689_),
    .C(net153),
    .X(_2220_));
 sky130_fd_sc_hd__or3b_2 _5510_ (.A(_2219_),
    .B(_2220_),
    .C_N(_1947_),
    .X(_2221_));
 sky130_fd_sc_hd__o211a_1 _5511_ (.A1(_2029_),
    .A2(_2212_),
    .B1(_2218_),
    .C1(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__nor2_1 _5512_ (.A(net93),
    .B(_2208_),
    .Y(_2223_));
 sky130_fd_sc_hd__nor2_1 _5513_ (.A(net68),
    .B(_2212_),
    .Y(_2224_));
 sky130_fd_sc_hd__a211o_1 _5514_ (.A1(net139),
    .A2(_2212_),
    .B1(_2223_),
    .C1(net145),
    .X(_2225_));
 sky130_fd_sc_hd__o221a_1 _5515_ (.A1(_2942_),
    .A2(net102),
    .B1(_2212_),
    .B2(net104),
    .C1(_2225_),
    .X(_2226_));
 sky130_fd_sc_hd__o21ai_1 _5516_ (.A1(net72),
    .A2(_2222_),
    .B1(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a21o_1 _5517_ (.A1(net67),
    .A2(_2227_),
    .B1(_1971_),
    .X(_2228_));
 sky130_fd_sc_hd__o221a_1 _5518_ (.A1(\as2650.pc[9] ),
    .A2(net45),
    .B1(_2224_),
    .B2(_2228_),
    .C1(net319),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_1 _5519_ (.A(\as2650.addr_buff[2] ),
    .B(_2220_),
    .Y(_2229_));
 sky130_fd_sc_hd__a21o_1 _5520_ (.A1(_1719_),
    .A2(_2188_),
    .B1(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(_2630_),
    .A1(_1734_),
    .S(net311),
    .X(_2231_));
 sky130_fd_sc_hd__xnor2_4 _5522_ (.A(net272),
    .B(_2210_),
    .Y(_2232_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(net342),
    .A1(\as2650.addr_buff[2] ),
    .S(net148),
    .X(_2233_));
 sky130_fd_sc_hd__a21oi_1 _5524_ (.A1(net157),
    .A2(_2233_),
    .B1(net100),
    .Y(_2234_));
 sky130_fd_sc_hd__o221a_1 _5525_ (.A1(net77),
    .A2(_2231_),
    .B1(_2232_),
    .B2(net63),
    .C1(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__a21o_1 _5526_ (.A1(_2680_),
    .A2(_2230_),
    .B1(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__xnor2_1 _5527_ (.A(net271),
    .B(_2215_),
    .Y(_2237_));
 sky130_fd_sc_hd__a22o_1 _5528_ (.A1(net132),
    .A2(_2236_),
    .B1(_2237_),
    .B2(_2009_),
    .X(_2238_));
 sky130_fd_sc_hd__a211o_1 _5529_ (.A1(_2028_),
    .A2(_2232_),
    .B1(_2238_),
    .C1(net146),
    .X(_2239_));
 sky130_fd_sc_hd__a221o_1 _5530_ (.A1(net64),
    .A2(_2231_),
    .B1(_2232_),
    .B2(_2826_),
    .C1(_0579_),
    .X(_2240_));
 sky130_fd_sc_hd__nand2_1 _5531_ (.A(_2239_),
    .B(_2240_),
    .Y(_2241_));
 sky130_fd_sc_hd__o2bb2a_1 _5532_ (.A1_N(_0814_),
    .A2_N(_2232_),
    .B1(net102),
    .B2(_2993_),
    .X(_2242_));
 sky130_fd_sc_hd__o21ai_1 _5533_ (.A1(net67),
    .A2(_2232_),
    .B1(net45),
    .Y(_2243_));
 sky130_fd_sc_hd__a31o_1 _5534_ (.A1(net67),
    .A2(_2241_),
    .A3(_2242_),
    .B1(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__o211a_1 _5535_ (.A1(net272),
    .A2(net45),
    .B1(_2244_),
    .C1(net319),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_1 _5536_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2220_),
    .B1(\as2650.addr_buff[3] ),
    .Y(_2245_));
 sky130_fd_sc_hd__and2_1 _5537_ (.A(_1768_),
    .B(_2220_),
    .X(_2246_));
 sky130_fd_sc_hd__o21ai_1 _5538_ (.A1(_2245_),
    .A2(_2246_),
    .B1(_2680_),
    .Y(_2247_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(net270),
    .A1(_1759_),
    .S(net311),
    .X(_2248_));
 sky130_fd_sc_hd__and3_1 _5540_ (.A(\as2650.pc[11] ),
    .B(net272),
    .C(_2210_),
    .X(_2249_));
 sky130_fd_sc_hd__a21oi_1 _5541_ (.A1(net272),
    .A2(_2210_),
    .B1(net270),
    .Y(_2250_));
 sky130_fd_sc_hd__or2_4 _5542_ (.A(_2249_),
    .B(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net341),
    .A1(\as2650.addr_buff[3] ),
    .S(net148),
    .X(_2252_));
 sky130_fd_sc_hd__a2bb2o_1 _5544_ (.A1_N(net63),
    .A2_N(_2251_),
    .B1(_2252_),
    .B2(net157),
    .X(_2253_));
 sky130_fd_sc_hd__a211o_1 _5545_ (.A1(_2741_),
    .A2(_2248_),
    .B1(_2253_),
    .C1(net100),
    .X(_2254_));
 sky130_fd_sc_hd__a21oi_1 _5546_ (.A1(_2247_),
    .A2(_2254_),
    .B1(net92),
    .Y(_2255_));
 sky130_fd_sc_hd__and3_1 _5547_ (.A(net270),
    .B(net271),
    .C(_2215_),
    .X(_2256_));
 sky130_fd_sc_hd__a21oi_1 _5548_ (.A1(net272),
    .A2(_2215_),
    .B1(net270),
    .Y(_2257_));
 sky130_fd_sc_hd__o21a_1 _5549_ (.A1(_2256_),
    .A2(_2257_),
    .B1(_2009_),
    .X(_2258_));
 sky130_fd_sc_hd__a2111o_1 _5550_ (.A1(_2028_),
    .A2(_2251_),
    .B1(_2255_),
    .C1(_2258_),
    .D1(net72),
    .X(_2259_));
 sky130_fd_sc_hd__nor2_1 _5551_ (.A(net92),
    .B(_2248_),
    .Y(_2260_));
 sky130_fd_sc_hd__a211o_1 _5552_ (.A1(net92),
    .A2(_2251_),
    .B1(_2260_),
    .C1(net144),
    .X(_2261_));
 sky130_fd_sc_hd__o221a_1 _5553_ (.A1(_0340_),
    .A2(net102),
    .B1(_2251_),
    .B2(net104),
    .C1(_2259_),
    .X(_2262_));
 sky130_fd_sc_hd__a21oi_1 _5554_ (.A1(_2261_),
    .A2(_2262_),
    .B1(net65),
    .Y(_2263_));
 sky130_fd_sc_hd__o21ai_1 _5555_ (.A1(net69),
    .A2(_2251_),
    .B1(net46),
    .Y(_2264_));
 sky130_fd_sc_hd__o221a_1 _5556_ (.A1(net270),
    .A2(net46),
    .B1(_2263_),
    .B2(_2264_),
    .C1(net315),
    .X(_0227_));
 sky130_fd_sc_hd__and2_2 _5557_ (.A(net269),
    .B(_2249_),
    .X(_2265_));
 sky130_fd_sc_hd__nor2_1 _5558_ (.A(\as2650.pc[12] ),
    .B(_2249_),
    .Y(_2266_));
 sky130_fd_sc_hd__nor2_2 _5559_ (.A(_2265_),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__xnor2_1 _5560_ (.A(\as2650.addr_buff[4] ),
    .B(_2246_),
    .Y(_2268_));
 sky130_fd_sc_hd__mux2_2 _5561_ (.A0(net269),
    .A1(_1783_),
    .S(net312),
    .X(_2269_));
 sky130_fd_sc_hd__o21ai_1 _5562_ (.A1(_2662_),
    .A2(net147),
    .B1(_2080_),
    .Y(_2270_));
 sky130_fd_sc_hd__a221o_1 _5563_ (.A1(_1396_),
    .A2(_2267_),
    .B1(_2270_),
    .B2(net157),
    .C1(net99),
    .X(_2271_));
 sky130_fd_sc_hd__a21oi_1 _5564_ (.A1(_2741_),
    .A2(_2269_),
    .B1(_2271_),
    .Y(_2272_));
 sky130_fd_sc_hd__a21oi_1 _5565_ (.A1(_2680_),
    .A2(_2268_),
    .B1(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__and2_1 _5566_ (.A(net269),
    .B(_2256_),
    .X(_2274_));
 sky130_fd_sc_hd__nor2_1 _5567_ (.A(net269),
    .B(_2256_),
    .Y(_2275_));
 sky130_fd_sc_hd__o21ai_1 _5568_ (.A1(_2274_),
    .A2(_2275_),
    .B1(_2009_),
    .Y(_2276_));
 sky130_fd_sc_hd__o211a_1 _5569_ (.A1(net137),
    .A2(_2273_),
    .B1(_2276_),
    .C1(_0579_),
    .X(_2277_));
 sky130_fd_sc_hd__or2_1 _5570_ (.A(net89),
    .B(_2267_),
    .X(_2278_));
 sky130_fd_sc_hd__o211a_1 _5571_ (.A1(net92),
    .A2(_2269_),
    .B1(_2278_),
    .C1(net146),
    .X(_2279_));
 sky130_fd_sc_hd__or2_1 _5572_ (.A(net67),
    .B(_2267_),
    .X(_2280_));
 sky130_fd_sc_hd__o32a_1 _5573_ (.A1(net66),
    .A2(_2277_),
    .A3(_2279_),
    .B1(_2029_),
    .B2(_2267_),
    .X(_2281_));
 sky130_fd_sc_hd__a21o_1 _5574_ (.A1(_0392_),
    .A2(_0830_),
    .B1(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__a221o_1 _5575_ (.A1(_0814_),
    .A2(_2267_),
    .B1(_2280_),
    .B2(_2282_),
    .C1(_1971_),
    .X(_2283_));
 sky130_fd_sc_hd__o211a_1 _5576_ (.A1(net269),
    .A2(_1970_),
    .B1(_2283_),
    .C1(net319),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_4 _5577_ (.A(\as2650.pc[13] ),
    .B(_2265_),
    .Y(_2284_));
 sky130_fd_sc_hd__or2_1 _5578_ (.A(\as2650.pc[13] ),
    .B(_2265_),
    .X(_2285_));
 sky130_fd_sc_hd__nand2_2 _5579_ (.A(_2284_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__a22o_1 _5581_ (.A1(_0443_),
    .A2(_0830_),
    .B1(_2287_),
    .B2(_0814_),
    .X(_2288_));
 sky130_fd_sc_hd__or2_1 _5582_ (.A(\as2650.pc[13] ),
    .B(_2274_),
    .X(_2289_));
 sky130_fd_sc_hd__nand2_1 _5583_ (.A(\as2650.pc[13] ),
    .B(_2274_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(_1861_),
    .B(_2286_),
    .Y(_2291_));
 sky130_fd_sc_hd__a31o_1 _5585_ (.A1(_1861_),
    .A2(_2289_),
    .A3(_2290_),
    .B1(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__a221o_1 _5586_ (.A1(\as2650.addr_buff[5] ),
    .A2(net155),
    .B1(_1396_),
    .B2(_2287_),
    .C1(_2676_),
    .X(_2293_));
 sky130_fd_sc_hd__a21o_1 _5587_ (.A1(net93),
    .A2(_2292_),
    .B1(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__a31o_1 _5588_ (.A1(\as2650.pc[13] ),
    .A2(net329),
    .A3(_2741_),
    .B1(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__a31o_1 _5589_ (.A1(net93),
    .A2(_2284_),
    .A3(_2285_),
    .B1(net144),
    .X(_2296_));
 sky130_fd_sc_hd__nor2_1 _5590_ (.A(net141),
    .B(_2286_),
    .Y(_2297_));
 sky130_fd_sc_hd__a32o_1 _5591_ (.A1(\as2650.pc[13] ),
    .A2(net329),
    .A3(_1393_),
    .B1(_2296_),
    .B2(net237),
    .X(_2298_));
 sky130_fd_sc_hd__a22o_1 _5592_ (.A1(\as2650.addr_buff[5] ),
    .A2(net147),
    .B1(_2246_),
    .B2(\as2650.addr_buff[4] ),
    .X(_2299_));
 sky130_fd_sc_hd__a211o_1 _5593_ (.A1(net141),
    .A2(_2299_),
    .B1(_2297_),
    .C1(net97),
    .X(_2300_));
 sky130_fd_sc_hd__a31o_1 _5594_ (.A1(_2295_),
    .A2(_2298_),
    .A3(_2300_),
    .B1(_2288_),
    .X(_2301_));
 sky130_fd_sc_hd__nor2_1 _5595_ (.A(net67),
    .B(_2286_),
    .Y(_2302_));
 sky130_fd_sc_hd__a21o_1 _5596_ (.A1(net67),
    .A2(_2301_),
    .B1(_1971_),
    .X(_2303_));
 sky130_fd_sc_hd__o221a_1 _5597_ (.A1(\as2650.pc[13] ),
    .A2(_1970_),
    .B1(_2302_),
    .B2(_2303_),
    .C1(net319),
    .X(_0229_));
 sky130_fd_sc_hd__xnor2_4 _5598_ (.A(\as2650.pc[14] ),
    .B(_2284_),
    .Y(_2304_));
 sky130_fd_sc_hd__and2_1 _5599_ (.A(\as2650.pc[14] ),
    .B(net330),
    .X(_2305_));
 sky130_fd_sc_hd__o221a_1 _5600_ (.A1(\as2650.addr_buff[6] ),
    .A2(net160),
    .B1(_2742_),
    .B2(_2305_),
    .C1(_2694_),
    .X(_2306_));
 sky130_fd_sc_hd__o21a_1 _5601_ (.A1(net63),
    .A2(_2304_),
    .B1(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__xnor2_1 _5602_ (.A(\as2650.pc[14] ),
    .B(_2290_),
    .Y(_2308_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(_2304_),
    .A1(_2308_),
    .S(_1861_),
    .X(_2309_));
 sky130_fd_sc_hd__a211o_1 _5604_ (.A1(net137),
    .A2(_2309_),
    .B1(_2307_),
    .C1(net100),
    .X(_2310_));
 sky130_fd_sc_hd__and3_1 _5605_ (.A(\as2650.addr_buff[6] ),
    .B(_2693_),
    .C(net141),
    .X(_2311_));
 sky130_fd_sc_hd__a211o_1 _5606_ (.A1(net143),
    .A2(_2304_),
    .B1(_2311_),
    .C1(net97),
    .X(_2312_));
 sky130_fd_sc_hd__a21o_1 _5607_ (.A1(_2310_),
    .A2(_2312_),
    .B1(net72),
    .X(_2313_));
 sky130_fd_sc_hd__a31o_1 _5608_ (.A1(\as2650.pc[14] ),
    .A2(net330),
    .A3(net135),
    .B1(net144),
    .X(_2314_));
 sky130_fd_sc_hd__a21o_1 _5609_ (.A1(net94),
    .A2(_2304_),
    .B1(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__o221a_1 _5610_ (.A1(_0496_),
    .A2(net102),
    .B1(_2304_),
    .B2(net104),
    .C1(net68),
    .X(_2316_));
 sky130_fd_sc_hd__and2_1 _5611_ (.A(_2315_),
    .B(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__a221o_1 _5612_ (.A1(net66),
    .A2(_2304_),
    .B1(_2313_),
    .B2(_2317_),
    .C1(_1971_),
    .X(_2318_));
 sky130_fd_sc_hd__o211a_1 _5613_ (.A1(\as2650.pc[14] ),
    .A2(_1970_),
    .B1(_2318_),
    .C1(net319),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _5614_ (.A(net150),
    .B(_2934_),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _5615_ (.A0(_2906_),
    .A1(_2912_),
    .S(net83),
    .X(_2320_));
 sky130_fd_sc_hd__o211a_1 _5616_ (.A1(net155),
    .A2(_2320_),
    .B1(_2319_),
    .C1(net81),
    .X(_2321_));
 sky130_fd_sc_hd__or3_1 _5617_ (.A(_2783_),
    .B(net197),
    .C(_0834_),
    .X(_2322_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(net204),
    .A2(_2782_),
    .B1(_2799_),
    .B2(_2692_),
    .X(_2323_));
 sky130_fd_sc_hd__o211a_1 _5619_ (.A1(net204),
    .A2(_2780_),
    .B1(_2648_),
    .C1(net85),
    .X(_2324_));
 sky130_fd_sc_hd__o21ai_1 _5620_ (.A1(_2323_),
    .A2(_2324_),
    .B1(net214),
    .Y(_2325_));
 sky130_fd_sc_hd__o21ai_1 _5621_ (.A1(_2815_),
    .A2(net71),
    .B1(_2796_),
    .Y(_2326_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(net204),
    .B(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__a31o_1 _5623_ (.A1(net298),
    .A2(net94),
    .A3(net205),
    .B1(_0580_),
    .X(_2328_));
 sky130_fd_sc_hd__a21o_1 _5624_ (.A1(_0587_),
    .A2(_2328_),
    .B1(_2646_),
    .X(_2329_));
 sky130_fd_sc_hd__or3_2 _5625_ (.A(net232),
    .B(_2698_),
    .C(_1347_),
    .X(_2330_));
 sky130_fd_sc_hd__nor2_1 _5626_ (.A(net127),
    .B(_2900_),
    .Y(_2331_));
 sky130_fd_sc_hd__and2_1 _5627_ (.A(\as2650.carry ),
    .B(_0759_),
    .X(_2332_));
 sky130_fd_sc_hd__a211o_1 _5628_ (.A1(\as2650.psu[0] ),
    .A2(_0758_),
    .B1(_2332_),
    .C1(_2813_),
    .X(_2333_));
 sky130_fd_sc_hd__o221a_1 _5629_ (.A1(net124),
    .A2(_0605_),
    .B1(_1956_),
    .B2(net73),
    .C1(net71),
    .X(_2334_));
 sky130_fd_sc_hd__a221o_1 _5630_ (.A1(_2758_),
    .A2(net120),
    .B1(_2333_),
    .B2(_2334_),
    .C1(net126),
    .X(_2335_));
 sky130_fd_sc_hd__o221a_1 _5631_ (.A1(net348),
    .A2(_2792_),
    .B1(_2331_),
    .B2(_2335_),
    .C1(net171),
    .X(_2336_));
 sky130_fd_sc_hd__and4_1 _5632_ (.A(_0839_),
    .B(_2325_),
    .C(_2327_),
    .D(_2329_),
    .X(_2337_));
 sky130_fd_sc_hd__a31o_2 _5633_ (.A1(\as2650.cycle[7] ),
    .A2(net213),
    .A3(net131),
    .B1(net294),
    .X(_2338_));
 sky130_fd_sc_hd__or4_1 _5634_ (.A(net231),
    .B(_0807_),
    .C(_0823_),
    .D(_0827_),
    .X(_2339_));
 sky130_fd_sc_hd__nor2_1 _5635_ (.A(net198),
    .B(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__or3b_1 _5636_ (.A(_2338_),
    .B(_2340_),
    .C_N(_1342_),
    .X(_2341_));
 sky130_fd_sc_hd__or3b_1 _5637_ (.A(_2341_),
    .B(_0819_),
    .C_N(_2337_),
    .X(_2342_));
 sky130_fd_sc_hd__and3_1 _5638_ (.A(_2677_),
    .B(net103),
    .C(_1796_),
    .X(_2343_));
 sky130_fd_sc_hd__and3_1 _5639_ (.A(_2740_),
    .B(_1793_),
    .C(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__and4b_1 _5640_ (.A_N(_2735_),
    .B(_0829_),
    .C(_1369_),
    .D(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__o2111a_1 _5641_ (.A1(net80),
    .A2(_2801_),
    .B1(_2322_),
    .C1(_2330_),
    .D1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__or3b_4 _5642_ (.A(_0828_),
    .B(_2342_),
    .C_N(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__o2111a_1 _5643_ (.A1(_2724_),
    .A2(_2801_),
    .B1(_2322_),
    .C1(_2329_),
    .D1(_2330_),
    .X(_2348_));
 sky130_fd_sc_hd__and3_1 _5644_ (.A(_0839_),
    .B(_2325_),
    .C(_2327_),
    .X(_2349_));
 sky130_fd_sc_hd__nor2_1 _5645_ (.A(_0828_),
    .B(_2341_),
    .Y(_2350_));
 sky130_fd_sc_hd__o31a_1 _5646_ (.A1(net236),
    .A2(net133),
    .A3(_2865_),
    .B1(_0821_),
    .X(_2351_));
 sky130_fd_sc_hd__and4b_1 _5647_ (.A_N(_2735_),
    .B(_2740_),
    .C(_0844_),
    .D(_2343_),
    .X(_2352_));
 sky130_fd_sc_hd__and4b_1 _5648_ (.A_N(_1791_),
    .B(_2350_),
    .C(_2351_),
    .D(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__and3_4 _5649_ (.A(_2348_),
    .B(_2349_),
    .C(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__a2111o_1 _5650_ (.A1(net121),
    .A2(net59),
    .B1(_2321_),
    .C1(_2336_),
    .D1(_2347_),
    .X(_2355_));
 sky130_fd_sc_hd__o21ba_1 _5651_ (.A1(net211),
    .A2(_2881_),
    .B1_N(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__a211oi_1 _5652_ (.A1(_2629_),
    .A2(_2347_),
    .B1(_2356_),
    .C1(net325),
    .Y(_0231_));
 sky130_fd_sc_hd__or2_1 _5653_ (.A(net150),
    .B(_2986_),
    .X(_2357_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(_2962_),
    .A1(_2965_),
    .S(net83),
    .X(_2358_));
 sky130_fd_sc_hd__o211a_1 _5655_ (.A1(net155),
    .A2(_2358_),
    .B1(_2357_),
    .C1(net82),
    .X(_2359_));
 sky130_fd_sc_hd__nor2_1 _5656_ (.A(_2623_),
    .B(_0773_),
    .Y(_2360_));
 sky130_fd_sc_hd__a21o_1 _5657_ (.A1(net226),
    .A2(_0758_),
    .B1(_2813_),
    .X(_2361_));
 sky130_fd_sc_hd__o21a_1 _5658_ (.A1(net124),
    .A2(_0608_),
    .B1(net71),
    .X(_2362_));
 sky130_fd_sc_hd__o221a_1 _5659_ (.A1(net73),
    .A2(_2001_),
    .B1(_2360_),
    .B2(_2361_),
    .C1(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__a221o_1 _5660_ (.A1(_2773_),
    .A2(net121),
    .B1(net116),
    .B2(_2758_),
    .C1(net126),
    .X(_2364_));
 sky130_fd_sc_hd__o221a_1 _5661_ (.A1(net2),
    .A2(_2792_),
    .B1(_2363_),
    .B2(_2364_),
    .C1(net171),
    .X(_2365_));
 sky130_fd_sc_hd__a211o_1 _5662_ (.A1(net120),
    .A2(net59),
    .B1(_2347_),
    .C1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__a211o_1 _5663_ (.A1(net173),
    .A2(_2947_),
    .B1(_2359_),
    .C1(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__o211a_1 _5664_ (.A1(net263),
    .A2(_2354_),
    .B1(_2367_),
    .C1(net320),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(_0312_),
    .A1(_0316_),
    .S(net83),
    .X(_2368_));
 sky130_fd_sc_hd__o21a_1 _5666_ (.A1(net156),
    .A2(_2368_),
    .B1(net82),
    .X(_2369_));
 sky130_fd_sc_hd__o21a_1 _5667_ (.A1(net151),
    .A2(_0333_),
    .B1(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__nor2_1 _5668_ (.A(_2625_),
    .B(_0773_),
    .Y(_2371_));
 sky130_fd_sc_hd__a21o_1 _5669_ (.A1(\as2650.psu[2] ),
    .A2(_0758_),
    .B1(_2813_),
    .X(_2372_));
 sky130_fd_sc_hd__o21a_1 _5670_ (.A1(net124),
    .A2(net187),
    .B1(net71),
    .X(_2373_));
 sky130_fd_sc_hd__o221a_1 _5671_ (.A1(net74),
    .A2(_2039_),
    .B1(_2371_),
    .B2(_2372_),
    .C1(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__a221o_1 _5672_ (.A1(_2773_),
    .A2(net120),
    .B1(net112),
    .B2(_2758_),
    .C1(net126),
    .X(_2375_));
 sky130_fd_sc_hd__o221a_1 _5673_ (.A1(net3),
    .A2(_2792_),
    .B1(_2374_),
    .B2(_2375_),
    .C1(net171),
    .X(_2376_));
 sky130_fd_sc_hd__a221o_1 _5674_ (.A1(net173),
    .A2(_0300_),
    .B1(net59),
    .B2(net116),
    .C1(_2347_),
    .X(_2377_));
 sky130_fd_sc_hd__or3_2 _5675_ (.A(_2370_),
    .B(_2376_),
    .C(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__o211a_1 _5676_ (.A1(net259),
    .A2(_2354_),
    .B1(_2378_),
    .C1(net320),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _5677_ (.A(net156),
    .B(_0382_),
    .Y(_2379_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(_0362_),
    .A1(_0364_),
    .S(net83),
    .X(_2380_));
 sky130_fd_sc_hd__o211a_1 _5679_ (.A1(net156),
    .A2(_2380_),
    .B1(_2379_),
    .C1(net82),
    .X(_2381_));
 sky130_fd_sc_hd__a21o_1 _5680_ (.A1(\as2650.psl[3] ),
    .A2(_0759_),
    .B1(_2813_),
    .X(_2382_));
 sky130_fd_sc_hd__a21o_1 _5681_ (.A1(\as2650.psu[3] ),
    .A2(_0758_),
    .B1(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__o221a_1 _5682_ (.A1(net124),
    .A2(net185),
    .B1(_2069_),
    .B2(net73),
    .C1(net71),
    .X(_2384_));
 sky130_fd_sc_hd__a221o_1 _5683_ (.A1(_2773_),
    .A2(net117),
    .B1(_0353_),
    .B2(_2758_),
    .C1(net126),
    .X(_2385_));
 sky130_fd_sc_hd__a21o_1 _5684_ (.A1(_2383_),
    .A2(_2384_),
    .B1(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__o211a_1 _5685_ (.A1(net4),
    .A2(_2792_),
    .B1(net171),
    .C1(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__a221o_1 _5686_ (.A1(net173),
    .A2(_0344_),
    .B1(net59),
    .B2(net112),
    .C1(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__or3_2 _5687_ (.A(_2347_),
    .B(_2381_),
    .C(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__o211a_1 _5688_ (.A1(net255),
    .A2(_2354_),
    .B1(_2389_),
    .C1(net320),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(_0413_),
    .A1(_0416_),
    .S(net83),
    .X(_2390_));
 sky130_fd_sc_hd__or2_1 _5690_ (.A(net156),
    .B(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__o211a_1 _5691_ (.A1(net151),
    .A2(_0434_),
    .B1(_2391_),
    .C1(net82),
    .X(_2392_));
 sky130_fd_sc_hd__nor2_1 _5692_ (.A(\as2650.psu[4] ),
    .B(_0759_),
    .Y(_2393_));
 sky130_fd_sc_hd__a211o_1 _5693_ (.A1(_2624_),
    .A2(_0759_),
    .B1(_2393_),
    .C1(_2807_),
    .X(_2394_));
 sky130_fd_sc_hd__o211a_1 _5694_ (.A1(net74),
    .A2(_2096_),
    .B1(_2394_),
    .C1(net124),
    .X(_2395_));
 sky130_fd_sc_hd__o21ai_1 _5695_ (.A1(net124),
    .A2(net183),
    .B1(net127),
    .Y(_2396_));
 sky130_fd_sc_hd__a2bb2o_1 _5696_ (.A1_N(_2395_),
    .A2_N(_2396_),
    .B1(_2773_),
    .B2(net113),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(net109),
    .A1(_2397_),
    .S(net128),
    .X(_2398_));
 sky130_fd_sc_hd__or2_1 _5698_ (.A(_2791_),
    .B(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__a21oi_1 _5699_ (.A1(_2655_),
    .A2(_2791_),
    .B1(_2794_),
    .Y(_2400_));
 sky130_fd_sc_hd__a221o_1 _5700_ (.A1(_2664_),
    .A2(_0402_),
    .B1(_2399_),
    .B2(_2400_),
    .C1(_2347_),
    .X(_2401_));
 sky130_fd_sc_hd__a211o_1 _5701_ (.A1(_0353_),
    .A2(_0824_),
    .B1(_2392_),
    .C1(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__o211a_1 _5702_ (.A1(net253),
    .A2(_2354_),
    .B1(_2402_),
    .C1(net320),
    .X(_0235_));
 sky130_fd_sc_hd__and2_1 _5703_ (.A(net83),
    .B(_0452_),
    .X(_2403_));
 sky130_fd_sc_hd__a211o_1 _5704_ (.A1(net86),
    .A2(_0469_),
    .B1(_2403_),
    .C1(net156),
    .X(_2404_));
 sky130_fd_sc_hd__o211a_1 _5705_ (.A1(net151),
    .A2(_0489_),
    .B1(_2404_),
    .C1(net82),
    .X(_2405_));
 sky130_fd_sc_hd__nor2_1 _5706_ (.A(net211),
    .B(_0455_),
    .Y(_2406_));
 sky130_fd_sc_hd__nor2_1 _5707_ (.A(net127),
    .B(net110),
    .Y(_2407_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(\as2650.psl[5] ),
    .A1(\as2650.psu[5] ),
    .S(_0773_),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(_2124_),
    .A1(_2408_),
    .S(net73),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(_0396_),
    .A1(_2409_),
    .S(net124),
    .X(_2410_));
 sky130_fd_sc_hd__a21o_1 _5711_ (.A1(net127),
    .A2(_2410_),
    .B1(_2407_),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(net106),
    .A1(_2411_),
    .S(net128),
    .X(_2412_));
 sky130_fd_sc_hd__or2_1 _5713_ (.A(_2791_),
    .B(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_2657_),
    .B(_2791_),
    .Y(_2414_));
 sky130_fd_sc_hd__a311o_1 _5715_ (.A1(net171),
    .A2(_2413_),
    .A3(_2414_),
    .B1(_2347_),
    .C1(_2406_),
    .X(_2415_));
 sky130_fd_sc_hd__a211o_2 _5716_ (.A1(net109),
    .A2(_0824_),
    .B1(_2405_),
    .C1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__o211a_1 _5717_ (.A1(net248),
    .A2(_2354_),
    .B1(_2416_),
    .C1(net321),
    .X(_0236_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(net156),
    .B(_0535_),
    .Y(_2417_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(_0515_),
    .A1(_0518_),
    .S(net84),
    .X(_2418_));
 sky130_fd_sc_hd__o211a_1 _5720_ (.A1(net156),
    .A2(_2418_),
    .B1(_2417_),
    .C1(net82),
    .X(_2419_));
 sky130_fd_sc_hd__nor2_1 _5721_ (.A(net211),
    .B(_0506_),
    .Y(_2420_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(\as2650.psl[6] ),
    .A1(net29),
    .S(_0773_),
    .X(_2421_));
 sky130_fd_sc_hd__o221a_1 _5723_ (.A1(net124),
    .A2(net179),
    .B1(_2155_),
    .B2(net73),
    .C1(net71),
    .X(_2422_));
 sky130_fd_sc_hd__o21ai_1 _5724_ (.A1(_2813_),
    .A2(_2421_),
    .B1(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__o221a_1 _5725_ (.A1(_2759_),
    .A2(_2896_),
    .B1(_0399_),
    .B2(_2774_),
    .C1(_2792_),
    .X(_2424_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(_2423_),
    .B(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__a32o_1 _5727_ (.A1(net171),
    .A2(_0862_),
    .A3(_2425_),
    .B1(net106),
    .B2(_0824_),
    .X(_2426_));
 sky130_fd_sc_hd__or4_2 _5728_ (.A(_2347_),
    .B(_2419_),
    .C(_2420_),
    .D(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__o211a_1 _5729_ (.A1(net245),
    .A2(_2354_),
    .B1(_2427_),
    .C1(net320),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _5730_ (.A(net151),
    .B(_0568_),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(_0550_),
    .A1(_0552_),
    .S(net84),
    .X(_2429_));
 sky130_fd_sc_hd__o211a_1 _5732_ (.A1(net156),
    .A2(_2429_),
    .B1(_2428_),
    .C1(net82),
    .X(_2430_));
 sky130_fd_sc_hd__nor2_1 _5733_ (.A(net211),
    .B(_0540_),
    .Y(_2431_));
 sky130_fd_sc_hd__or2_1 _5734_ (.A(net73),
    .B(_2183_),
    .X(_2432_));
 sky130_fd_sc_hd__mux2_1 _5735_ (.A0(\as2650.psl[7] ),
    .A1(\as2650.psu[7] ),
    .S(_0773_),
    .X(_2433_));
 sky130_fd_sc_hd__o221a_1 _5736_ (.A1(net124),
    .A2(_2893_),
    .B1(_2433_),
    .B2(_2813_),
    .C1(_2432_),
    .X(_2434_));
 sky130_fd_sc_hd__o21ai_1 _5737_ (.A1(_0749_),
    .A2(_2434_),
    .B1(_0867_),
    .Y(_2435_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_0860_),
    .B(_2435_),
    .Y(_2436_));
 sky130_fd_sc_hd__a221o_1 _5739_ (.A1(net118),
    .A2(_0824_),
    .B1(_2436_),
    .B2(_2793_),
    .C1(_2347_),
    .X(_2437_));
 sky130_fd_sc_hd__or3_2 _5740_ (.A(_2430_),
    .B(_2431_),
    .C(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__o211a_1 _5741_ (.A1(net241),
    .A2(_2354_),
    .B1(_2438_),
    .C1(net320),
    .X(_0238_));
 sky130_fd_sc_hd__nor3_4 _5742_ (.A(_2627_),
    .B(net190),
    .C(net56),
    .Y(_2439_));
 sky130_fd_sc_hd__or3_4 _5743_ (.A(net219),
    .B(net191),
    .C(net55),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(net288),
    .A1(\as2650.stack[6][0] ),
    .S(_0600_),
    .X(_2441_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(net265),
    .A1(_2441_),
    .S(_2440_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _5746_ (.A(\as2650.stack[6][1] ),
    .B(_0599_),
    .X(_2442_));
 sky130_fd_sc_hd__o21a_1 _5747_ (.A1(net285),
    .A2(_0600_),
    .B1(_2440_),
    .X(_2443_));
 sky130_fd_sc_hd__a22o_1 _5748_ (.A1(net261),
    .A2(_2439_),
    .B1(_2442_),
    .B2(_2443_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _5749_ (.A(\as2650.stack[6][2] ),
    .B(_0599_),
    .X(_2444_));
 sky130_fd_sc_hd__a21oi_1 _5750_ (.A1(_2634_),
    .A2(_0599_),
    .B1(_2439_),
    .Y(_2445_));
 sky130_fd_sc_hd__a22o_1 _5751_ (.A1(net257),
    .A2(_2439_),
    .B1(_2444_),
    .B2(_2445_),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _5752_ (.A(\as2650.stack[6][3] ),
    .B(_0599_),
    .X(_2446_));
 sky130_fd_sc_hd__a21oi_1 _5753_ (.A1(_2633_),
    .A2(_0599_),
    .B1(_2439_),
    .Y(_2447_));
 sky130_fd_sc_hd__a22o_1 _5754_ (.A1(net254),
    .A2(_2439_),
    .B1(_2446_),
    .B2(_2447_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _5755_ (.A(\as2650.stack[6][4] ),
    .B(_0599_),
    .X(_2448_));
 sky130_fd_sc_hd__a21oi_1 _5756_ (.A1(_2632_),
    .A2(_0599_),
    .B1(_2439_),
    .Y(_2449_));
 sky130_fd_sc_hd__a22o_1 _5757_ (.A1(net251),
    .A2(_2439_),
    .B1(_2448_),
    .B2(_2449_),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _5758_ (.A(\as2650.stack[6][5] ),
    .B(_0599_),
    .X(_2450_));
 sky130_fd_sc_hd__o21a_1 _5759_ (.A1(net280),
    .A2(_0600_),
    .B1(_2440_),
    .X(_2451_));
 sky130_fd_sc_hd__a22o_1 _5760_ (.A1(net247),
    .A2(_2439_),
    .B1(_2450_),
    .B2(_2451_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5761_ (.A0(net277),
    .A1(\as2650.stack[6][6] ),
    .S(_0600_),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(net243),
    .A1(_2452_),
    .S(_2440_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _5763_ (.A(\as2650.stack[6][7] ),
    .B(_0599_),
    .X(_2453_));
 sky130_fd_sc_hd__o21a_1 _5764_ (.A1(net275),
    .A2(_0600_),
    .B1(_2440_),
    .X(_2454_));
 sky130_fd_sc_hd__a22o_1 _5765_ (.A1(net239),
    .A2(_2439_),
    .B1(_2453_),
    .B2(_2454_),
    .X(_0246_));
 sky130_fd_sc_hd__nor3_4 _5766_ (.A(net219),
    .B(net189),
    .C(_0584_),
    .Y(_2455_));
 sky130_fd_sc_hd__or3_4 _5767_ (.A(net219),
    .B(net189),
    .C(net49),
    .X(_2456_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net288),
    .A1(\as2650.stack[7][0] ),
    .S(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_1 _5769_ (.A0(net265),
    .A1(_2457_),
    .S(_1080_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _5770_ (.A(\as2650.stack[7][1] ),
    .B(_2455_),
    .X(_2458_));
 sky130_fd_sc_hd__o21a_1 _5771_ (.A1(net285),
    .A2(_2456_),
    .B1(_1080_),
    .X(_2459_));
 sky130_fd_sc_hd__a22o_1 _5772_ (.A1(net261),
    .A2(_1079_),
    .B1(_2458_),
    .B2(_2459_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _5773_ (.A(\as2650.stack[7][2] ),
    .B(_2455_),
    .X(_2460_));
 sky130_fd_sc_hd__a21oi_1 _5774_ (.A1(_2634_),
    .A2(_2455_),
    .B1(_1079_),
    .Y(_2461_));
 sky130_fd_sc_hd__a22o_1 _5775_ (.A1(net257),
    .A2(_1079_),
    .B1(_2460_),
    .B2(_2461_),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _5776_ (.A(\as2650.stack[7][3] ),
    .B(_2455_),
    .X(_2462_));
 sky130_fd_sc_hd__a21oi_1 _5777_ (.A1(_2633_),
    .A2(_2455_),
    .B1(_1079_),
    .Y(_2463_));
 sky130_fd_sc_hd__a22o_1 _5778_ (.A1(net254),
    .A2(_1079_),
    .B1(_2462_),
    .B2(_2463_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _5779_ (.A(\as2650.stack[7][4] ),
    .B(_2455_),
    .X(_2464_));
 sky130_fd_sc_hd__a21oi_1 _5780_ (.A1(_2632_),
    .A2(_2455_),
    .B1(_1079_),
    .Y(_2465_));
 sky130_fd_sc_hd__a22o_1 _5781_ (.A1(net251),
    .A2(_1079_),
    .B1(_2464_),
    .B2(_2465_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _5782_ (.A(\as2650.stack[7][5] ),
    .B(_2455_),
    .X(_2466_));
 sky130_fd_sc_hd__o21a_1 _5783_ (.A1(net280),
    .A2(_2456_),
    .B1(_1080_),
    .X(_2467_));
 sky130_fd_sc_hd__a22o_1 _5784_ (.A1(net247),
    .A2(_1079_),
    .B1(_2466_),
    .B2(_2467_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _5785_ (.A(\as2650.stack[7][6] ),
    .B(_2455_),
    .X(_2468_));
 sky130_fd_sc_hd__o21a_1 _5786_ (.A1(net277),
    .A2(_2456_),
    .B1(_1080_),
    .X(_2469_));
 sky130_fd_sc_hd__a22o_1 _5787_ (.A1(net243),
    .A2(_1079_),
    .B1(_2468_),
    .B2(_2469_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _5788_ (.A(\as2650.stack[7][7] ),
    .B(_2455_),
    .X(_2470_));
 sky130_fd_sc_hd__o21a_1 _5789_ (.A1(net276),
    .A2(_2456_),
    .B1(_1080_),
    .X(_2471_));
 sky130_fd_sc_hd__a22o_1 _5790_ (.A1(net239),
    .A2(_1079_),
    .B1(_2470_),
    .B2(_2471_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_8 _5791_ (.A(_2440_),
    .B(_2456_),
    .Y(_2472_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(\as2650.stack[7][8] ),
    .A1(_0607_),
    .S(_2472_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(\as2650.stack[7][9] ),
    .A1(_0610_),
    .S(_2472_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5794_ (.A0(\as2650.stack[7][10] ),
    .A1(_0612_),
    .S(_2472_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(\as2650.stack[7][11] ),
    .A1(_0614_),
    .S(_2472_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(\as2650.stack[7][12] ),
    .A1(_0616_),
    .S(_2472_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(\as2650.stack[7][13] ),
    .A1(_0618_),
    .S(_2472_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5798_ (.A0(\as2650.stack[7][14] ),
    .A1(_0620_),
    .S(_2472_),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_4 _5799_ (.A(net321),
    .B(_2867_),
    .Y(_2473_));
 sky130_fd_sc_hd__nor2_8 _5800_ (.A(net308),
    .B(_2831_),
    .Y(_2474_));
 sky130_fd_sc_hd__nor2_4 _5801_ (.A(_2473_),
    .B(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__a32o_1 _5802_ (.A1(net266),
    .A2(net62),
    .A3(net176),
    .B1(_2474_),
    .B2(_2935_),
    .X(_2476_));
 sky130_fd_sc_hd__a21o_1 _5803_ (.A1(\as2650.r123[1][0] ),
    .A2(_2475_),
    .B1(_2476_),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _5804_ (.A1(_2987_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][1] ),
    .X(_2477_));
 sky130_fd_sc_hd__a21o_1 _5805_ (.A1(net62),
    .A2(_0921_),
    .B1(_2477_),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _5806_ (.A1(_0334_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][2] ),
    .X(_2478_));
 sky130_fd_sc_hd__a21o_1 _5807_ (.A1(net61),
    .A2(_0932_),
    .B1(_2478_),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _5808_ (.A1(_0386_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][3] ),
    .X(_2479_));
 sky130_fd_sc_hd__a21o_1 _5809_ (.A1(net61),
    .A2(_0944_),
    .B1(_2479_),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _5810_ (.A1(_0437_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][4] ),
    .X(_2480_));
 sky130_fd_sc_hd__a21o_1 _5811_ (.A1(net62),
    .A2(_0967_),
    .B1(_2480_),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _5812_ (.A1(_0490_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][5] ),
    .X(_2481_));
 sky130_fd_sc_hd__a21o_1 _5813_ (.A1(net62),
    .A2(_0996_),
    .B1(_2481_),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _5814_ (.A1(_0536_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][6] ),
    .X(_2482_));
 sky130_fd_sc_hd__a21o_1 _5815_ (.A1(net62),
    .A2(_1028_),
    .B1(_2482_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _5816_ (.A1(_0571_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(\as2650.r123[1][7] ),
    .X(_2483_));
 sky130_fd_sc_hd__a21o_1 _5817_ (.A1(net62),
    .A2(_1068_),
    .B1(_2483_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_8 _5818_ (.A(net207),
    .B(_2831_),
    .Y(_2484_));
 sky130_fd_sc_hd__nor2_8 _5819_ (.A(_2473_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__a22o_1 _5820_ (.A1(net61),
    .A2(_1115_),
    .B1(_2485_),
    .B2(\as2650.r123[2][0] ),
    .X(_2486_));
 sky130_fd_sc_hd__a21o_1 _5821_ (.A1(_2935_),
    .A2(_2484_),
    .B1(_2486_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _5822_ (.A1(net61),
    .A2(_1152_),
    .B1(_2485_),
    .B2(\as2650.r123[2][1] ),
    .X(_2487_));
 sky130_fd_sc_hd__a21o_1 _5823_ (.A1(_2987_),
    .A2(_2484_),
    .B1(_2487_),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _5824_ (.A1(net61),
    .A2(_1179_),
    .B1(_2485_),
    .B2(\as2650.r123[2][2] ),
    .X(_2488_));
 sky130_fd_sc_hd__a21o_1 _5825_ (.A1(_0334_),
    .A2(_2484_),
    .B1(_2488_),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _5826_ (.A1(net61),
    .A2(_1203_),
    .B1(_2485_),
    .B2(\as2650.r123[2][3] ),
    .X(_2489_));
 sky130_fd_sc_hd__a21o_1 _5827_ (.A1(_0386_),
    .A2(_2484_),
    .B1(_2489_),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _5828_ (.A1(net61),
    .A2(_1223_),
    .B1(_2485_),
    .B2(\as2650.r123[2][4] ),
    .X(_2490_));
 sky130_fd_sc_hd__a21o_1 _5829_ (.A1(_0437_),
    .A2(_2484_),
    .B1(_2490_),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _5830_ (.A1(net61),
    .A2(_1237_),
    .B1(_2485_),
    .B2(\as2650.r123[2][5] ),
    .X(_2491_));
 sky130_fd_sc_hd__a21o_1 _5831_ (.A1(_0490_),
    .A2(_2484_),
    .B1(_2491_),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _5832_ (.A1(_0536_),
    .A2(_2484_),
    .B1(_2485_),
    .B2(\as2650.r123[2][6] ),
    .X(_2492_));
 sky130_fd_sc_hd__a21o_1 _5833_ (.A1(net61),
    .A2(_1248_),
    .B1(_2492_),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _5834_ (.A1(_0571_),
    .A2(_2484_),
    .B1(_2485_),
    .B2(\as2650.r123[2][7] ),
    .X(_2493_));
 sky130_fd_sc_hd__a21o_1 _5835_ (.A1(net61),
    .A2(_1251_),
    .B1(_2493_),
    .X(_0277_));
 sky130_fd_sc_hd__o211a_1 _5836_ (.A1(_2765_),
    .A2(net171),
    .B1(net103),
    .C1(_1796_),
    .X(_2494_));
 sky130_fd_sc_hd__o2111a_1 _5837_ (.A1(net136),
    .A2(_0836_),
    .B1(_1329_),
    .C1(_2494_),
    .D1(_2730_),
    .X(_2495_));
 sky130_fd_sc_hd__nor2_1 _5838_ (.A(_1794_),
    .B(_2338_),
    .Y(_2496_));
 sky130_fd_sc_hd__and4_4 _5839_ (.A(_1324_),
    .B(_2330_),
    .C(_2495_),
    .D(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__nor2_4 _5840_ (.A(net233),
    .B(_2780_),
    .Y(_2498_));
 sky130_fd_sc_hd__mux2_8 _5841_ (.A0(_2879_),
    .A1(_2629_),
    .S(net162),
    .X(_2499_));
 sky130_fd_sc_hd__o21ai_1 _5842_ (.A1(net11),
    .A2(net43),
    .B1(net313),
    .Y(_2500_));
 sky130_fd_sc_hd__a21oi_1 _5843_ (.A1(net43),
    .A2(_2499_),
    .B1(_2500_),
    .Y(_0278_));
 sky130_fd_sc_hd__mux2_8 _5844_ (.A0(_2887_),
    .A1(net261),
    .S(net162),
    .X(_2501_));
 sky130_fd_sc_hd__inv_2 _5845_ (.A(_2501_),
    .Y(_2502_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(net43),
    .B(_2502_),
    .Y(_2503_));
 sky130_fd_sc_hd__o211a_1 _5847_ (.A1(net22),
    .A2(net43),
    .B1(_2503_),
    .C1(net313),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_8 _5848_ (.A0(net117),
    .A1(net257),
    .S(net162),
    .X(_2504_));
 sky130_fd_sc_hd__inv_2 _5849_ (.A(_2504_),
    .Y(_2505_));
 sky130_fd_sc_hd__nand2_1 _5850_ (.A(net43),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__o211a_1 _5851_ (.A1(net30),
    .A2(net43),
    .B1(_2506_),
    .C1(net313),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_8 _5852_ (.A0(net113),
    .A1(net254),
    .S(net162),
    .X(_2507_));
 sky130_fd_sc_hd__inv_2 _5853_ (.A(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__nand2_1 _5854_ (.A(net43),
    .B(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__o211a_1 _5855_ (.A1(net31),
    .A2(net43),
    .B1(_2509_),
    .C1(net313),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(net251),
    .B(net162),
    .Y(_2510_));
 sky130_fd_sc_hd__o211ai_4 _5857_ (.A1(_0352_),
    .A2(net162),
    .B1(_2510_),
    .C1(net44),
    .Y(_2511_));
 sky130_fd_sc_hd__o211a_1 _5858_ (.A1(net32),
    .A2(net43),
    .B1(_2511_),
    .C1(net313),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(net250),
    .B(net162),
    .Y(_2512_));
 sky130_fd_sc_hd__o211ai_4 _5860_ (.A1(_0399_),
    .A2(net162),
    .B1(_2512_),
    .C1(net44),
    .Y(_2513_));
 sky130_fd_sc_hd__o211a_1 _5861_ (.A1(net33),
    .A2(net44),
    .B1(_2513_),
    .C1(net313),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _5862_ (.A(net246),
    .B(net162),
    .Y(_2514_));
 sky130_fd_sc_hd__o211ai_4 _5863_ (.A1(_0463_),
    .A2(net162),
    .B1(_2514_),
    .C1(net44),
    .Y(_2515_));
 sky130_fd_sc_hd__o211a_1 _5864_ (.A1(net34),
    .A2(net43),
    .B1(_2515_),
    .C1(net313),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_8 _5865_ (.A0(_2896_),
    .A1(_2628_),
    .S(_2498_),
    .X(_2516_));
 sky130_fd_sc_hd__o21ai_1 _5866_ (.A1(net35),
    .A2(net44),
    .B1(net313),
    .Y(_2517_));
 sky130_fd_sc_hd__a21oi_1 _5867_ (.A1(net44),
    .A2(_2516_),
    .B1(_2517_),
    .Y(_0285_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(net235),
    .A1(net340),
    .S(_0904_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(net230),
    .A1(net339),
    .S(_0904_),
    .X(_0287_));
 sky130_fd_sc_hd__or3b_1 _5870_ (.A(net158),
    .B(_1342_),
    .C_N(net105),
    .X(_2518_));
 sky130_fd_sc_hd__and4_1 _5871_ (.A(_1354_),
    .B(_1369_),
    .C(net53),
    .D(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__o211a_1 _5872_ (.A1(net236),
    .A2(_2790_),
    .B1(net103),
    .C1(_0841_),
    .X(_2520_));
 sky130_fd_sc_hd__o211a_1 _5873_ (.A1(_2672_),
    .A2(_1323_),
    .B1(_2520_),
    .C1(_0835_),
    .X(_2521_));
 sky130_fd_sc_hd__and3_1 _5874_ (.A(_0822_),
    .B(_2519_),
    .C(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__a211o_1 _5875_ (.A1(\as2650.psl[3] ),
    .A2(net140),
    .B1(net128),
    .C1(net238),
    .X(_2523_));
 sky130_fd_sc_hd__and3_1 _5876_ (.A(_1325_),
    .B(_1364_),
    .C(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__a21o_1 _5877_ (.A1(\as2650.psl[3] ),
    .A2(_0838_),
    .B1(_2776_),
    .X(_2525_));
 sky130_fd_sc_hd__and4_1 _5878_ (.A(_1361_),
    .B(_2522_),
    .C(_2524_),
    .D(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__o31a_1 _5879_ (.A1(net337),
    .A2(net70),
    .A3(_0838_),
    .B1(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__a21o_1 _5880_ (.A1(net247),
    .A2(net138),
    .B1(_0764_),
    .X(_2528_));
 sky130_fd_sc_hd__a31o_1 _5881_ (.A1(net127),
    .A2(_1857_),
    .A3(_2528_),
    .B1(_2407_),
    .X(_2529_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(net106),
    .A1(_2529_),
    .S(_2759_),
    .X(_2530_));
 sky130_fd_sc_hd__and2_1 _5883_ (.A(net234),
    .B(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__a21bo_1 _5884_ (.A1(net214),
    .A2(_0434_),
    .B1_N(_2527_),
    .X(_2532_));
 sky130_fd_sc_hd__o221a_1 _5885_ (.A1(\as2650.psl[5] ),
    .A2(_2527_),
    .B1(_2531_),
    .B2(_2532_),
    .C1(net320),
    .X(_0288_));
 sky130_fd_sc_hd__nor2_1 _5886_ (.A(_0568_),
    .B(_0788_),
    .Y(_2533_));
 sky130_fd_sc_hd__nand2_1 _5887_ (.A(_0484_),
    .B(_0489_),
    .Y(_2534_));
 sky130_fd_sc_hd__nor2_1 _5888_ (.A(_0484_),
    .B(_0489_),
    .Y(_2535_));
 sky130_fd_sc_hd__or2_1 _5889_ (.A(_2920_),
    .B(_2934_),
    .X(_2536_));
 sky130_fd_sc_hd__o21a_1 _5890_ (.A1(_2982_),
    .A2(_2536_),
    .B1(_2984_),
    .X(_2537_));
 sky130_fd_sc_hd__a21oi_1 _5891_ (.A1(_2986_),
    .A2(_2536_),
    .B1(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__o21ba_1 _5892_ (.A1(_0369_),
    .A2(_2538_),
    .B1_N(_0333_),
    .X(_2539_));
 sky130_fd_sc_hd__a221o_1 _5893_ (.A1(_0376_),
    .A2(_0382_),
    .B1(_2538_),
    .B2(_0369_),
    .C1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__o22a_1 _5894_ (.A1(_0376_),
    .A2(_0382_),
    .B1(_0418_),
    .B2(_0433_),
    .X(_2541_));
 sky130_fd_sc_hd__a2bb2o_1 _5895_ (.A1_N(_0417_),
    .A2_N(_0434_),
    .B1(_2540_),
    .B2(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__a21oi_1 _5896_ (.A1(_2534_),
    .A2(_2542_),
    .B1(_2535_),
    .Y(_2543_));
 sky130_fd_sc_hd__nor2_1 _5897_ (.A(_0530_),
    .B(_0535_),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _5898_ (.A(_0530_),
    .B(_0535_),
    .Y(_2545_));
 sky130_fd_sc_hd__o221a_1 _5899_ (.A1(_0568_),
    .A2(_0788_),
    .B1(_2543_),
    .B2(_2544_),
    .C1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__and2_1 _5900_ (.A(_0568_),
    .B(_0788_),
    .X(_2547_));
 sky130_fd_sc_hd__o31a_1 _5901_ (.A1(net347),
    .A2(net70),
    .A3(_0838_),
    .B1(_2526_),
    .X(_2548_));
 sky130_fd_sc_hd__a21o_1 _5902_ (.A1(net268),
    .A2(net140),
    .B1(_0764_),
    .X(_2549_));
 sky130_fd_sc_hd__nand3_1 _5903_ (.A(_2774_),
    .B(_1844_),
    .C(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__a21oi_1 _5904_ (.A1(_2773_),
    .A2(net118),
    .B1(_2758_),
    .Y(_2551_));
 sky130_fd_sc_hd__a221o_1 _5905_ (.A1(_2758_),
    .A2(_2879_),
    .B1(_2550_),
    .B2(_2551_),
    .C1(net213),
    .X(_2552_));
 sky130_fd_sc_hd__o311a_1 _5906_ (.A1(net234),
    .A2(_2546_),
    .A3(_2547_),
    .B1(_2548_),
    .C1(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__o21ai_1 _5907_ (.A1(\as2650.carry ),
    .A2(_2548_),
    .B1(net317),
    .Y(_2554_));
 sky130_fd_sc_hd__nor2_1 _5908_ (.A(_2553_),
    .B(_2554_),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_1 _5909_ (.A(_0816_),
    .B(_0830_),
    .Y(_2555_));
 sky130_fd_sc_hd__o221a_1 _5910_ (.A1(_1576_),
    .A2(_1958_),
    .B1(_2555_),
    .B2(net92),
    .C1(_1815_),
    .X(_2556_));
 sky130_fd_sc_hd__or4_1 _5911_ (.A(net238),
    .B(_0747_),
    .C(net70),
    .D(_0757_),
    .X(_2557_));
 sky130_fd_sc_hd__o22a_1 _5912_ (.A1(net172),
    .A2(_2702_),
    .B1(_0767_),
    .B2(_1341_),
    .X(_2558_));
 sky130_fd_sc_hd__a31o_1 _5913_ (.A1(net216),
    .A2(net125),
    .A3(_0752_),
    .B1(net88),
    .X(_2559_));
 sky130_fd_sc_hd__o221a_1 _5914_ (.A1(net292),
    .A2(_2669_),
    .B1(net198),
    .B2(_2788_),
    .C1(net218),
    .X(_2560_));
 sky130_fd_sc_hd__a21oi_1 _5915_ (.A1(net299),
    .A2(net154),
    .B1(net98),
    .Y(_2561_));
 sky130_fd_sc_hd__a31oi_1 _5916_ (.A1(net236),
    .A2(net98),
    .A3(_0581_),
    .B1(_2561_),
    .Y(_2562_));
 sky130_fd_sc_hd__o221a_1 _5917_ (.A1(net236),
    .A2(net71),
    .B1(_1404_),
    .B2(_1799_),
    .C1(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__o211a_1 _5918_ (.A1(net158),
    .A2(_0764_),
    .B1(_2560_),
    .C1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__and3_1 _5919_ (.A(_1369_),
    .B(_2559_),
    .C(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__and4bb_1 _5920_ (.A_N(_1961_),
    .B_N(_1964_),
    .C(_2558_),
    .D(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__and3_4 _5921_ (.A(_2556_),
    .B(_2557_),
    .C(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__o21a_1 _5922_ (.A1(net343),
    .A2(_1341_),
    .B1(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__a21o_1 _5923_ (.A1(net343),
    .A2(_0775_),
    .B1(net139),
    .X(_2569_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(net228),
    .B(net192),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2_1 _5925_ (.A(_0897_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(net257),
    .A1(_2571_),
    .S(_0586_),
    .X(_2572_));
 sky130_fd_sc_hd__o31a_1 _5927_ (.A1(net90),
    .A2(net76),
    .A3(_2572_),
    .B1(_2569_),
    .X(_2573_));
 sky130_fd_sc_hd__nor2_2 _5928_ (.A(_2845_),
    .B(net163),
    .Y(_2574_));
 sky130_fd_sc_hd__o221a_1 _5929_ (.A1(net163),
    .A2(_2573_),
    .B1(_2574_),
    .B2(net122),
    .C1(net215),
    .X(_2575_));
 sky130_fd_sc_hd__a21oi_1 _5930_ (.A1(net237),
    .A2(_2571_),
    .B1(_2575_),
    .Y(_2576_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(net219),
    .A1(_2576_),
    .S(_2568_),
    .X(_2577_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(net325),
    .B(_2577_),
    .Y(_0290_));
 sky130_fd_sc_hd__o21a_1 _5933_ (.A1(net346),
    .A2(_1341_),
    .B1(_2567_),
    .X(_2578_));
 sky130_fd_sc_hd__nor2_1 _5934_ (.A(net138),
    .B(_0775_),
    .Y(_2579_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(net261),
    .A1(_2855_),
    .S(_0586_),
    .X(_2580_));
 sky130_fd_sc_hd__or3_1 _5936_ (.A(net90),
    .B(net76),
    .C(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__o211a_1 _5937_ (.A1(net139),
    .A2(_0775_),
    .B1(_1845_),
    .C1(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__o221a_1 _5938_ (.A1(_2856_),
    .A2(_2574_),
    .B1(_2582_),
    .B2(net163),
    .C1(net215),
    .X(_2583_));
 sky130_fd_sc_hd__a21o_1 _5939_ (.A1(net237),
    .A2(_2855_),
    .B1(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(net226),
    .A1(_2584_),
    .S(_2578_),
    .X(_2585_));
 sky130_fd_sc_hd__and2_1 _5941_ (.A(net319),
    .B(_2585_),
    .X(_0291_));
 sky130_fd_sc_hd__o21a_1 _5942_ (.A1(net348),
    .A2(_1341_),
    .B1(_2567_),
    .X(_2586_));
 sky130_fd_sc_hd__or3_1 _5943_ (.A(net76),
    .B(_0586_),
    .C(net104),
    .X(_2587_));
 sky130_fd_sc_hd__o311a_2 _5944_ (.A1(net304),
    .A2(net199),
    .A3(_2806_),
    .B1(net138),
    .C1(net265),
    .X(_2588_));
 sky130_fd_sc_hd__a31o_1 _5945_ (.A1(net348),
    .A2(net135),
    .A3(_0775_),
    .B1(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__a32o_1 _5946_ (.A1(_2626_),
    .A2(_1341_),
    .A3(_2587_),
    .B1(_2589_),
    .B2(_0814_),
    .X(_2590_));
 sky130_fd_sc_hd__mux2_1 _5947_ (.A0(\as2650.psu[0] ),
    .A1(_2590_),
    .S(_2586_),
    .X(_2591_));
 sky130_fd_sc_hd__and2_1 _5948_ (.A(net319),
    .B(_2591_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _5949_ (.A(_2533_),
    .B(_2547_),
    .X(_2592_));
 sky130_fd_sc_hd__o221a_1 _5950_ (.A1(net238),
    .A2(_0748_),
    .B1(_0838_),
    .B2(net344),
    .C1(_1325_),
    .X(_2593_));
 sky130_fd_sc_hd__nand3_2 _5951_ (.A(_0756_),
    .B(_2522_),
    .C(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__a21o_1 _5952_ (.A1(net260),
    .A2(net138),
    .B1(_0764_),
    .X(_2595_));
 sky130_fd_sc_hd__a31o_1 _5953_ (.A1(net234),
    .A2(_1848_),
    .A3(_2595_),
    .B1(_2594_),
    .X(_2596_));
 sky130_fd_sc_hd__a31o_1 _5954_ (.A1(net214),
    .A2(_0556_),
    .A3(_2592_),
    .B1(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__nand2_1 _5955_ (.A(_2625_),
    .B(_2594_),
    .Y(_2598_));
 sky130_fd_sc_hd__and3_1 _5956_ (.A(net320),
    .B(_2597_),
    .C(_2598_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _5957_ (.A(net305),
    .B(net140),
    .Y(_2599_));
 sky130_fd_sc_hd__a211o_1 _5958_ (.A1(net161),
    .A2(net105),
    .B1(net142),
    .C1(net296),
    .X(_2600_));
 sky130_fd_sc_hd__nor2_1 _5959_ (.A(net88),
    .B(_0771_),
    .Y(_2601_));
 sky130_fd_sc_hd__a211o_1 _5960_ (.A1(net161),
    .A2(net105),
    .B1(net142),
    .C1(net296),
    .X(_2602_));
 sky130_fd_sc_hd__or4_1 _5961_ (.A(_0774_),
    .B(_0833_),
    .C(_2599_),
    .D(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__a21o_4 _5962_ (.A1(net138),
    .A2(_0820_),
    .B1(_2603_),
    .X(_2604_));
 sky130_fd_sc_hd__inv_2 _5963_ (.A(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__o21ai_1 _5964_ (.A1(_1853_),
    .A2(_2604_),
    .B1(net223),
    .Y(_2606_));
 sky130_fd_sc_hd__o31a_1 _5965_ (.A1(_2655_),
    .A2(net138),
    .A3(_0763_),
    .B1(_1854_),
    .X(_2607_));
 sky130_fd_sc_hd__or2_1 _5966_ (.A(_2604_),
    .B(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__a21oi_1 _5967_ (.A1(_2606_),
    .A2(_2608_),
    .B1(net323),
    .Y(_0294_));
 sky130_fd_sc_hd__o21ai_1 _5968_ (.A1(_1849_),
    .A2(_2604_),
    .B1(\as2650.psl[3] ),
    .Y(_2609_));
 sky130_fd_sc_hd__o31a_1 _5969_ (.A1(_2654_),
    .A2(net136),
    .A3(_0763_),
    .B1(_1850_),
    .X(_2610_));
 sky130_fd_sc_hd__or2_1 _5970_ (.A(_2604_),
    .B(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__a21oi_1 _5971_ (.A1(_2609_),
    .A2(_2611_),
    .B1(net323),
    .Y(_0295_));
 sky130_fd_sc_hd__a21o_1 _5972_ (.A1(_1845_),
    .A2(_2605_),
    .B1(\as2650.psl[1] ),
    .X(_2612_));
 sky130_fd_sc_hd__o31a_1 _5973_ (.A1(_2652_),
    .A2(net139),
    .A3(_0764_),
    .B1(_1846_),
    .X(_2613_));
 sky130_fd_sc_hd__o211a_1 _5974_ (.A1(_2604_),
    .A2(_2613_),
    .B1(_2612_),
    .C1(net320),
    .X(_0296_));
 sky130_fd_sc_hd__o21ai_1 _5975_ (.A1(net88),
    .A2(_0759_),
    .B1(_2803_),
    .Y(_2614_));
 sky130_fd_sc_hd__or4_4 _5976_ (.A(net305),
    .B(_2600_),
    .C(_2601_),
    .D(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__a21oi_1 _5977_ (.A1(_2658_),
    .A2(net88),
    .B1(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__or2_1 _5978_ (.A(net29),
    .B(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__o2bb2a_1 _5979_ (.A1_N(net335),
    .A2_N(_2579_),
    .B1(net88),
    .B2(net246),
    .X(_2618_));
 sky130_fd_sc_hd__o211a_1 _5980_ (.A1(_2615_),
    .A2(_2618_),
    .B1(_2617_),
    .C1(net317),
    .X(_0297_));
 sky130_fd_sc_hd__o21ai_1 _5981_ (.A1(_1853_),
    .A2(_2615_),
    .B1(\as2650.psu[4] ),
    .Y(_2619_));
 sky130_fd_sc_hd__or3_1 _5982_ (.A(_1855_),
    .B(_2579_),
    .C(_2615_),
    .X(_2620_));
 sky130_fd_sc_hd__a21oi_1 _5983_ (.A1(_2619_),
    .A2(_2620_),
    .B1(net323),
    .Y(_0298_));
 sky130_fd_sc_hd__o21ai_1 _5984_ (.A1(_1849_),
    .A2(_2615_),
    .B1(\as2650.psu[3] ),
    .Y(_2621_));
 sky130_fd_sc_hd__or3_1 _5985_ (.A(_1851_),
    .B(_2579_),
    .C(_2615_),
    .X(_2622_));
 sky130_fd_sc_hd__a21oi_1 _5986_ (.A1(_2621_),
    .A2(_2622_),
    .B1(net323),
    .Y(_0299_));
 sky130_fd_sc_hd__clkbuf_2 _5987_ (.A(\as2650.r123_2[3][0] ),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_2 _5988_ (.A(\as2650.r123_2[3][1] ),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_2 _5989_ (.A(\as2650.r123_2[3][2] ),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_2 _5990_ (.A(\as2650.r123_2[3][3] ),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_2 _5991_ (.A(\as2650.r123_2[3][4] ),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_2 _5992_ (.A(\as2650.r123_2[3][5] ),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_2 _5993_ (.A(\as2650.r123_2[3][6] ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_2 _5994_ (.A(\as2650.r123_2[3][7] ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _5995_ (.A(\as2650.r123[3][0] ),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_2 _5996_ (.A(\as2650.r123[3][1] ),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_2 _5997_ (.A(\as2650.r123[3][2] ),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_2 _5998_ (.A(\as2650.r123[3][3] ),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_2 _5999_ (.A(\as2650.r123[3][4] ),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_2 _6000_ (.A(\as2650.r123[3][5] ),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_2 _6001_ (.A(\as2650.r123[3][6] ),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_2 _6002_ (.A(\as2650.r123[3][7] ),
    .X(_0145_));
 sky130_fd_sc_hd__dfxtp_2 _6003_ (.CLK(clknet_leaf_6_clk),
    .D(_0000_),
    .Q(\as2650.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6004_ (.CLK(clknet_leaf_4_clk),
    .D(_0001_),
    .Q(\as2650.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6005_ (.CLK(clknet_leaf_4_clk),
    .D(_0002_),
    .Q(\as2650.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6006_ (.CLK(clknet_leaf_4_clk),
    .D(_0003_),
    .Q(\as2650.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6007_ (.CLK(clknet_leaf_4_clk),
    .D(_0004_),
    .Q(\as2650.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6008_ (.CLK(clknet_leaf_9_clk),
    .D(_0005_),
    .Q(\as2650.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6009_ (.CLK(clknet_leaf_9_clk),
    .D(_0006_),
    .Q(\as2650.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6010_ (.CLK(clknet_leaf_6_clk),
    .D(_0007_),
    .Q(\as2650.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_4 _6011_ (.CLK(clknet_leaf_25_clk),
    .D(_0008_),
    .Q(\as2650.r123[0][0] ));
 sky130_fd_sc_hd__dfxtp_4 _6012_ (.CLK(clknet_leaf_24_clk),
    .D(_0009_),
    .Q(\as2650.r123[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _6013_ (.CLK(clknet_leaf_26_clk),
    .D(_0010_),
    .Q(\as2650.r123[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _6014_ (.CLK(clknet_leaf_25_clk),
    .D(_0011_),
    .Q(\as2650.r123[0][3] ));
 sky130_fd_sc_hd__dfxtp_4 _6015_ (.CLK(clknet_leaf_25_clk),
    .D(_0012_),
    .Q(\as2650.r123[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _6016_ (.CLK(clknet_leaf_25_clk),
    .D(_0013_),
    .Q(\as2650.r123[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _6017_ (.CLK(clknet_leaf_25_clk),
    .D(_0014_),
    .Q(\as2650.r123[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6018_ (.CLK(clknet_leaf_24_clk),
    .D(_0015_),
    .Q(\as2650.r123[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6019_ (.CLK(clknet_leaf_41_clk),
    .D(_0016_),
    .Q(\as2650.stack[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6020_ (.CLK(clknet_leaf_48_clk),
    .D(_0017_),
    .Q(\as2650.stack[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6021_ (.CLK(clknet_leaf_47_clk),
    .D(_0018_),
    .Q(\as2650.stack[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6022_ (.CLK(clknet_leaf_50_clk),
    .D(_0019_),
    .Q(\as2650.stack[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6023_ (.CLK(clknet_leaf_47_clk),
    .D(_0020_),
    .Q(\as2650.stack[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6024_ (.CLK(clknet_leaf_41_clk),
    .D(_0021_),
    .Q(\as2650.stack[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6025_ (.CLK(clknet_leaf_38_clk),
    .D(_0022_),
    .Q(\as2650.stack[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6026_ (.CLK(clknet_leaf_48_clk),
    .D(_0023_),
    .Q(\as2650.stack[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6027_ (.CLK(clknet_leaf_43_clk),
    .D(_0024_),
    .Q(\as2650.stack[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6028_ (.CLK(clknet_leaf_44_clk),
    .D(_0025_),
    .Q(\as2650.stack[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6029_ (.CLK(clknet_leaf_42_clk),
    .D(_0026_),
    .Q(\as2650.stack[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6030_ (.CLK(clknet_leaf_30_clk),
    .D(_0027_),
    .Q(\as2650.stack[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6031_ (.CLK(clknet_leaf_43_clk),
    .D(_0028_),
    .Q(\as2650.stack[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6032_ (.CLK(clknet_leaf_25_clk),
    .D(_0029_),
    .Q(\as2650.stack[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6033_ (.CLK(clknet_leaf_30_clk),
    .D(_0030_),
    .Q(\as2650.stack[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6034_ (.CLK(clknet_leaf_26_clk),
    .D(_0031_),
    .Q(\as2650.r123_2[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6035_ (.CLK(clknet_leaf_21_clk),
    .D(_0032_),
    .Q(\as2650.r123_2[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6036_ (.CLK(clknet_leaf_26_clk),
    .D(_0033_),
    .Q(\as2650.r123_2[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6037_ (.CLK(clknet_leaf_26_clk),
    .D(_0034_),
    .Q(\as2650.r123_2[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6038_ (.CLK(clknet_leaf_27_clk),
    .D(_0035_),
    .Q(\as2650.r123_2[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6039_ (.CLK(clknet_leaf_24_clk),
    .D(_0036_),
    .Q(\as2650.r123_2[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6040_ (.CLK(clknet_leaf_22_clk),
    .D(_0037_),
    .Q(\as2650.r123_2[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6041_ (.CLK(clknet_leaf_24_clk),
    .D(_0038_),
    .Q(\as2650.r123_2[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6042_ (.CLK(clknet_leaf_12_clk),
    .D(_0039_),
    .Q(\as2650.psu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6043_ (.CLK(clknet_leaf_43_clk),
    .D(_0040_),
    .Q(\as2650.stack[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6044_ (.CLK(clknet_leaf_44_clk),
    .D(_0041_),
    .Q(\as2650.stack[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6045_ (.CLK(clknet_leaf_41_clk),
    .D(_0042_),
    .Q(\as2650.stack[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6046_ (.CLK(clknet_leaf_42_clk),
    .D(_0043_),
    .Q(\as2650.stack[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6047_ (.CLK(clknet_leaf_44_clk),
    .D(_0044_),
    .Q(\as2650.stack[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6048_ (.CLK(clknet_leaf_43_clk),
    .D(_0045_),
    .Q(\as2650.stack[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6049_ (.CLK(clknet_leaf_36_clk),
    .D(_0046_),
    .Q(\as2650.stack[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6050_ (.CLK(clknet_leaf_42_clk),
    .D(_0047_),
    .Q(\as2650.stack[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6051_ (.CLK(clknet_leaf_41_clk),
    .D(_0048_),
    .Q(\as2650.stack[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6052_ (.CLK(clknet_leaf_42_clk),
    .D(_0049_),
    .Q(\as2650.stack[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6053_ (.CLK(clknet_leaf_35_clk),
    .D(_0050_),
    .Q(\as2650.stack[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6054_ (.CLK(clknet_leaf_42_clk),
    .D(_0051_),
    .Q(\as2650.stack[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6055_ (.CLK(clknet_leaf_25_clk),
    .D(_0052_),
    .Q(\as2650.stack[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6056_ (.CLK(clknet_leaf_36_clk),
    .D(_0053_),
    .Q(\as2650.stack[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _6057_ (.CLK(clknet_leaf_15_clk),
    .D(_0054_),
    .Q(\as2650.psl[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6058_ (.CLK(clknet_leaf_11_clk),
    .D(_0055_),
    .Q(\as2650.psl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6059_ (.CLK(clknet_leaf_36_clk),
    .D(_0056_),
    .Q(\as2650.stack[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6060_ (.CLK(clknet_leaf_38_clk),
    .D(_0057_),
    .Q(\as2650.stack[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6061_ (.CLK(clknet_leaf_37_clk),
    .D(_0058_),
    .Q(\as2650.stack[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6062_ (.CLK(clknet_leaf_34_clk),
    .D(_0059_),
    .Q(\as2650.stack[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6063_ (.CLK(clknet_leaf_40_clk),
    .D(_0060_),
    .Q(\as2650.stack[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6064_ (.CLK(clknet_leaf_35_clk),
    .D(_0061_),
    .Q(\as2650.stack[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6065_ (.CLK(clknet_leaf_34_clk),
    .D(_0062_),
    .Q(\as2650.stack[3][14] ));
 sky130_fd_sc_hd__dfxtp_4 _6066_ (.CLK(clknet_leaf_8_clk),
    .D(_0063_),
    .Q(\as2650.ins_reg[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6067_ (.CLK(clknet_leaf_9_clk),
    .D(_0064_),
    .Q(\as2650.ins_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6068_ (.CLK(clknet_leaf_8_clk),
    .D(_0065_),
    .Q(\as2650.ins_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6069_ (.CLK(clknet_leaf_9_clk),
    .D(_0066_),
    .Q(\as2650.ins_reg[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6070_ (.CLK(clknet_leaf_8_clk),
    .D(_0067_),
    .Q(\as2650.ins_reg[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6071_ (.CLK(clknet_leaf_9_clk),
    .D(_0068_),
    .Q(\as2650.ins_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6072_ (.CLK(clknet_leaf_36_clk),
    .D(_0069_),
    .Q(\as2650.stack[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6073_ (.CLK(clknet_leaf_38_clk),
    .D(_0070_),
    .Q(\as2650.stack[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6074_ (.CLK(clknet_leaf_37_clk),
    .D(_0071_),
    .Q(\as2650.stack[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6075_ (.CLK(clknet_leaf_36_clk),
    .D(_0072_),
    .Q(\as2650.stack[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6076_ (.CLK(clknet_leaf_42_clk),
    .D(_0073_),
    .Q(\as2650.stack[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6077_ (.CLK(clknet_leaf_35_clk),
    .D(_0074_),
    .Q(\as2650.stack[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6078_ (.CLK(clknet_leaf_34_clk),
    .D(_0075_),
    .Q(\as2650.stack[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6079_ (.CLK(clknet_leaf_22_clk),
    .D(_0076_),
    .Q(\as2650.r123_2[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6080_ (.CLK(clknet_leaf_19_clk),
    .D(_0077_),
    .Q(\as2650.r123_2[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6081_ (.CLK(clknet_leaf_19_clk),
    .D(_0078_),
    .Q(\as2650.r123_2[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6082_ (.CLK(clknet_leaf_20_clk),
    .D(_0079_),
    .Q(\as2650.r123_2[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6083_ (.CLK(clknet_leaf_19_clk),
    .D(_0080_),
    .Q(\as2650.r123_2[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6084_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0081_),
    .Q(\as2650.r123_2[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6085_ (.CLK(clknet_leaf_21_clk),
    .D(_0082_),
    .Q(\as2650.r123_2[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6086_ (.CLK(clknet_leaf_19_clk),
    .D(_0083_),
    .Q(\as2650.r123_2[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6087_ (.CLK(clknet_leaf_36_clk),
    .D(_0084_),
    .Q(\as2650.stack[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6088_ (.CLK(clknet_leaf_38_clk),
    .D(_0085_),
    .Q(\as2650.stack[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6089_ (.CLK(clknet_leaf_37_clk),
    .D(_0086_),
    .Q(\as2650.stack[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6090_ (.CLK(clknet_leaf_34_clk),
    .D(_0087_),
    .Q(\as2650.stack[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6091_ (.CLK(clknet_leaf_38_clk),
    .D(_0088_),
    .Q(\as2650.stack[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6092_ (.CLK(clknet_leaf_36_clk),
    .D(_0089_),
    .Q(\as2650.stack[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6093_ (.CLK(clknet_leaf_34_clk),
    .D(_0090_),
    .Q(\as2650.stack[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6094_ (.CLK(clknet_leaf_36_clk),
    .D(_0091_),
    .Q(\as2650.stack[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6095_ (.CLK(clknet_leaf_37_clk),
    .D(_0092_),
    .Q(\as2650.stack[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6096_ (.CLK(clknet_leaf_37_clk),
    .D(_0093_),
    .Q(\as2650.stack[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6097_ (.CLK(clknet_leaf_37_clk),
    .D(_0094_),
    .Q(\as2650.stack[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6098_ (.CLK(clknet_leaf_37_clk),
    .D(_0095_),
    .Q(\as2650.stack[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6099_ (.CLK(clknet_leaf_36_clk),
    .D(_0096_),
    .Q(\as2650.stack[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6100_ (.CLK(clknet_leaf_36_clk),
    .D(_0097_),
    .Q(\as2650.stack[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6101_ (.CLK(clknet_leaf_54_clk),
    .D(_0098_),
    .Q(\as2650.r123_2[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6102_ (.CLK(clknet_leaf_32_clk),
    .D(_0099_),
    .Q(\as2650.r123_2[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6103_ (.CLK(clknet_leaf_54_clk),
    .D(_0100_),
    .Q(\as2650.r123_2[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6104_ (.CLK(clknet_leaf_32_clk),
    .D(_0101_),
    .Q(\as2650.r123_2[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6105_ (.CLK(clknet_leaf_32_clk),
    .D(_0102_),
    .Q(\as2650.r123_2[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6106_ (.CLK(clknet_leaf_32_clk),
    .D(_0103_),
    .Q(\as2650.r123_2[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6107_ (.CLK(clknet_leaf_32_clk),
    .D(_0104_),
    .Q(\as2650.r123_2[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6108_ (.CLK(clknet_leaf_33_clk),
    .D(_0105_),
    .Q(\as2650.r123_2[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6109_ (.CLK(clknet_leaf_20_clk),
    .D(_0106_),
    .Q(\as2650.r123_2[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6110_ (.CLK(clknet_leaf_20_clk),
    .D(_0107_),
    .Q(\as2650.r123_2[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_28_clk),
    .D(_0108_),
    .Q(\as2650.r123_2[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6112_ (.CLK(clknet_leaf_28_clk),
    .D(_0109_),
    .Q(\as2650.r123_2[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6113_ (.CLK(clknet_leaf_28_clk),
    .D(_0110_),
    .Q(\as2650.r123_2[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6114_ (.CLK(clknet_leaf_26_clk),
    .D(_0111_),
    .Q(\as2650.r123_2[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6115_ (.CLK(clknet_leaf_27_clk),
    .D(_0112_),
    .Q(\as2650.r123_2[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6116_ (.CLK(clknet_leaf_27_clk),
    .D(_0113_),
    .Q(\as2650.r123_2[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6117_ (.CLK(clknet_leaf_40_clk),
    .D(_0114_),
    .Q(\as2650.stack[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6118_ (.CLK(clknet_leaf_39_clk),
    .D(_0115_),
    .Q(\as2650.stack[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6119_ (.CLK(clknet_leaf_49_clk),
    .D(_0116_),
    .Q(\as2650.stack[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6120_ (.CLK(clknet_leaf_49_clk),
    .D(_0117_),
    .Q(\as2650.stack[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6121_ (.CLK(clknet_leaf_47_clk),
    .D(_0118_),
    .Q(\as2650.stack[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6122_ (.CLK(clknet_leaf_40_clk),
    .D(_0119_),
    .Q(\as2650.stack[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6123_ (.CLK(clknet_leaf_38_clk),
    .D(_0120_),
    .Q(\as2650.stack[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6124_ (.CLK(clknet_leaf_48_clk),
    .D(_0121_),
    .Q(\as2650.stack[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6125_ (.CLK(clknet_leaf_46_clk),
    .D(_0122_),
    .Q(\as2650.stack[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6126_ (.CLK(clknet_leaf_49_clk),
    .D(_0123_),
    .Q(\as2650.stack[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6127_ (.CLK(clknet_leaf_51_clk),
    .D(_0124_),
    .Q(\as2650.stack[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6128_ (.CLK(clknet_leaf_51_clk),
    .D(_0125_),
    .Q(\as2650.stack[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6129_ (.CLK(clknet_leaf_50_clk),
    .D(_0126_),
    .Q(\as2650.stack[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6130_ (.CLK(clknet_leaf_50_clk),
    .D(_0127_),
    .Q(\as2650.stack[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6131_ (.CLK(clknet_leaf_49_clk),
    .D(_0128_),
    .Q(\as2650.stack[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6132_ (.CLK(clknet_leaf_52_clk),
    .D(_0129_),
    .Q(\as2650.stack[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6133_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0130_),
    .Q(\as2650.stack[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6134_ (.CLK(clknet_leaf_53_clk),
    .D(_0131_),
    .Q(\as2650.stack[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6135_ (.CLK(clknet_leaf_55_clk),
    .D(_0132_),
    .Q(\as2650.stack[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6136_ (.CLK(clknet_leaf_52_clk),
    .D(_0133_),
    .Q(\as2650.stack[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6137_ (.CLK(clknet_leaf_51_clk),
    .D(_0134_),
    .Q(\as2650.stack[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6138_ (.CLK(clknet_leaf_54_clk),
    .D(_0135_),
    .Q(\as2650.stack[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6139_ (.CLK(clknet_leaf_53_clk),
    .D(_0136_),
    .Q(\as2650.stack[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6140_ (.CLK(clknet_leaf_54_clk),
    .D(_0137_),
    .Q(\as2650.stack[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6141_ (.CLK(clknet_leaf_33_clk),
    .D(_0138_),
    .Q(\as2650.r123[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_54_clk),
    .D(_0139_),
    .Q(\as2650.r123[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6143_ (.CLK(clknet_leaf_32_clk),
    .D(_0140_),
    .Q(\as2650.r123[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_33_clk),
    .D(_0141_),
    .Q(\as2650.r123[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6145_ (.CLK(clknet_leaf_54_clk),
    .D(_0142_),
    .Q(\as2650.r123[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(clknet_leaf_54_clk),
    .D(_0143_),
    .Q(\as2650.r123[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(clknet_leaf_54_clk),
    .D(_0144_),
    .Q(\as2650.r123[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(clknet_leaf_54_clk),
    .D(_0145_),
    .Q(\as2650.r123[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_50_clk),
    .D(_0146_),
    .Q(\as2650.stack[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6150_ (.CLK(clknet_leaf_49_clk),
    .D(_0147_),
    .Q(\as2650.stack[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6151_ (.CLK(clknet_leaf_50_clk),
    .D(_0148_),
    .Q(\as2650.stack[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6152_ (.CLK(clknet_leaf_52_clk),
    .D(_0149_),
    .Q(\as2650.stack[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6153_ (.CLK(clknet_leaf_50_clk),
    .D(_0150_),
    .Q(\as2650.stack[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6154_ (.CLK(clknet_leaf_50_clk),
    .D(_0151_),
    .Q(\as2650.stack[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6155_ (.CLK(clknet_leaf_49_clk),
    .D(_0152_),
    .Q(\as2650.stack[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6156_ (.CLK(clknet_leaf_53_clk),
    .D(_0153_),
    .Q(\as2650.stack[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _6157_ (.CLK(clknet_leaf_30_clk),
    .D(_0154_),
    .Q(\lfsr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6158_ (.CLK(clknet_leaf_30_clk),
    .D(_0155_),
    .Q(\lfsr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6159_ (.CLK(clknet_leaf_30_clk),
    .D(_0156_),
    .Q(\lfsr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6160_ (.CLK(clknet_leaf_30_clk),
    .D(_0157_),
    .Q(\lfsr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6161_ (.CLK(clknet_leaf_30_clk),
    .D(_0158_),
    .Q(\lfsr[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6162_ (.CLK(clknet_leaf_29_clk),
    .D(_0159_),
    .Q(\as2650.sense ));
 sky130_fd_sc_hd__dfxtp_1 _6163_ (.CLK(clknet_leaf_29_clk),
    .D(_0160_),
    .Q(\lfsr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6164_ (.CLK(clknet_leaf_29_clk),
    .D(_0161_),
    .Q(\lfsr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6165_ (.CLK(clknet_leaf_30_clk),
    .D(_0162_),
    .Q(\lfsr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6166_ (.CLK(clknet_leaf_31_clk),
    .D(_0163_),
    .Q(\lfsr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6167_ (.CLK(clknet_leaf_31_clk),
    .D(_0164_),
    .Q(\lfsr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6168_ (.CLK(clknet_leaf_31_clk),
    .D(_0165_),
    .Q(\lfsr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6169_ (.CLK(clknet_leaf_31_clk),
    .D(_0166_),
    .Q(\lfsr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6170_ (.CLK(clknet_leaf_31_clk),
    .D(_0167_),
    .Q(\lfsr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6171_ (.CLK(clknet_leaf_35_clk),
    .D(_0168_),
    .Q(\lfsr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6172_ (.CLK(clknet_leaf_35_clk),
    .D(_0169_),
    .Q(\lfsr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6173_ (.CLK(clknet_leaf_51_clk),
    .D(_0170_),
    .Q(\as2650.stack[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6174_ (.CLK(clknet_leaf_53_clk),
    .D(_0171_),
    .Q(\as2650.stack[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6175_ (.CLK(clknet_leaf_55_clk),
    .D(_0172_),
    .Q(\as2650.stack[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6176_ (.CLK(clknet_leaf_52_clk),
    .D(_0173_),
    .Q(\as2650.stack[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6177_ (.CLK(clknet_leaf_51_clk),
    .D(_0174_),
    .Q(\as2650.stack[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6178_ (.CLK(clknet_leaf_55_clk),
    .D(_0175_),
    .Q(\as2650.stack[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6179_ (.CLK(clknet_leaf_53_clk),
    .D(_0176_),
    .Q(\as2650.stack[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6180_ (.CLK(clknet_leaf_54_clk),
    .D(_0177_),
    .Q(\as2650.stack[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6181_ (.CLK(clknet_leaf_7_clk),
    .D(_0178_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _6182_ (.CLK(clknet_leaf_8_clk),
    .D(_0179_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _6183_ (.CLK(clknet_leaf_8_clk),
    .D(_0180_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_4 _6184_ (.CLK(clknet_leaf_5_clk),
    .D(_0181_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_4 _6185_ (.CLK(clknet_leaf_0_clk),
    .D(_0182_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _6186_ (.CLK(clknet_leaf_1_clk),
    .D(_0183_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_2 _6187_ (.CLK(clknet_leaf_5_clk),
    .D(_0184_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_2 _6188_ (.CLK(clknet_leaf_5_clk),
    .D(_0185_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_4 _6189_ (.CLK(clknet_leaf_0_clk),
    .D(_0186_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_4 _6190_ (.CLK(clknet_leaf_0_clk),
    .D(_0187_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_4 _6191_ (.CLK(clknet_leaf_6_clk),
    .D(_0188_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_4 _6192_ (.CLK(clknet_leaf_0_clk),
    .D(_0189_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_2 _6193_ (.CLK(clknet_leaf_5_clk),
    .D(_0190_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_4 _6194_ (.CLK(clknet_leaf_0_clk),
    .D(_0191_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_4 _6195_ (.CLK(clknet_leaf_0_clk),
    .D(_0192_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_4 _6196_ (.CLK(clknet_leaf_1_clk),
    .D(_0193_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_2 _6197_ (.CLK(clknet_leaf_8_clk),
    .D(_0194_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_4 _6198_ (.CLK(clknet_leaf_6_clk),
    .D(_0195_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 _6199_ (.CLK(clknet_leaf_10_clk),
    .D(_0196_),
    .Q(\as2650.idx_ctrl[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6200_ (.CLK(clknet_leaf_10_clk),
    .D(_0197_),
    .Q(\as2650.idx_ctrl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6201_ (.CLK(clknet_leaf_15_clk),
    .D(_0198_),
    .Q(\as2650.holding_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6202_ (.CLK(clknet_leaf_16_clk),
    .D(_0199_),
    .Q(\as2650.holding_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6203_ (.CLK(clknet_leaf_15_clk),
    .D(_0200_),
    .Q(\as2650.holding_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6204_ (.CLK(clknet_leaf_15_clk),
    .D(_0201_),
    .Q(\as2650.holding_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6205_ (.CLK(clknet_leaf_10_clk),
    .D(_0202_),
    .Q(\as2650.holding_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6206_ (.CLK(clknet_leaf_15_clk),
    .D(_0203_),
    .Q(\as2650.holding_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6207_ (.CLK(clknet_leaf_10_clk),
    .D(_0204_),
    .Q(\as2650.holding_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6208_ (.CLK(clknet_leaf_10_clk),
    .D(_0205_),
    .Q(\as2650.holding_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6209_ (.CLK(clknet_leaf_9_clk),
    .D(_0206_),
    .Q(\as2650.halted ));
 sky130_fd_sc_hd__dfxtp_1 _6210_ (.CLK(clknet_leaf_7_clk),
    .D(_0207_),
    .Q(\as2650.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6211_ (.CLK(clknet_leaf_7_clk),
    .D(_0208_),
    .Q(\as2650.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6212_ (.CLK(clknet_leaf_7_clk),
    .D(_0209_),
    .Q(\as2650.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6213_ (.CLK(clknet_leaf_7_clk),
    .D(_0210_),
    .Q(\as2650.cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6214_ (.CLK(clknet_leaf_7_clk),
    .D(_0211_),
    .Q(\as2650.cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6215_ (.CLK(clknet_leaf_6_clk),
    .D(_0212_),
    .Q(\as2650.cycle[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6216_ (.CLK(clknet_leaf_6_clk),
    .D(_0213_),
    .Q(\as2650.cycle[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6217_ (.CLK(clknet_leaf_6_clk),
    .D(_0214_),
    .Q(\as2650.cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6218_ (.CLK(clknet_leaf_12_clk),
    .D(_0215_),
    .Q(\as2650.psu[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6219_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0216_),
    .Q(\as2650.pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6220_ (.CLK(clknet_leaf_45_clk),
    .D(_0217_),
    .Q(\as2650.pc[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6221_ (.CLK(clknet_leaf_46_clk),
    .D(_0218_),
    .Q(\as2650.pc[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6222_ (.CLK(clknet_leaf_46_clk),
    .D(_0219_),
    .Q(\as2650.pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6223_ (.CLK(clknet_leaf_47_clk),
    .D(_0220_),
    .Q(\as2650.pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6224_ (.CLK(clknet_leaf_46_clk),
    .D(_0221_),
    .Q(\as2650.pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6225_ (.CLK(clknet_leaf_44_clk),
    .D(_0222_),
    .Q(\as2650.pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6226_ (.CLK(clknet_leaf_47_clk),
    .D(_0223_),
    .Q(\as2650.pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6227_ (.CLK(clknet_leaf_46_clk),
    .D(_0224_),
    .Q(\as2650.pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6228_ (.CLK(clknet_leaf_44_clk),
    .D(_0225_),
    .Q(\as2650.pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6229_ (.CLK(clknet_leaf_44_clk),
    .D(_0226_),
    .Q(\as2650.pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6230_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0227_),
    .Q(\as2650.pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6231_ (.CLK(clknet_leaf_45_clk),
    .D(_0228_),
    .Q(\as2650.pc[12] ));
 sky130_fd_sc_hd__dfxtp_4 _6232_ (.CLK(clknet_leaf_45_clk),
    .D(_0229_),
    .Q(\as2650.pc[13] ));
 sky130_fd_sc_hd__dfxtp_4 _6233_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0230_),
    .Q(\as2650.pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6234_ (.CLK(clknet_leaf_16_clk),
    .D(_0231_),
    .Q(\as2650.r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6235_ (.CLK(clknet_leaf_18_clk),
    .D(_0232_),
    .Q(\as2650.r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6236_ (.CLK(clknet_leaf_17_clk),
    .D(_0233_),
    .Q(\as2650.r0[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6237_ (.CLK(clknet_leaf_17_clk),
    .D(_0234_),
    .Q(\as2650.r0[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6238_ (.CLK(clknet_leaf_18_clk),
    .D(_0235_),
    .Q(\as2650.r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6239_ (.CLK(clknet_leaf_18_clk),
    .D(_0236_),
    .Q(\as2650.r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6240_ (.CLK(clknet_leaf_17_clk),
    .D(_0237_),
    .Q(\as2650.r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6241_ (.CLK(clknet_leaf_17_clk),
    .D(_0238_),
    .Q(\as2650.r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6242_ (.CLK(clknet_leaf_41_clk),
    .D(_0239_),
    .Q(\as2650.stack[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6243_ (.CLK(clknet_leaf_39_clk),
    .D(_0240_),
    .Q(\as2650.stack[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6244_ (.CLK(clknet_leaf_47_clk),
    .D(_0241_),
    .Q(\as2650.stack[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6245_ (.CLK(clknet_leaf_47_clk),
    .D(_0242_),
    .Q(\as2650.stack[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6246_ (.CLK(clknet_leaf_47_clk),
    .D(_0243_),
    .Q(\as2650.stack[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6247_ (.CLK(clknet_leaf_47_clk),
    .D(_0244_),
    .Q(\as2650.stack[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6248_ (.CLK(clknet_leaf_38_clk),
    .D(_0245_),
    .Q(\as2650.stack[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6249_ (.CLK(clknet_leaf_48_clk),
    .D(_0246_),
    .Q(\as2650.stack[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6250_ (.CLK(clknet_leaf_40_clk),
    .D(_0247_),
    .Q(\as2650.stack[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6251_ (.CLK(clknet_leaf_39_clk),
    .D(_0248_),
    .Q(\as2650.stack[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6252_ (.CLK(clknet_leaf_48_clk),
    .D(_0249_),
    .Q(\as2650.stack[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6253_ (.CLK(clknet_leaf_48_clk),
    .D(_0250_),
    .Q(\as2650.stack[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6254_ (.CLK(clknet_leaf_47_clk),
    .D(_0251_),
    .Q(\as2650.stack[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6255_ (.CLK(clknet_leaf_39_clk),
    .D(_0252_),
    .Q(\as2650.stack[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6256_ (.CLK(clknet_leaf_39_clk),
    .D(_0253_),
    .Q(\as2650.stack[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6257_ (.CLK(clknet_leaf_48_clk),
    .D(_0254_),
    .Q(\as2650.stack[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6258_ (.CLK(clknet_leaf_25_clk),
    .D(_0255_),
    .Q(\as2650.stack[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6259_ (.CLK(clknet_leaf_42_clk),
    .D(_0256_),
    .Q(\as2650.stack[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6260_ (.CLK(clknet_leaf_36_clk),
    .D(_0257_),
    .Q(\as2650.stack[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6261_ (.CLK(clknet_leaf_30_clk),
    .D(_0258_),
    .Q(\as2650.stack[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6262_ (.CLK(clknet_leaf_43_clk),
    .D(_0259_),
    .Q(\as2650.stack[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6263_ (.CLK(clknet_leaf_30_clk),
    .D(_0260_),
    .Q(\as2650.stack[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6264_ (.CLK(clknet_leaf_35_clk),
    .D(_0261_),
    .Q(\as2650.stack[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6265_ (.CLK(clknet_leaf_21_clk),
    .D(_0262_),
    .Q(\as2650.r123[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6266_ (.CLK(clknet_leaf_19_clk),
    .D(_0263_),
    .Q(\as2650.r123[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6267_ (.CLK(clknet_leaf_20_clk),
    .D(_0264_),
    .Q(\as2650.r123[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6268_ (.CLK(clknet_leaf_20_clk),
    .D(_0265_),
    .Q(\as2650.r123[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6269_ (.CLK(clknet_leaf_19_clk),
    .D(_0266_),
    .Q(\as2650.r123[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6270_ (.CLK(clknet_leaf_18_clk),
    .D(_0267_),
    .Q(\as2650.r123[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6271_ (.CLK(clknet_leaf_20_clk),
    .D(_0268_),
    .Q(\as2650.r123[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6272_ (.CLK(clknet_leaf_19_clk),
    .D(_0269_),
    .Q(\as2650.r123[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6273_ (.CLK(clknet_leaf_27_clk),
    .D(_0270_),
    .Q(\as2650.r123[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6274_ (.CLK(clknet_leaf_20_clk),
    .D(_0271_),
    .Q(\as2650.r123[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6275_ (.CLK(clknet_leaf_27_clk),
    .D(_0272_),
    .Q(\as2650.r123[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6276_ (.CLK(clknet_leaf_27_clk),
    .D(_0273_),
    .Q(\as2650.r123[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6277_ (.CLK(clknet_leaf_29_clk),
    .D(_0274_),
    .Q(\as2650.r123[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6278_ (.CLK(clknet_leaf_26_clk),
    .D(_0275_),
    .Q(\as2650.r123[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6279_ (.CLK(clknet_leaf_29_clk),
    .D(_0276_),
    .Q(\as2650.r123[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6280_ (.CLK(clknet_leaf_27_clk),
    .D(_0277_),
    .Q(\as2650.r123[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6281_ (.CLK(clknet_leaf_55_clk),
    .D(_0278_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _6282_ (.CLK(clknet_leaf_55_clk),
    .D(_0279_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _6283_ (.CLK(clknet_leaf_55_clk),
    .D(_0280_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _6284_ (.CLK(clknet_leaf_55_clk),
    .D(_0281_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _6285_ (.CLK(clknet_leaf_56_clk),
    .D(_0282_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _6286_ (.CLK(clknet_leaf_56_clk),
    .D(_0283_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _6287_ (.CLK(clknet_leaf_0_clk),
    .D(_0284_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _6288_ (.CLK(clknet_leaf_0_clk),
    .D(_0285_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _6289_ (.CLK(clknet_leaf_8_clk),
    .D(_0286_),
    .Q(\as2650.ins_reg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6290_ (.CLK(clknet_leaf_8_clk),
    .D(_0287_),
    .Q(\as2650.ins_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6291_ (.CLK(clknet_leaf_14_clk),
    .D(_0288_),
    .Q(\as2650.psl[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6292_ (.CLK(clknet_leaf_10_clk),
    .D(_0289_),
    .Q(\as2650.carry ));
 sky130_fd_sc_hd__dfxtp_4 _6293_ (.CLK(clknet_leaf_41_clk),
    .D(_0290_),
    .Q(\as2650.psu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6294_ (.CLK(clknet_leaf_44_clk),
    .D(_0291_),
    .Q(\as2650.psu[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6295_ (.CLK(clknet_leaf_44_clk),
    .D(_0292_),
    .Q(\as2650.psu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6296_ (.CLK(clknet_leaf_11_clk),
    .D(_0293_),
    .Q(\as2650.overflow ));
 sky130_fd_sc_hd__dfxtp_1 _6297_ (.CLK(clknet_leaf_11_clk),
    .D(_0294_),
    .Q(\as2650.psl[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6298_ (.CLK(clknet_leaf_10_clk),
    .D(_0295_),
    .Q(\as2650.psl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6299_ (.CLK(clknet_leaf_14_clk),
    .D(_0296_),
    .Q(\as2650.psl[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6300_ (.CLK(clknet_leaf_10_clk),
    .D(_0297_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _6301_ (.CLK(clknet_leaf_11_clk),
    .D(_0298_),
    .Q(\as2650.psu[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6302_ (.CLK(clknet_leaf_10_clk),
    .D(_0299_),
    .Q(\as2650.psu[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(_2678_),
    .X(net101));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(_0831_),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(_0831_),
    .X(net103));
 sky130_fd_sc_hd__buf_4 fanout104 (.A(_0815_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_0762_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(_0464_),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(_0464_),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(_0400_),
    .X(net109));
 sky130_fd_sc_hd__buf_12 fanout110 (.A(_0352_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_16 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_6 fanout113 (.A(_0307_),
    .X(net113));
 sky130_fd_sc_hd__buf_12 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(_2952_),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout118 (.A(_2897_),
    .X(net118));
 sky130_fd_sc_hd__buf_12 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_12 fanout120 (.A(_2887_),
    .X(net120));
 sky130_fd_sc_hd__buf_12 fanout121 (.A(_2880_),
    .X(net121));
 sky130_fd_sc_hd__buf_12 fanout122 (.A(_2858_),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(_2858_),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_6 fanout125 (.A(_2811_),
    .X(net125));
 sky130_fd_sc_hd__buf_6 fanout126 (.A(_2791_),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(_2774_),
    .X(net127));
 sky130_fd_sc_hd__buf_6 fanout128 (.A(_2759_),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(_2732_),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(_2731_),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(_2714_),
    .X(net131));
 sky130_fd_sc_hd__buf_12 fanout132 (.A(_2705_),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(_2705_),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(_2705_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_8 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_16 fanout137 (.A(net140),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(_2704_),
    .X(net140));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(_2699_),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(_2699_),
    .X(net142));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(_2698_),
    .X(net143));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_8 fanout145 (.A(_2697_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_16 fanout146 (.A(_2696_),
    .X(net146));
 sky130_fd_sc_hd__buf_8 fanout147 (.A(_2693_),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(_2692_),
    .X(net148));
 sky130_fd_sc_hd__buf_12 fanout149 (.A(net152),
    .X(net149));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(net152),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(_2691_),
    .X(net152));
 sky130_fd_sc_hd__buf_12 fanout153 (.A(_2690_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(_2690_),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(_2690_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(_2690_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_16 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_8 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_6 fanout159 (.A(_2671_),
    .X(net159));
 sky130_fd_sc_hd__buf_12 fanout160 (.A(_2670_),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(_2670_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_16 fanout162 (.A(_2498_),
    .X(net162));
 sky130_fd_sc_hd__buf_8 fanout163 (.A(_0737_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net167),
    .X(net164));
 sky130_fd_sc_hd__buf_6 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_2853_),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(_2852_),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(_2852_),
    .X(net170));
 sky130_fd_sc_hd__buf_6 fanout171 (.A(_2793_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 fanout172 (.A(_2677_),
    .X(net172));
 sky130_fd_sc_hd__buf_8 fanout173 (.A(_2664_),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(_0608_),
    .X(net175));
 sky130_fd_sc_hd__buf_6 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(_0605_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_16 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(_0460_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(_0396_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_16 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_8 fanout183 (.A(_0349_),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(_0304_),
    .X(net185));
 sky130_fd_sc_hd__buf_6 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_6 fanout187 (.A(_2949_),
    .X(net187));
 sky130_fd_sc_hd__buf_8 fanout188 (.A(_2893_),
    .X(net188));
 sky130_fd_sc_hd__buf_6 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout190 (.A(_2854_),
    .X(net190));
 sky130_fd_sc_hd__buf_6 fanout191 (.A(_2854_),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(_2854_),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout193 (.A(_2848_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(_2848_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_16 fanout195 (.A(_2847_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_2785_),
    .X(net197));
 sky130_fd_sc_hd__buf_8 fanout198 (.A(net200),
    .X(net198));
 sky130_fd_sc_hd__buf_8 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(_2761_),
    .X(net200));
 sky130_fd_sc_hd__buf_6 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_6 fanout202 (.A(_2760_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(_2750_),
    .X(net204));
 sky130_fd_sc_hd__buf_8 fanout205 (.A(_2749_),
    .X(net205));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(_2745_),
    .X(net206));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(_2675_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_16 fanout209 (.A(_2674_),
    .X(net209));
 sky130_fd_sc_hd__buf_6 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(_2665_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(_2646_),
    .X(net212));
 sky130_fd_sc_hd__buf_8 fanout213 (.A(_2646_),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(_2646_),
    .X(net214));
 sky130_fd_sc_hd__buf_12 fanout215 (.A(_2645_),
    .X(net215));
 sky130_fd_sc_hd__buf_6 fanout216 (.A(_2645_),
    .X(net216));
 sky130_fd_sc_hd__buf_6 fanout217 (.A(_2638_),
    .X(net217));
 sky130_fd_sc_hd__buf_8 fanout218 (.A(_2636_),
    .X(net218));
 sky130_fd_sc_hd__buf_8 fanout219 (.A(_2627_),
    .X(net219));
 sky130_fd_sc_hd__buf_8 fanout220 (.A(net222),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_16 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_6 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_8 fanout223 (.A(\as2650.psl[4] ),
    .X(net223));
 sky130_fd_sc_hd__buf_12 fanout224 (.A(\as2650.psu[0] ),
    .X(net224));
 sky130_fd_sc_hd__buf_8 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(\as2650.psu[1] ),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(\as2650.psu[2] ),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(\as2650.psu[2] ),
    .X(net228));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net232),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_16 fanout230 (.A(net232),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_6 fanout232 (.A(\as2650.ins_reg[4] ),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_16 fanout233 (.A(\as2650.ins_reg[4] ),
    .X(net233));
 sky130_fd_sc_hd__buf_6 fanout234 (.A(\as2650.ins_reg[4] ),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_6 fanout236 (.A(net238),
    .X(net236));
 sky130_fd_sc_hd__buf_12 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(\as2650.ins_reg[3] ),
    .X(net238));
 sky130_fd_sc_hd__buf_8 fanout239 (.A(net242),
    .X(net239));
 sky130_fd_sc_hd__buf_6 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_16 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_6 fanout242 (.A(\as2650.r0[7] ),
    .X(net242));
 sky130_fd_sc_hd__buf_8 fanout243 (.A(net246),
    .X(net243));
 sky130_fd_sc_hd__buf_8 fanout244 (.A(net246),
    .X(net244));
 sky130_fd_sc_hd__buf_6 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_16 fanout246 (.A(\as2650.r0[6] ),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(net250),
    .X(net247));
 sky130_fd_sc_hd__buf_8 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_12 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout250 (.A(\as2650.r0[5] ),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(\as2650.r0[4] ),
    .X(net251));
 sky130_fd_sc_hd__buf_8 fanout252 (.A(\as2650.r0[4] ),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(\as2650.r0[4] ),
    .X(net253));
 sky130_fd_sc_hd__buf_8 fanout254 (.A(\as2650.r0[3] ),
    .X(net254));
 sky130_fd_sc_hd__buf_8 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__buf_12 fanout256 (.A(\as2650.r0[3] ),
    .X(net256));
 sky130_fd_sc_hd__buf_6 fanout257 (.A(net260),
    .X(net257));
 sky130_fd_sc_hd__buf_8 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_12 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_6 fanout260 (.A(\as2650.r0[2] ),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout261 (.A(net264),
    .X(net261));
 sky130_fd_sc_hd__buf_6 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_6 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_12 fanout264 (.A(\as2650.r0[1] ),
    .X(net264));
 sky130_fd_sc_hd__buf_6 fanout265 (.A(net268),
    .X(net265));
 sky130_fd_sc_hd__buf_6 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_8 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(\as2650.r0[0] ),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(\as2650.pc[12] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(\as2650.pc[11] ),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_6 fanout272 (.A(\as2650.pc[10] ),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_16 fanout273 (.A(\as2650.pc[9] ),
    .X(net273));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(\as2650.pc[8] ),
    .X(net274));
 sky130_fd_sc_hd__buf_6 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 fanout276 (.A(\as2650.pc[7] ),
    .X(net276));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_16 fanout278 (.A(\as2650.pc[6] ),
    .X(net278));
 sky130_fd_sc_hd__buf_6 fanout279 (.A(\as2650.pc[5] ),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(\as2650.pc[5] ),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_16 fanout281 (.A(\as2650.pc[4] ),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(\as2650.pc[4] ),
    .X(net282));
 sky130_fd_sc_hd__buf_8 fanout283 (.A(\as2650.pc[3] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(\as2650.pc[1] ),
    .X(net284));
 sky130_fd_sc_hd__buf_6 fanout285 (.A(\as2650.pc[1] ),
    .X(net285));
 sky130_fd_sc_hd__buf_8 fanout286 (.A(net288),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(\as2650.pc[0] ),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(\as2650.cycle[3] ),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(\as2650.cycle[2] ),
    .X(net290));
 sky130_fd_sc_hd__buf_6 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_6 fanout292 (.A(\as2650.cycle[1] ),
    .X(net292));
 sky130_fd_sc_hd__buf_8 fanout293 (.A(\as2650.cycle[0] ),
    .X(net293));
 sky130_fd_sc_hd__buf_8 fanout294 (.A(net296),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(\as2650.halted ),
    .X(net296));
 sky130_fd_sc_hd__buf_12 fanout297 (.A(\as2650.ins_reg[7] ),
    .X(net297));
 sky130_fd_sc_hd__buf_12 fanout298 (.A(\as2650.ins_reg[6] ),
    .X(net298));
 sky130_fd_sc_hd__buf_12 fanout299 (.A(\as2650.ins_reg[5] ),
    .X(net299));
 sky130_fd_sc_hd__buf_8 fanout300 (.A(\as2650.ins_reg[5] ),
    .X(net300));
 sky130_fd_sc_hd__buf_6 fanout301 (.A(net303),
    .X(net301));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_12 fanout303 (.A(\as2650.ins_reg[2] ),
    .X(net303));
 sky130_fd_sc_hd__buf_12 fanout304 (.A(\as2650.ins_reg[1] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_8 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(\as2650.ins_reg[0] ),
    .X(net306));
 sky130_fd_sc_hd__buf_8 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__buf_6 fanout308 (.A(\as2650.ins_reg[0] ),
    .X(net308));
 sky130_fd_sc_hd__buf_12 fanout309 (.A(\as2650.addr_buff[7] ),
    .X(net309));
 sky130_fd_sc_hd__buf_6 fanout310 (.A(\as2650.addr_buff[0] ),
    .X(net310));
 sky130_fd_sc_hd__buf_6 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_8 fanout312 (.A(_2650_),
    .X(net312));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_4 fanout315 (.A(_2649_),
    .X(net315));
 sky130_fd_sc_hd__buf_6 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_6 fanout317 (.A(_2649_),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_8 fanout318 (.A(net321),
    .X(net318));
 sky130_fd_sc_hd__buf_4 fanout319 (.A(net321),
    .X(net319));
 sky130_fd_sc_hd__buf_6 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_8 fanout321 (.A(_2649_),
    .X(net321));
 sky130_fd_sc_hd__buf_8 fanout322 (.A(net9),
    .X(net322));
 sky130_fd_sc_hd__buf_2 fanout323 (.A(net9),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_6 fanout325 (.A(net9),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_6 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__buf_8 fanout328 (.A(net8),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_4 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__buf_6 fanout331 (.A(net8),
    .X(net331));
 sky130_fd_sc_hd__buf_8 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_6 fanout333 (.A(net335),
    .X(net333));
 sky130_fd_sc_hd__buf_8 fanout334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_16 fanout335 (.A(net7),
    .X(net335));
 sky130_fd_sc_hd__buf_6 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_12 fanout337 (.A(net6),
    .X(net337));
 sky130_fd_sc_hd__buf_6 fanout338 (.A(net5),
    .X(net338));
 sky130_fd_sc_hd__buf_12 fanout339 (.A(net5),
    .X(net339));
 sky130_fd_sc_hd__buf_6 fanout340 (.A(net4),
    .X(net340));
 sky130_fd_sc_hd__buf_12 fanout341 (.A(net4),
    .X(net341));
 sky130_fd_sc_hd__buf_8 fanout342 (.A(net3),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 fanout343 (.A(net3),
    .X(net343));
 sky130_fd_sc_hd__buf_8 fanout344 (.A(net3),
    .X(net344));
 sky130_fd_sc_hd__buf_8 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_12 fanout346 (.A(net2),
    .X(net346));
 sky130_fd_sc_hd__buf_6 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_6 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_16 fanout349 (.A(net1),
    .X(net349));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(_1380_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 fanout41 (.A(_0916_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_0916_),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_8 fanout44 (.A(_2497_),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(_1970_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(_1077_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(_1071_),
    .X(net48));
 sky130_fd_sc_hd__buf_6 fanout49 (.A(_0584_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(_1073_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(_0908_),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(_1409_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(_0624_),
    .X(net54));
 sky130_fd_sc_hd__buf_8 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_16 fanout56 (.A(_0588_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_2816_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(_2797_),
    .X(net58));
 sky130_fd_sc_hd__buf_6 fanout59 (.A(_0824_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(_0636_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_2866_),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(_2866_),
    .X(net62));
 sky130_fd_sc_hd__buf_6 fanout63 (.A(_1397_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(_1393_),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(_1356_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(_1356_),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 fanout69 (.A(_1355_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(_0749_),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(_0748_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 fanout72 (.A(_0580_),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_2808_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(_2808_),
    .X(net74));
 sky130_fd_sc_hd__buf_4 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(_2807_),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(_2742_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 fanout78 (.A(_2736_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(_2736_),
    .X(net79));
 sky130_fd_sc_hd__buf_6 fanout80 (.A(_2724_),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout81 (.A(_2723_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(_2723_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_16 fanout84 (.A(_2712_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_16 fanout85 (.A(_2711_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(_2711_),
    .X(net86));
 sky130_fd_sc_hd__buf_6 fanout87 (.A(net89),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(_2701_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_8 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__buf_12 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(_2700_),
    .X(net94));
 sky130_fd_sc_hd__buf_6 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(_2700_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 fanout97 (.A(_2679_),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(_2679_),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_8 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_8 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input9 (.A(rst),
    .X(net9));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output17 (.A(net17),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 output36 (.A(net36),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_4 output37 (.A(net37),
    .X(io_out[9]));
endmodule

