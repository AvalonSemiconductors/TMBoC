VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO posit_unit
  CLASS BLOCK ;
  FOREIGN posit_unit ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.820 4.000 175.020 ;
    END
  END io_in[2]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 0.000 44.210 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.050 0.000 131.610 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.450 0.000 219.010 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 0.000 306.410 4.000 ;
    END
  END io_out[3]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.540 4.000 313.740 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 344.080 337.520 ;
      LAYER met2 ;
        RECT 7.000 4.280 341.680 337.465 ;
        RECT 7.000 4.000 43.370 4.280 ;
        RECT 44.490 4.000 130.770 4.280 ;
        RECT 131.890 4.000 218.170 4.280 ;
        RECT 219.290 4.000 305.570 4.280 ;
        RECT 306.690 4.000 341.680 4.280 ;
      LAYER met3 ;
        RECT 4.000 314.140 329.830 337.445 ;
        RECT 4.400 312.140 329.830 314.140 ;
        RECT 4.000 244.780 329.830 312.140 ;
        RECT 4.400 242.780 329.830 244.780 ;
        RECT 4.000 175.420 329.830 242.780 ;
        RECT 4.400 173.420 329.830 175.420 ;
        RECT 4.000 106.060 329.830 173.420 ;
        RECT 4.400 104.060 329.830 106.060 ;
        RECT 4.000 36.700 329.830 104.060 ;
        RECT 4.400 34.700 329.830 36.700 ;
        RECT 4.000 10.715 329.830 34.700 ;
      LAYER met4 ;
        RECT 15.935 17.175 20.640 290.185 ;
        RECT 23.040 17.175 97.440 290.185 ;
        RECT 99.840 17.175 174.240 290.185 ;
        RECT 176.640 17.175 251.040 290.185 ;
        RECT 253.440 17.175 289.505 290.185 ;
  END
END posit_unit
END LIBRARY

