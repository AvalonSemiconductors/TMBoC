magic
tech sky130B
magscale 1 2
timestamp 1684334855
<< obsli1 >>
rect 1104 2159 10856 15793
<< obsm1 >>
rect 566 2128 11394 15824
<< metal2 >>
rect 2962 17200 3018 18000
rect 8942 17200 8998 18000
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
rect 11334 0 11390 800
<< obsm2 >>
rect 572 17144 2906 17200
rect 3074 17144 8886 17200
rect 9054 17144 11388 17200
rect 572 856 11388 17144
rect 682 800 1710 856
rect 1878 800 2906 856
rect 3074 800 4102 856
rect 4270 800 5298 856
rect 5466 800 6494 856
rect 6662 800 7690 856
rect 7858 800 8886 856
rect 9054 800 10082 856
rect 10250 800 11278 856
<< metal3 >>
rect 11200 15920 12000 16040
rect 11200 12384 12000 12504
rect 11200 8848 12000 8968
rect 11200 5312 12000 5432
rect 11200 1776 12000 1896
<< obsm3 >>
rect 2165 15840 11120 16013
rect 2165 12584 11346 15840
rect 2165 12304 11120 12584
rect 2165 9048 11346 12304
rect 2165 8768 11120 9048
rect 2165 5512 11346 8768
rect 2165 5232 11120 5512
rect 2165 1976 11346 5232
rect 2165 1803 11120 1976
<< metal4 >>
rect 2163 2128 2483 15824
rect 3382 2128 3702 15824
rect 4601 2128 4921 15824
rect 5820 2128 6140 15824
rect 7039 2128 7359 15824
rect 8258 2128 8578 15824
rect 9477 2128 9797 15824
rect 10696 2128 11016 15824
<< labels >>
rlabel metal2 s 2962 17200 3018 18000 6 clk
port 1 nsew signal input
rlabel metal3 s 11200 1776 12000 1896 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 11200 5312 12000 5432 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 11200 8848 12000 8968 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 11200 12384 12000 12504 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 11200 15920 12000 16040 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 io_oeb
port 7 nsew signal output
rlabel metal2 s 570 0 626 800 6 io_out[0]
port 8 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 io_out[1]
port 9 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 io_out[2]
port 10 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 io_out[3]
port 11 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 io_out[4]
port 12 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 io_out[5]
port 13 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 io_out[6]
port 14 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 io_out[8]
port 16 nsew signal output
rlabel metal2 s 8942 17200 8998 18000 6 rst
port 17 nsew signal input
rlabel metal4 s 2163 2128 2483 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 15824 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 3382 2128 3702 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 5820 2128 6140 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 8258 2128 8578 15824 6 vssd1
port 19 nsew ground bidirectional
rlabel metal4 s 10696 2128 11016 15824 6 vssd1
port 19 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 466022
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MC14500/runs/23_05_17_16_45/results/signoff/wrapped_MC14500.magic.gds
string GDS_START 205780
<< end >>

