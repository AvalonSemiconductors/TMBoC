magic
tech sky130B
magscale 1 2
timestamp 1680008481
<< nwell >>
rect 1066 41605 43922 42171
rect 1066 40517 43922 41083
rect 1066 39429 43922 39995
rect 1066 38341 43922 38907
rect 1066 37253 43922 37819
rect 1066 36165 43922 36731
rect 1066 35077 43922 35643
rect 1066 33989 43922 34555
rect 1066 32901 43922 33467
rect 1066 31813 43922 32379
rect 1066 30725 43922 31291
rect 1066 29637 43922 30203
rect 1066 28549 43922 29115
rect 1066 27461 43922 28027
rect 1066 26373 43922 26939
rect 1066 25285 43922 25851
rect 1066 24197 43922 24763
rect 1066 23109 43922 23675
rect 1066 22021 43922 22587
rect 1066 20933 43922 21499
rect 1066 19845 43922 20411
rect 1066 18757 43922 19323
rect 1066 17669 43922 18235
rect 1066 16581 43922 17147
rect 1066 15493 43922 16059
rect 1066 14405 43922 14971
rect 1066 13317 43922 13883
rect 1066 12229 43922 12795
rect 1066 11141 43922 11707
rect 1066 10053 43922 10619
rect 1066 8965 43922 9531
rect 1066 7877 43922 8443
rect 1066 6789 43922 7355
rect 1066 5701 43922 6267
rect 1066 4613 43922 5179
rect 1066 3525 43922 4091
rect 1066 2437 43922 3003
<< obsli1 >>
rect 1104 2159 43884 42449
<< obsm1 >>
rect 1104 2128 44054 44124
<< metal2 >>
rect 2226 44200 2282 45000
rect 5906 44200 5962 45000
rect 9586 44200 9642 45000
rect 13266 44200 13322 45000
rect 16946 44200 17002 45000
rect 20626 44200 20682 45000
rect 24306 44200 24362 45000
rect 27986 44200 28042 45000
rect 31666 44200 31722 45000
rect 35346 44200 35402 45000
rect 39026 44200 39082 45000
rect 42706 44200 42762 45000
<< obsm2 >>
rect 2338 44144 5850 44200
rect 6018 44144 9530 44200
rect 9698 44144 13210 44200
rect 13378 44144 16890 44200
rect 17058 44144 20570 44200
rect 20738 44144 24250 44200
rect 24418 44144 27930 44200
rect 28098 44144 31610 44200
rect 31778 44144 35290 44200
rect 35458 44144 38970 44200
rect 39138 44144 42650 44200
rect 42818 44144 44050 44200
rect 2228 2139 44050 44144
<< metal3 >>
rect 44200 42576 45000 42696
rect 44200 41080 45000 41200
rect 44200 39584 45000 39704
rect 44200 38088 45000 38208
rect 44200 36592 45000 36712
rect 44200 35096 45000 35216
rect 44200 33600 45000 33720
rect 44200 32104 45000 32224
rect 44200 30608 45000 30728
rect 44200 29112 45000 29232
rect 44200 27616 45000 27736
rect 44200 26120 45000 26240
rect 44200 24624 45000 24744
rect 44200 23128 45000 23248
rect 44200 21632 45000 21752
rect 44200 20136 45000 20256
rect 44200 18640 45000 18760
rect 44200 17144 45000 17264
rect 44200 15648 45000 15768
rect 44200 14152 45000 14272
rect 44200 12656 45000 12776
rect 44200 11160 45000 11280
rect 44200 9664 45000 9784
rect 44200 8168 45000 8288
rect 44200 6672 45000 6792
rect 44200 5176 45000 5296
rect 44200 3680 45000 3800
rect 44200 2184 45000 2304
<< obsm3 >>
rect 4210 42496 44120 42669
rect 4210 41280 44200 42496
rect 4210 41000 44120 41280
rect 4210 39784 44200 41000
rect 4210 39504 44120 39784
rect 4210 38288 44200 39504
rect 4210 38008 44120 38288
rect 4210 36792 44200 38008
rect 4210 36512 44120 36792
rect 4210 35296 44200 36512
rect 4210 35016 44120 35296
rect 4210 33800 44200 35016
rect 4210 33520 44120 33800
rect 4210 32304 44200 33520
rect 4210 32024 44120 32304
rect 4210 30808 44200 32024
rect 4210 30528 44120 30808
rect 4210 29312 44200 30528
rect 4210 29032 44120 29312
rect 4210 27816 44200 29032
rect 4210 27536 44120 27816
rect 4210 26320 44200 27536
rect 4210 26040 44120 26320
rect 4210 24824 44200 26040
rect 4210 24544 44120 24824
rect 4210 23328 44200 24544
rect 4210 23048 44120 23328
rect 4210 21832 44200 23048
rect 4210 21552 44120 21832
rect 4210 20336 44200 21552
rect 4210 20056 44120 20336
rect 4210 18840 44200 20056
rect 4210 18560 44120 18840
rect 4210 17344 44200 18560
rect 4210 17064 44120 17344
rect 4210 15848 44200 17064
rect 4210 15568 44120 15848
rect 4210 14352 44200 15568
rect 4210 14072 44120 14352
rect 4210 12856 44200 14072
rect 4210 12576 44120 12856
rect 4210 11360 44200 12576
rect 4210 11080 44120 11360
rect 4210 9864 44200 11080
rect 4210 9584 44120 9864
rect 4210 8368 44200 9584
rect 4210 8088 44120 8368
rect 4210 6872 44200 8088
rect 4210 6592 44120 6872
rect 4210 5376 44200 6592
rect 4210 5096 44120 5376
rect 4210 3880 44200 5096
rect 4210 3600 44120 3880
rect 4210 2384 44200 3600
rect 4210 2143 44120 2384
<< metal4 >>
rect 4208 2128 4528 42480
rect 19568 2128 19888 42480
rect 34928 2128 35248 42480
<< obsm4 >>
rect 8155 17851 19488 41445
rect 19968 17851 34848 41445
rect 35328 17851 39133 41445
<< labels >>
rlabel metal2 s 39026 44200 39082 45000 6 clk
port 1 nsew signal input
rlabel metal2 s 2226 44200 2282 45000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 5906 44200 5962 45000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 9586 44200 9642 45000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 13266 44200 13322 45000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 16946 44200 17002 45000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 20626 44200 20682 45000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 24306 44200 24362 45000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 27986 44200 28042 45000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 31666 44200 31722 45000 6 io_in[8]
port 10 nsew signal input
rlabel metal2 s 35346 44200 35402 45000 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 44200 42576 45000 42696 6 io_oeb
port 12 nsew signal output
rlabel metal3 s 44200 2184 45000 2304 6 io_out[0]
port 13 nsew signal output
rlabel metal3 s 44200 17144 45000 17264 6 io_out[10]
port 14 nsew signal output
rlabel metal3 s 44200 18640 45000 18760 6 io_out[11]
port 15 nsew signal output
rlabel metal3 s 44200 20136 45000 20256 6 io_out[12]
port 16 nsew signal output
rlabel metal3 s 44200 21632 45000 21752 6 io_out[13]
port 17 nsew signal output
rlabel metal3 s 44200 23128 45000 23248 6 io_out[14]
port 18 nsew signal output
rlabel metal3 s 44200 24624 45000 24744 6 io_out[15]
port 19 nsew signal output
rlabel metal3 s 44200 26120 45000 26240 6 io_out[16]
port 20 nsew signal output
rlabel metal3 s 44200 27616 45000 27736 6 io_out[17]
port 21 nsew signal output
rlabel metal3 s 44200 29112 45000 29232 6 io_out[18]
port 22 nsew signal output
rlabel metal3 s 44200 30608 45000 30728 6 io_out[19]
port 23 nsew signal output
rlabel metal3 s 44200 3680 45000 3800 6 io_out[1]
port 24 nsew signal output
rlabel metal3 s 44200 32104 45000 32224 6 io_out[20]
port 25 nsew signal output
rlabel metal3 s 44200 33600 45000 33720 6 io_out[21]
port 26 nsew signal output
rlabel metal3 s 44200 35096 45000 35216 6 io_out[22]
port 27 nsew signal output
rlabel metal3 s 44200 36592 45000 36712 6 io_out[23]
port 28 nsew signal output
rlabel metal3 s 44200 38088 45000 38208 6 io_out[24]
port 29 nsew signal output
rlabel metal3 s 44200 39584 45000 39704 6 io_out[25]
port 30 nsew signal output
rlabel metal3 s 44200 41080 45000 41200 6 io_out[26]
port 31 nsew signal output
rlabel metal3 s 44200 5176 45000 5296 6 io_out[2]
port 32 nsew signal output
rlabel metal3 s 44200 6672 45000 6792 6 io_out[3]
port 33 nsew signal output
rlabel metal3 s 44200 8168 45000 8288 6 io_out[4]
port 34 nsew signal output
rlabel metal3 s 44200 9664 45000 9784 6 io_out[5]
port 35 nsew signal output
rlabel metal3 s 44200 11160 45000 11280 6 io_out[6]
port 36 nsew signal output
rlabel metal3 s 44200 12656 45000 12776 6 io_out[7]
port 37 nsew signal output
rlabel metal3 s 44200 14152 45000 14272 6 io_out[8]
port 38 nsew signal output
rlabel metal3 s 44200 15648 45000 15768 6 io_out[9]
port 39 nsew signal output
rlabel metal2 s 42706 44200 42762 45000 6 rst
port 40 nsew signal input
rlabel metal4 s 4208 2128 4528 42480 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 42480 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 42480 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4219484
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MOS6502/runs/23_03_28_14_58/results/signoff/wrapped_6502.magic.gds
string GDS_START 1065482
<< end >>

