module bitmap(
	input [14:0] addr,
	output val
);

reg [3:0] res;

assign val = res >> addr[1:0];

always @(*) begin
case(addr[14:2])
	0: res <= 0;
	1: res <= 0;
	2: res <= 0;
	3: res <= 0;
	4: res <= 0;
	5: res <= 0;
	6: res <= 0;
	7: res <= 0;
	8: res <= 0;
	9: res <= 0;
	10: res <= 0;
	11: res <= 0;
	12: res <= 0;
	13: res <= 0;
	14: res <= 0;
	15: res <= 0;
	16: res <= 0;
	17: res <= 0;
	18: res <= 0;
	19: res <= 0;
	20: res <= 0;
	21: res <= 0;
	22: res <= 0;
	23: res <= 0;
	24: res <= 0;
	25: res <= 0;
	26: res <= 0;
	27: res <= 0;
	28: res <= 0;
	29: res <= 0;
	30: res <= 0;
	31: res <= 0;
	32: res <= 0;
	33: res <= 0;
	34: res <= 0;
	35: res <= 0;
	36: res <= 0;
	37: res <= 0;
	38: res <= 0;
	39: res <= 0;
	40: res <= 0;
	41: res <= 0;
	42: res <= 0;
	43: res <= 0;
	44: res <= 0;
	45: res <= 0;
	46: res <= 0;
	47: res <= 0;
	48: res <= 0;
	49: res <= 0;
	50: res <= 0;
	51: res <= 0;
	52: res <= 0;
	53: res <= 0;
	54: res <= 0;
	55: res <= 0;
	56: res <= 0;
	57: res <= 0;
	58: res <= 0;
	59: res <= 0;
	60: res <= 0;
	61: res <= 0;
	62: res <= 0;
	63: res <= 0;
	64: res <= 0;
	65: res <= 0;
	66: res <= 0;
	67: res <= 0;
	68: res <= 0;
	69: res <= 0;
	70: res <= 0;
	71: res <= 0;
	72: res <= 0;
	73: res <= 0;
	74: res <= 0;
	75: res <= 0;
	76: res <= 0;
	77: res <= 0;
	78: res <= 0;
	79: res <= 0;
	80: res <= 0;
	81: res <= 0;
	82: res <= 0;
	83: res <= 0;
	84: res <= 0;
	85: res <= 0;
	86: res <= 0;
	87: res <= 0;
	88: res <= 0;
	89: res <= 0;
	90: res <= 0;
	91: res <= 0;
	92: res <= 0;
	93: res <= 0;
	94: res <= 0;
	95: res <= 0;
	96: res <= 0;
	97: res <= 0;
	98: res <= 0;
	99: res <= 0;
	100: res <= 0;
	101: res <= 0;
	102: res <= 0;
	103: res <= 0;
	104: res <= 0;
	105: res <= 0;
	106: res <= 0;
	107: res <= 0;
	108: res <= 0;
	109: res <= 0;
	110: res <= 0;
	111: res <= 0;
	112: res <= 0;
	113: res <= 0;
	114: res <= 0;
	115: res <= 0;
	116: res <= 0;
	117: res <= 0;
	118: res <= 0;
	119: res <= 0;
	120: res <= 0;
	121: res <= 0;
	122: res <= 0;
	123: res <= 0;
	124: res <= 0;
	125: res <= 0;
	126: res <= 0;
	127: res <= 0;
	128: res <= 0;
	129: res <= 0;
	130: res <= 0;
	131: res <= 0;
	132: res <= 0;
	133: res <= 0;
	134: res <= 0;
	135: res <= 0;
	136: res <= 7;
	137: res <= 0;
	138: res <= 0;
	139: res <= 7;
	140: res <= 8;
	141: res <= 15;
	142: res <= 15;
	143: res <= 0;
	144: res <= 8;
	145: res <= 3;
	146: res <= 0;
	147: res <= 8;
	148: res <= 3;
	149: res <= 0;
	150: res <= 0;
	151: res <= 0;
	152: res <= 0;
	153: res <= 12;
	154: res <= 15;
	155: res <= 0;
	156: res <= 0;
	157: res <= 0;
	158: res <= 0;
	159: res <= 0;
	160: res <= 0;
	161: res <= 0;
	162: res <= 0;
	163: res <= 0;
	164: res <= 0;
	165: res <= 0;
	166: res <= 0;
	167: res <= 0;
	168: res <= 0;
	169: res <= 0;
	170: res <= 0;
	171: res <= 0;
	172: res <= 0;
	173: res <= 0;
	174: res <= 0;
	175: res <= 0;
	176: res <= 0;
	177: res <= 0;
	178: res <= 0;
	179: res <= 0;
	180: res <= 0;
	181: res <= 7;
	182: res <= 0;
	183: res <= 0;
	184: res <= 7;
	185: res <= 8;
	186: res <= 15;
	187: res <= 15;
	188: res <= 0;
	189: res <= 8;
	190: res <= 3;
	191: res <= 0;
	192: res <= 8;
	193: res <= 3;
	194: res <= 0;
	195: res <= 0;
	196: res <= 0;
	197: res <= 0;
	198: res <= 12;
	199: res <= 15;
	200: res <= 0;
	201: res <= 0;
	202: res <= 0;
	203: res <= 0;
	204: res <= 0;
	205: res <= 0;
	206: res <= 0;
	207: res <= 0;
	208: res <= 6;
	209: res <= 0;
	210: res <= 0;
	211: res <= 0;
	212: res <= 0;
	213: res <= 0;
	214: res <= 0;
	215: res <= 0;
	216: res <= 0;
	217: res <= 0;
	218: res <= 0;
	219: res <= 0;
	220: res <= 0;
	221: res <= 0;
	222: res <= 0;
	223: res <= 0;
	224: res <= 0;
	225: res <= 0;
	226: res <= 7;
	227: res <= 0;
	228: res <= 0;
	229: res <= 7;
	230: res <= 8;
	231: res <= 15;
	232: res <= 15;
	233: res <= 0;
	234: res <= 8;
	235: res <= 3;
	236: res <= 0;
	237: res <= 8;
	238: res <= 3;
	239: res <= 0;
	240: res <= 0;
	241: res <= 0;
	242: res <= 0;
	243: res <= 12;
	244: res <= 15;
	245: res <= 0;
	246: res <= 0;
	247: res <= 0;
	248: res <= 0;
	249: res <= 0;
	250: res <= 0;
	251: res <= 0;
	252: res <= 0;
	253: res <= 6;
	254: res <= 0;
	255: res <= 0;
	256: res <= 0;
	257: res <= 0;
	258: res <= 0;
	259: res <= 0;
	260: res <= 0;
	261: res <= 15;
	262: res <= 15;
	263: res <= 15;
	264: res <= 7;
	265: res <= 0;
	266: res <= 0;
	267: res <= 0;
	268: res <= 0;
	269: res <= 0;
	270: res <= 0;
	271: res <= 15;
	272: res <= 3;
	273: res <= 14;
	274: res <= 7;
	275: res <= 8;
	276: res <= 3;
	277: res <= 0;
	278: res <= 7;
	279: res <= 8;
	280: res <= 3;
	281: res <= 0;
	282: res <= 8;
	283: res <= 3;
	284: res <= 0;
	285: res <= 0;
	286: res <= 0;
	287: res <= 8;
	288: res <= 3;
	289: res <= 0;
	290: res <= 7;
	291: res <= 0;
	292: res <= 0;
	293: res <= 0;
	294: res <= 0;
	295: res <= 0;
	296: res <= 0;
	297: res <= 0;
	298: res <= 15;
	299: res <= 0;
	300: res <= 0;
	301: res <= 0;
	302: res <= 0;
	303: res <= 0;
	304: res <= 0;
	305: res <= 0;
	306: res <= 15;
	307: res <= 15;
	308: res <= 15;
	309: res <= 7;
	310: res <= 0;
	311: res <= 0;
	312: res <= 0;
	313: res <= 0;
	314: res <= 0;
	315: res <= 0;
	316: res <= 15;
	317: res <= 3;
	318: res <= 14;
	319: res <= 7;
	320: res <= 8;
	321: res <= 3;
	322: res <= 0;
	323: res <= 7;
	324: res <= 8;
	325: res <= 3;
	326: res <= 0;
	327: res <= 8;
	328: res <= 3;
	329: res <= 0;
	330: res <= 0;
	331: res <= 0;
	332: res <= 8;
	333: res <= 3;
	334: res <= 0;
	335: res <= 7;
	336: res <= 0;
	337: res <= 0;
	338: res <= 0;
	339: res <= 0;
	340: res <= 0;
	341: res <= 0;
	342: res <= 8;
	343: res <= 15;
	344: res <= 0;
	345: res <= 0;
	346: res <= 0;
	347: res <= 0;
	348: res <= 0;
	349: res <= 0;
	350: res <= 0;
	351: res <= 15;
	352: res <= 15;
	353: res <= 15;
	354: res <= 7;
	355: res <= 0;
	356: res <= 0;
	357: res <= 0;
	358: res <= 0;
	359: res <= 0;
	360: res <= 0;
	361: res <= 15;
	362: res <= 15;
	363: res <= 15;
	364: res <= 7;
	365: res <= 8;
	366: res <= 3;
	367: res <= 0;
	368: res <= 7;
	369: res <= 8;
	370: res <= 3;
	371: res <= 0;
	372: res <= 8;
	373: res <= 3;
	374: res <= 0;
	375: res <= 0;
	376: res <= 0;
	377: res <= 8;
	378: res <= 3;
	379: res <= 0;
	380: res <= 7;
	381: res <= 0;
	382: res <= 0;
	383: res <= 0;
	384: res <= 0;
	385: res <= 0;
	386: res <= 0;
	387: res <= 12;
	388: res <= 15;
	389: res <= 0;
	390: res <= 0;
	391: res <= 0;
	392: res <= 0;
	393: res <= 0;
	394: res <= 0;
	395: res <= 0;
	396: res <= 0;
	397: res <= 12;
	398: res <= 1;
	399: res <= 0;
	400: res <= 0;
	401: res <= 0;
	402: res <= 0;
	403: res <= 0;
	404: res <= 0;
	405: res <= 0;
	406: res <= 7;
	407: res <= 12;
	408: res <= 1;
	409: res <= 7;
	410: res <= 8;
	411: res <= 15;
	412: res <= 15;
	413: res <= 0;
	414: res <= 8;
	415: res <= 3;
	416: res <= 0;
	417: res <= 8;
	418: res <= 3;
	419: res <= 0;
	420: res <= 0;
	421: res <= 0;
	422: res <= 8;
	423: res <= 3;
	424: res <= 0;
	425: res <= 7;
	426: res <= 0;
	427: res <= 0;
	428: res <= 0;
	429: res <= 0;
	430: res <= 0;
	431: res <= 0;
	432: res <= 12;
	433: res <= 15;
	434: res <= 1;
	435: res <= 0;
	436: res <= 0;
	437: res <= 0;
	438: res <= 0;
	439: res <= 0;
	440: res <= 0;
	441: res <= 0;
	442: res <= 12;
	443: res <= 1;
	444: res <= 0;
	445: res <= 0;
	446: res <= 0;
	447: res <= 0;
	448: res <= 0;
	449: res <= 0;
	450: res <= 0;
	451: res <= 7;
	452: res <= 12;
	453: res <= 1;
	454: res <= 7;
	455: res <= 8;
	456: res <= 15;
	457: res <= 15;
	458: res <= 0;
	459: res <= 8;
	460: res <= 3;
	461: res <= 0;
	462: res <= 8;
	463: res <= 3;
	464: res <= 12;
	465: res <= 15;
	466: res <= 7;
	467: res <= 8;
	468: res <= 3;
	469: res <= 0;
	470: res <= 7;
	471: res <= 0;
	472: res <= 0;
	473: res <= 0;
	474: res <= 0;
	475: res <= 0;
	476: res <= 0;
	477: res <= 14;
	478: res <= 15;
	479: res <= 1;
	480: res <= 0;
	481: res <= 0;
	482: res <= 0;
	483: res <= 0;
	484: res <= 0;
	485: res <= 0;
	486: res <= 0;
	487: res <= 12;
	488: res <= 1;
	489: res <= 0;
	490: res <= 0;
	491: res <= 0;
	492: res <= 0;
	493: res <= 0;
	494: res <= 0;
	495: res <= 0;
	496: res <= 7;
	497: res <= 0;
	498: res <= 0;
	499: res <= 7;
	500: res <= 8;
	501: res <= 15;
	502: res <= 15;
	503: res <= 0;
	504: res <= 8;
	505: res <= 3;
	506: res <= 14;
	507: res <= 8;
	508: res <= 3;
	509: res <= 12;
	510: res <= 15;
	511: res <= 7;
	512: res <= 8;
	513: res <= 3;
	514: res <= 0;
	515: res <= 7;
	516: res <= 0;
	517: res <= 0;
	518: res <= 0;
	519: res <= 0;
	520: res <= 0;
	521: res <= 0;
	522: res <= 15;
	523: res <= 15;
	524: res <= 1;
	525: res <= 0;
	526: res <= 0;
	527: res <= 0;
	528: res <= 0;
	529: res <= 0;
	530: res <= 0;
	531: res <= 0;
	532: res <= 12;
	533: res <= 1;
	534: res <= 0;
	535: res <= 0;
	536: res <= 0;
	537: res <= 0;
	538: res <= 0;
	539: res <= 0;
	540: res <= 0;
	541: res <= 7;
	542: res <= 0;
	543: res <= 0;
	544: res <= 7;
	545: res <= 8;
	546: res <= 3;
	547: res <= 0;
	548: res <= 0;
	549: res <= 8;
	550: res <= 3;
	551: res <= 14;
	552: res <= 8;
	553: res <= 3;
	554: res <= 12;
	555: res <= 15;
	556: res <= 7;
	557: res <= 0;
	558: res <= 12;
	559: res <= 15;
	560: res <= 7;
	561: res <= 0;
	562: res <= 0;
	563: res <= 0;
	564: res <= 0;
	565: res <= 0;
	566: res <= 8;
	567: res <= 15;
	568: res <= 15;
	569: res <= 1;
	570: res <= 0;
	571: res <= 0;
	572: res <= 0;
	573: res <= 0;
	574: res <= 0;
	575: res <= 0;
	576: res <= 0;
	577: res <= 12;
	578: res <= 1;
	579: res <= 0;
	580: res <= 0;
	581: res <= 0;
	582: res <= 0;
	583: res <= 0;
	584: res <= 0;
	585: res <= 0;
	586: res <= 7;
	587: res <= 0;
	588: res <= 0;
	589: res <= 7;
	590: res <= 8;
	591: res <= 3;
	592: res <= 0;
	593: res <= 0;
	594: res <= 8;
	595: res <= 3;
	596: res <= 14;
	597: res <= 8;
	598: res <= 3;
	599: res <= 0;
	600: res <= 0;
	601: res <= 0;
	602: res <= 0;
	603: res <= 12;
	604: res <= 15;
	605: res <= 7;
	606: res <= 0;
	607: res <= 0;
	608: res <= 0;
	609: res <= 0;
	610: res <= 0;
	611: res <= 12;
	612: res <= 15;
	613: res <= 15;
	614: res <= 1;
	615: res <= 0;
	616: res <= 0;
	617: res <= 0;
	618: res <= 0;
	619: res <= 0;
	620: res <= 0;
	621: res <= 0;
	622: res <= 12;
	623: res <= 1;
	624: res <= 0;
	625: res <= 0;
	626: res <= 0;
	627: res <= 0;
	628: res <= 0;
	629: res <= 0;
	630: res <= 0;
	631: res <= 7;
	632: res <= 0;
	633: res <= 0;
	634: res <= 7;
	635: res <= 8;
	636: res <= 3;
	637: res <= 0;
	638: res <= 0;
	639: res <= 8;
	640: res <= 15;
	641: res <= 1;
	642: res <= 15;
	643: res <= 3;
	644: res <= 0;
	645: res <= 0;
	646: res <= 0;
	647: res <= 0;
	648: res <= 12;
	649: res <= 15;
	650: res <= 7;
	651: res <= 0;
	652: res <= 0;
	653: res <= 0;
	654: res <= 0;
	655: res <= 0;
	656: res <= 12;
	657: res <= 15;
	658: res <= 15;
	659: res <= 1;
	660: res <= 0;
	661: res <= 0;
	662: res <= 0;
	663: res <= 0;
	664: res <= 0;
	665: res <= 0;
	666: res <= 0;
	667: res <= 12;
	668: res <= 1;
	669: res <= 0;
	670: res <= 0;
	671: res <= 0;
	672: res <= 0;
	673: res <= 0;
	674: res <= 0;
	675: res <= 0;
	676: res <= 7;
	677: res <= 0;
	678: res <= 0;
	679: res <= 7;
	680: res <= 8;
	681: res <= 3;
	682: res <= 0;
	683: res <= 0;
	684: res <= 8;
	685: res <= 15;
	686: res <= 1;
	687: res <= 15;
	688: res <= 3;
	689: res <= 0;
	690: res <= 0;
	691: res <= 0;
	692: res <= 0;
	693: res <= 0;
	694: res <= 0;
	695: res <= 7;
	696: res <= 0;
	697: res <= 0;
	698: res <= 0;
	699: res <= 0;
	700: res <= 0;
	701: res <= 14;
	702: res <= 15;
	703: res <= 15;
	704: res <= 1;
	705: res <= 0;
	706: res <= 0;
	707: res <= 0;
	708: res <= 0;
	709: res <= 0;
	710: res <= 0;
	711: res <= 0;
	712: res <= 12;
	713: res <= 1;
	714: res <= 0;
	715: res <= 0;
	716: res <= 0;
	717: res <= 0;
	718: res <= 0;
	719: res <= 0;
	720: res <= 0;
	721: res <= 7;
	722: res <= 0;
	723: res <= 0;
	724: res <= 7;
	725: res <= 8;
	726: res <= 3;
	727: res <= 0;
	728: res <= 0;
	729: res <= 8;
	730: res <= 15;
	731: res <= 1;
	732: res <= 15;
	733: res <= 3;
	734: res <= 0;
	735: res <= 0;
	736: res <= 0;
	737: res <= 0;
	738: res <= 0;
	739: res <= 0;
	740: res <= 7;
	741: res <= 0;
	742: res <= 0;
	743: res <= 0;
	744: res <= 0;
	745: res <= 0;
	746: res <= 15;
	747: res <= 15;
	748: res <= 15;
	749: res <= 1;
	750: res <= 0;
	751: res <= 0;
	752: res <= 0;
	753: res <= 0;
	754: res <= 0;
	755: res <= 0;
	756: res <= 0;
	757: res <= 12;
	758: res <= 1;
	759: res <= 0;
	760: res <= 0;
	761: res <= 0;
	762: res <= 0;
	763: res <= 0;
	764: res <= 0;
	765: res <= 0;
	766: res <= 7;
	767: res <= 0;
	768: res <= 0;
	769: res <= 7;
	770: res <= 8;
	771: res <= 3;
	772: res <= 0;
	773: res <= 0;
	774: res <= 8;
	775: res <= 3;
	776: res <= 0;
	777: res <= 8;
	778: res <= 3;
	779: res <= 0;
	780: res <= 0;
	781: res <= 0;
	782: res <= 0;
	783: res <= 0;
	784: res <= 0;
	785: res <= 7;
	786: res <= 0;
	787: res <= 0;
	788: res <= 0;
	789: res <= 0;
	790: res <= 8;
	791: res <= 15;
	792: res <= 15;
	793: res <= 15;
	794: res <= 1;
	795: res <= 0;
	796: res <= 0;
	797: res <= 0;
	798: res <= 0;
	799: res <= 0;
	800: res <= 0;
	801: res <= 0;
	802: res <= 12;
	803: res <= 1;
	804: res <= 0;
	805: res <= 0;
	806: res <= 0;
	807: res <= 0;
	808: res <= 0;
	809: res <= 0;
	810: res <= 0;
	811: res <= 7;
	812: res <= 0;
	813: res <= 0;
	814: res <= 7;
	815: res <= 8;
	816: res <= 3;
	817: res <= 0;
	818: res <= 0;
	819: res <= 8;
	820: res <= 3;
	821: res <= 0;
	822: res <= 8;
	823: res <= 3;
	824: res <= 0;
	825: res <= 0;
	826: res <= 0;
	827: res <= 0;
	828: res <= 12;
	829: res <= 15;
	830: res <= 0;
	831: res <= 0;
	832: res <= 0;
	833: res <= 0;
	834: res <= 0;
	835: res <= 8;
	836: res <= 15;
	837: res <= 15;
	838: res <= 15;
	839: res <= 1;
	840: res <= 0;
	841: res <= 0;
	842: res <= 0;
	843: res <= 0;
	844: res <= 0;
	845: res <= 0;
	846: res <= 0;
	847: res <= 12;
	848: res <= 1;
	849: res <= 0;
	850: res <= 0;
	851: res <= 0;
	852: res <= 0;
	853: res <= 0;
	854: res <= 0;
	855: res <= 0;
	856: res <= 7;
	857: res <= 0;
	858: res <= 0;
	859: res <= 7;
	860: res <= 8;
	861: res <= 3;
	862: res <= 0;
	863: res <= 0;
	864: res <= 8;
	865: res <= 3;
	866: res <= 0;
	867: res <= 8;
	868: res <= 3;
	869: res <= 0;
	870: res <= 0;
	871: res <= 0;
	872: res <= 0;
	873: res <= 12;
	874: res <= 15;
	875: res <= 0;
	876: res <= 0;
	877: res <= 0;
	878: res <= 0;
	879: res <= 0;
	880: res <= 12;
	881: res <= 15;
	882: res <= 15;
	883: res <= 15;
	884: res <= 1;
	885: res <= 0;
	886: res <= 0;
	887: res <= 0;
	888: res <= 0;
	889: res <= 0;
	890: res <= 0;
	891: res <= 0;
	892: res <= 12;
	893: res <= 1;
	894: res <= 0;
	895: res <= 0;
	896: res <= 0;
	897: res <= 0;
	898: res <= 0;
	899: res <= 0;
	900: res <= 0;
	901: res <= 0;
	902: res <= 0;
	903: res <= 0;
	904: res <= 0;
	905: res <= 0;
	906: res <= 0;
	907: res <= 0;
	908: res <= 0;
	909: res <= 0;
	910: res <= 0;
	911: res <= 0;
	912: res <= 0;
	913: res <= 0;
	914: res <= 0;
	915: res <= 0;
	916: res <= 0;
	917: res <= 0;
	918: res <= 12;
	919: res <= 15;
	920: res <= 0;
	921: res <= 0;
	922: res <= 0;
	923: res <= 0;
	924: res <= 0;
	925: res <= 14;
	926: res <= 15;
	927: res <= 15;
	928: res <= 15;
	929: res <= 0;
	930: res <= 0;
	931: res <= 0;
	932: res <= 0;
	933: res <= 0;
	934: res <= 0;
	935: res <= 0;
	936: res <= 0;
	937: res <= 0;
	938: res <= 0;
	939: res <= 0;
	940: res <= 0;
	941: res <= 0;
	942: res <= 0;
	943: res <= 0;
	944: res <= 0;
	945: res <= 0;
	946: res <= 0;
	947: res <= 0;
	948: res <= 0;
	949: res <= 0;
	950: res <= 0;
	951: res <= 0;
	952: res <= 0;
	953: res <= 0;
	954: res <= 0;
	955: res <= 0;
	956: res <= 0;
	957: res <= 0;
	958: res <= 0;
	959: res <= 0;
	960: res <= 0;
	961: res <= 0;
	962: res <= 0;
	963: res <= 0;
	964: res <= 0;
	965: res <= 0;
	966: res <= 0;
	967: res <= 0;
	968: res <= 0;
	969: res <= 0;
	970: res <= 15;
	971: res <= 15;
	972: res <= 15;
	973: res <= 15;
	974: res <= 0;
	975: res <= 0;
	976: res <= 0;
	977: res <= 0;
	978: res <= 0;
	979: res <= 0;
	980: res <= 0;
	981: res <= 0;
	982: res <= 0;
	983: res <= 0;
	984: res <= 0;
	985: res <= 0;
	986: res <= 0;
	987: res <= 0;
	988: res <= 0;
	989: res <= 0;
	990: res <= 0;
	991: res <= 0;
	992: res <= 0;
	993: res <= 0;
	994: res <= 0;
	995: res <= 0;
	996: res <= 0;
	997: res <= 0;
	998: res <= 0;
	999: res <= 0;
	1000: res <= 0;
	1001: res <= 0;
	1002: res <= 0;
	1003: res <= 0;
	1004: res <= 0;
	1005: res <= 0;
	1006: res <= 0;
	1007: res <= 0;
	1008: res <= 0;
	1009: res <= 0;
	1010: res <= 0;
	1011: res <= 0;
	1012: res <= 0;
	1013: res <= 0;
	1014: res <= 0;
	1015: res <= 15;
	1016: res <= 15;
	1017: res <= 15;
	1018: res <= 15;
	1019: res <= 0;
	1020: res <= 0;
	1021: res <= 0;
	1022: res <= 0;
	1023: res <= 0;
	1024: res <= 0;
	1025: res <= 0;
	1026: res <= 0;
	1027: res <= 0;
	1028: res <= 0;
	1029: res <= 0;
	1030: res <= 0;
	1031: res <= 0;
	1032: res <= 0;
	1033: res <= 0;
	1034: res <= 0;
	1035: res <= 0;
	1036: res <= 0;
	1037: res <= 0;
	1038: res <= 0;
	1039: res <= 0;
	1040: res <= 0;
	1041: res <= 0;
	1042: res <= 0;
	1043: res <= 0;
	1044: res <= 0;
	1045: res <= 0;
	1046: res <= 0;
	1047: res <= 0;
	1048: res <= 0;
	1049: res <= 0;
	1050: res <= 0;
	1051: res <= 0;
	1052: res <= 0;
	1053: res <= 0;
	1054: res <= 0;
	1055: res <= 0;
	1056: res <= 0;
	1057: res <= 0;
	1058: res <= 0;
	1059: res <= 8;
	1060: res <= 15;
	1061: res <= 15;
	1062: res <= 15;
	1063: res <= 7;
	1064: res <= 0;
	1065: res <= 0;
	1066: res <= 0;
	1067: res <= 0;
	1068: res <= 0;
	1069: res <= 0;
	1070: res <= 12;
	1071: res <= 1;
	1072: res <= 0;
	1073: res <= 12;
	1074: res <= 1;
	1075: res <= 0;
	1076: res <= 0;
	1077: res <= 0;
	1078: res <= 0;
	1079: res <= 0;
	1080: res <= 0;
	1081: res <= 0;
	1082: res <= 0;
	1083: res <= 0;
	1084: res <= 0;
	1085: res <= 0;
	1086: res <= 0;
	1087: res <= 0;
	1088: res <= 0;
	1089: res <= 0;
	1090: res <= 0;
	1091: res <= 0;
	1092: res <= 0;
	1093: res <= 0;
	1094: res <= 0;
	1095: res <= 0;
	1096: res <= 0;
	1097: res <= 0;
	1098: res <= 0;
	1099: res <= 0;
	1100: res <= 0;
	1101: res <= 0;
	1102: res <= 0;
	1103: res <= 0;
	1104: res <= 12;
	1105: res <= 15;
	1106: res <= 15;
	1107: res <= 15;
	1108: res <= 7;
	1109: res <= 0;
	1110: res <= 0;
	1111: res <= 0;
	1112: res <= 0;
	1113: res <= 0;
	1114: res <= 0;
	1115: res <= 12;
	1116: res <= 1;
	1117: res <= 0;
	1118: res <= 12;
	1119: res <= 1;
	1120: res <= 0;
	1121: res <= 0;
	1122: res <= 0;
	1123: res <= 0;
	1124: res <= 0;
	1125: res <= 0;
	1126: res <= 0;
	1127: res <= 0;
	1128: res <= 0;
	1129: res <= 0;
	1130: res <= 0;
	1131: res <= 0;
	1132: res <= 0;
	1133: res <= 0;
	1134: res <= 0;
	1135: res <= 0;
	1136: res <= 0;
	1137: res <= 0;
	1138: res <= 0;
	1139: res <= 0;
	1140: res <= 0;
	1141: res <= 0;
	1142: res <= 0;
	1143: res <= 0;
	1144: res <= 0;
	1145: res <= 0;
	1146: res <= 0;
	1147: res <= 0;
	1148: res <= 0;
	1149: res <= 14;
	1150: res <= 15;
	1151: res <= 15;
	1152: res <= 15;
	1153: res <= 7;
	1154: res <= 0;
	1155: res <= 0;
	1156: res <= 0;
	1157: res <= 0;
	1158: res <= 0;
	1159: res <= 0;
	1160: res <= 12;
	1161: res <= 1;
	1162: res <= 0;
	1163: res <= 12;
	1164: res <= 1;
	1165: res <= 0;
	1166: res <= 0;
	1167: res <= 0;
	1168: res <= 0;
	1169: res <= 0;
	1170: res <= 0;
	1171: res <= 0;
	1172: res <= 0;
	1173: res <= 0;
	1174: res <= 0;
	1175: res <= 0;
	1176: res <= 0;
	1177: res <= 0;
	1178: res <= 0;
	1179: res <= 0;
	1180: res <= 0;
	1181: res <= 0;
	1182: res <= 0;
	1183: res <= 0;
	1184: res <= 0;
	1185: res <= 0;
	1186: res <= 0;
	1187: res <= 0;
	1188: res <= 0;
	1189: res <= 0;
	1190: res <= 0;
	1191: res <= 0;
	1192: res <= 0;
	1193: res <= 0;
	1194: res <= 14;
	1195: res <= 15;
	1196: res <= 15;
	1197: res <= 15;
	1198: res <= 7;
	1199: res <= 0;
	1200: res <= 0;
	1201: res <= 0;
	1202: res <= 0;
	1203: res <= 0;
	1204: res <= 0;
	1205: res <= 12;
	1206: res <= 15;
	1207: res <= 8;
	1208: res <= 15;
	1209: res <= 1;
	1210: res <= 0;
	1211: res <= 0;
	1212: res <= 0;
	1213: res <= 0;
	1214: res <= 0;
	1215: res <= 8;
	1216: res <= 15;
	1217: res <= 15;
	1218: res <= 8;
	1219: res <= 3;
	1220: res <= 14;
	1221: res <= 8;
	1222: res <= 15;
	1223: res <= 7;
	1224: res <= 14;
	1225: res <= 0;
	1226: res <= 14;
	1227: res <= 12;
	1228: res <= 1;
	1229: res <= 12;
	1230: res <= 1;
	1231: res <= 0;
	1232: res <= 0;
	1233: res <= 0;
	1234: res <= 0;
	1235: res <= 0;
	1236: res <= 0;
	1237: res <= 0;
	1238: res <= 0;
	1239: res <= 15;
	1240: res <= 15;
	1241: res <= 15;
	1242: res <= 15;
	1243: res <= 3;
	1244: res <= 0;
	1245: res <= 0;
	1246: res <= 0;
	1247: res <= 0;
	1248: res <= 0;
	1249: res <= 0;
	1250: res <= 12;
	1251: res <= 15;
	1252: res <= 8;
	1253: res <= 15;
	1254: res <= 1;
	1255: res <= 0;
	1256: res <= 0;
	1257: res <= 0;
	1258: res <= 0;
	1259: res <= 0;
	1260: res <= 8;
	1261: res <= 15;
	1262: res <= 15;
	1263: res <= 8;
	1264: res <= 3;
	1265: res <= 14;
	1266: res <= 8;
	1267: res <= 15;
	1268: res <= 7;
	1269: res <= 14;
	1270: res <= 0;
	1271: res <= 14;
	1272: res <= 12;
	1273: res <= 1;
	1274: res <= 12;
	1275: res <= 1;
	1276: res <= 0;
	1277: res <= 0;
	1278: res <= 0;
	1279: res <= 0;
	1280: res <= 0;
	1281: res <= 0;
	1282: res <= 0;
	1283: res <= 8;
	1284: res <= 15;
	1285: res <= 15;
	1286: res <= 15;
	1287: res <= 15;
	1288: res <= 3;
	1289: res <= 0;
	1290: res <= 0;
	1291: res <= 0;
	1292: res <= 0;
	1293: res <= 0;
	1294: res <= 0;
	1295: res <= 12;
	1296: res <= 15;
	1297: res <= 8;
	1298: res <= 15;
	1299: res <= 1;
	1300: res <= 0;
	1301: res <= 0;
	1302: res <= 0;
	1303: res <= 0;
	1304: res <= 0;
	1305: res <= 8;
	1306: res <= 15;
	1307: res <= 15;
	1308: res <= 8;
	1309: res <= 3;
	1310: res <= 14;
	1311: res <= 8;
	1312: res <= 15;
	1313: res <= 7;
	1314: res <= 14;
	1315: res <= 0;
	1316: res <= 14;
	1317: res <= 12;
	1318: res <= 15;
	1319: res <= 12;
	1320: res <= 1;
	1321: res <= 0;
	1322: res <= 0;
	1323: res <= 0;
	1324: res <= 0;
	1325: res <= 0;
	1326: res <= 0;
	1327: res <= 0;
	1328: res <= 8;
	1329: res <= 15;
	1330: res <= 15;
	1331: res <= 15;
	1332: res <= 15;
	1333: res <= 3;
	1334: res <= 0;
	1335: res <= 0;
	1336: res <= 0;
	1337: res <= 0;
	1338: res <= 0;
	1339: res <= 0;
	1340: res <= 12;
	1341: res <= 1;
	1342: res <= 7;
	1343: res <= 12;
	1344: res <= 1;
	1345: res <= 0;
	1346: res <= 0;
	1347: res <= 0;
	1348: res <= 0;
	1349: res <= 0;
	1350: res <= 0;
	1351: res <= 12;
	1352: res <= 1;
	1353: res <= 8;
	1354: res <= 3;
	1355: res <= 14;
	1356: res <= 8;
	1357: res <= 3;
	1358: res <= 7;
	1359: res <= 14;
	1360: res <= 0;
	1361: res <= 14;
	1362: res <= 12;
	1363: res <= 15;
	1364: res <= 12;
	1365: res <= 1;
	1366: res <= 0;
	1367: res <= 0;
	1368: res <= 0;
	1369: res <= 0;
	1370: res <= 0;
	1371: res <= 0;
	1372: res <= 0;
	1373: res <= 12;
	1374: res <= 15;
	1375: res <= 15;
	1376: res <= 15;
	1377: res <= 15;
	1378: res <= 1;
	1379: res <= 0;
	1380: res <= 0;
	1381: res <= 0;
	1382: res <= 0;
	1383: res <= 0;
	1384: res <= 0;
	1385: res <= 12;
	1386: res <= 1;
	1387: res <= 7;
	1388: res <= 12;
	1389: res <= 1;
	1390: res <= 0;
	1391: res <= 0;
	1392: res <= 0;
	1393: res <= 0;
	1394: res <= 0;
	1395: res <= 0;
	1396: res <= 12;
	1397: res <= 1;
	1398: res <= 8;
	1399: res <= 15;
	1400: res <= 15;
	1401: res <= 8;
	1402: res <= 3;
	1403: res <= 7;
	1404: res <= 14;
	1405: res <= 0;
	1406: res <= 14;
	1407: res <= 12;
	1408: res <= 15;
	1409: res <= 12;
	1410: res <= 1;
	1411: res <= 0;
	1412: res <= 0;
	1413: res <= 0;
	1414: res <= 0;
	1415: res <= 0;
	1416: res <= 0;
	1417: res <= 0;
	1418: res <= 14;
	1419: res <= 15;
	1420: res <= 15;
	1421: res <= 15;
	1422: res <= 15;
	1423: res <= 1;
	1424: res <= 0;
	1425: res <= 0;
	1426: res <= 0;
	1427: res <= 3;
	1428: res <= 0;
	1429: res <= 0;
	1430: res <= 12;
	1431: res <= 1;
	1432: res <= 7;
	1433: res <= 12;
	1434: res <= 1;
	1435: res <= 0;
	1436: res <= 0;
	1437: res <= 0;
	1438: res <= 0;
	1439: res <= 0;
	1440: res <= 0;
	1441: res <= 12;
	1442: res <= 1;
	1443: res <= 8;
	1444: res <= 15;
	1445: res <= 15;
	1446: res <= 8;
	1447: res <= 3;
	1448: res <= 7;
	1449: res <= 14;
	1450: res <= 0;
	1451: res <= 14;
	1452: res <= 12;
	1453: res <= 9;
	1454: res <= 15;
	1455: res <= 1;
	1456: res <= 0;
	1457: res <= 0;
	1458: res <= 0;
	1459: res <= 0;
	1460: res <= 15;
	1461: res <= 15;
	1462: res <= 1;
	1463: res <= 14;
	1464: res <= 15;
	1465: res <= 15;
	1466: res <= 15;
	1467: res <= 15;
	1468: res <= 0;
	1469: res <= 0;
	1470: res <= 0;
	1471: res <= 12;
	1472: res <= 3;
	1473: res <= 0;
	1474: res <= 0;
	1475: res <= 12;
	1476: res <= 1;
	1477: res <= 0;
	1478: res <= 12;
	1479: res <= 1;
	1480: res <= 0;
	1481: res <= 0;
	1482: res <= 0;
	1483: res <= 0;
	1484: res <= 0;
	1485: res <= 0;
	1486: res <= 12;
	1487: res <= 1;
	1488: res <= 8;
	1489: res <= 15;
	1490: res <= 15;
	1491: res <= 8;
	1492: res <= 3;
	1493: res <= 7;
	1494: res <= 14;
	1495: res <= 0;
	1496: res <= 14;
	1497: res <= 12;
	1498: res <= 9;
	1499: res <= 15;
	1500: res <= 1;
	1501: res <= 0;
	1502: res <= 0;
	1503: res <= 0;
	1504: res <= 15;
	1505: res <= 15;
	1506: res <= 15;
	1507: res <= 7;
	1508: res <= 15;
	1509: res <= 15;
	1510: res <= 15;
	1511: res <= 15;
	1512: res <= 15;
	1513: res <= 0;
	1514: res <= 0;
	1515: res <= 0;
	1516: res <= 14;
	1517: res <= 3;
	1518: res <= 0;
	1519: res <= 0;
	1520: res <= 12;
	1521: res <= 1;
	1522: res <= 0;
	1523: res <= 12;
	1524: res <= 1;
	1525: res <= 0;
	1526: res <= 0;
	1527: res <= 0;
	1528: res <= 0;
	1529: res <= 0;
	1530: res <= 0;
	1531: res <= 12;
	1532: res <= 1;
	1533: res <= 8;
	1534: res <= 3;
	1535: res <= 14;
	1536: res <= 8;
	1537: res <= 15;
	1538: res <= 7;
	1539: res <= 14;
	1540: res <= 7;
	1541: res <= 14;
	1542: res <= 12;
	1543: res <= 9;
	1544: res <= 15;
	1545: res <= 1;
	1546: res <= 0;
	1547: res <= 0;
	1548: res <= 15;
	1549: res <= 15;
	1550: res <= 15;
	1551: res <= 15;
	1552: res <= 3;
	1553: res <= 15;
	1554: res <= 15;
	1555: res <= 15;
	1556: res <= 15;
	1557: res <= 7;
	1558: res <= 0;
	1559: res <= 0;
	1560: res <= 8;
	1561: res <= 15;
	1562: res <= 3;
	1563: res <= 0;
	1564: res <= 0;
	1565: res <= 12;
	1566: res <= 1;
	1567: res <= 0;
	1568: res <= 12;
	1569: res <= 1;
	1570: res <= 0;
	1571: res <= 0;
	1572: res <= 0;
	1573: res <= 0;
	1574: res <= 0;
	1575: res <= 0;
	1576: res <= 12;
	1577: res <= 1;
	1578: res <= 8;
	1579: res <= 3;
	1580: res <= 14;
	1581: res <= 8;
	1582: res <= 15;
	1583: res <= 7;
	1584: res <= 14;
	1585: res <= 7;
	1586: res <= 14;
	1587: res <= 12;
	1588: res <= 1;
	1589: res <= 12;
	1590: res <= 1;
	1591: res <= 0;
	1592: res <= 12;
	1593: res <= 15;
	1594: res <= 15;
	1595: res <= 15;
	1596: res <= 15;
	1597: res <= 11;
	1598: res <= 15;
	1599: res <= 15;
	1600: res <= 15;
	1601: res <= 15;
	1602: res <= 7;
	1603: res <= 0;
	1604: res <= 0;
	1605: res <= 14;
	1606: res <= 15;
	1607: res <= 3;
	1608: res <= 0;
	1609: res <= 0;
	1610: res <= 12;
	1611: res <= 1;
	1612: res <= 0;
	1613: res <= 12;
	1614: res <= 1;
	1615: res <= 0;
	1616: res <= 0;
	1617: res <= 0;
	1618: res <= 0;
	1619: res <= 0;
	1620: res <= 0;
	1621: res <= 12;
	1622: res <= 1;
	1623: res <= 8;
	1624: res <= 3;
	1625: res <= 14;
	1626: res <= 8;
	1627: res <= 15;
	1628: res <= 7;
	1629: res <= 14;
	1630: res <= 7;
	1631: res <= 14;
	1632: res <= 12;
	1633: res <= 1;
	1634: res <= 12;
	1635: res <= 1;
	1636: res <= 0;
	1637: res <= 15;
	1638: res <= 15;
	1639: res <= 15;
	1640: res <= 15;
	1641: res <= 15;
	1642: res <= 13;
	1643: res <= 15;
	1644: res <= 15;
	1645: res <= 15;
	1646: res <= 15;
	1647: res <= 7;
	1648: res <= 0;
	1649: res <= 0;
	1650: res <= 15;
	1651: res <= 15;
	1652: res <= 3;
	1653: res <= 0;
	1654: res <= 0;
	1655: res <= 12;
	1656: res <= 1;
	1657: res <= 0;
	1658: res <= 12;
	1659: res <= 1;
	1660: res <= 0;
	1661: res <= 0;
	1662: res <= 0;
	1663: res <= 0;
	1664: res <= 0;
	1665: res <= 0;
	1666: res <= 0;
	1667: res <= 0;
	1668: res <= 0;
	1669: res <= 0;
	1670: res <= 0;
	1671: res <= 0;
	1672: res <= 0;
	1673: res <= 0;
	1674: res <= 0;
	1675: res <= 0;
	1676: res <= 0;
	1677: res <= 0;
	1678: res <= 0;
	1679: res <= 0;
	1680: res <= 0;
	1681: res <= 8;
	1682: res <= 15;
	1683: res <= 15;
	1684: res <= 15;
	1685: res <= 15;
	1686: res <= 15;
	1687: res <= 13;
	1688: res <= 15;
	1689: res <= 15;
	1690: res <= 15;
	1691: res <= 15;
	1692: res <= 3;
	1693: res <= 0;
	1694: res <= 8;
	1695: res <= 15;
	1696: res <= 15;
	1697: res <= 3;
	1698: res <= 0;
	1699: res <= 0;
	1700: res <= 12;
	1701: res <= 1;
	1702: res <= 0;
	1703: res <= 12;
	1704: res <= 1;
	1705: res <= 0;
	1706: res <= 0;
	1707: res <= 0;
	1708: res <= 0;
	1709: res <= 0;
	1710: res <= 0;
	1711: res <= 0;
	1712: res <= 0;
	1713: res <= 0;
	1714: res <= 0;
	1715: res <= 0;
	1716: res <= 0;
	1717: res <= 0;
	1718: res <= 0;
	1719: res <= 0;
	1720: res <= 0;
	1721: res <= 0;
	1722: res <= 0;
	1723: res <= 0;
	1724: res <= 0;
	1725: res <= 0;
	1726: res <= 14;
	1727: res <= 15;
	1728: res <= 15;
	1729: res <= 15;
	1730: res <= 1;
	1731: res <= 0;
	1732: res <= 12;
	1733: res <= 15;
	1734: res <= 15;
	1735: res <= 15;
	1736: res <= 15;
	1737: res <= 3;
	1738: res <= 0;
	1739: res <= 12;
	1740: res <= 15;
	1741: res <= 15;
	1742: res <= 3;
	1743: res <= 0;
	1744: res <= 0;
	1745: res <= 0;
	1746: res <= 0;
	1747: res <= 0;
	1748: res <= 0;
	1749: res <= 0;
	1750: res <= 0;
	1751: res <= 0;
	1752: res <= 0;
	1753: res <= 0;
	1754: res <= 0;
	1755: res <= 0;
	1756: res <= 0;
	1757: res <= 0;
	1758: res <= 0;
	1759: res <= 0;
	1760: res <= 0;
	1761: res <= 0;
	1762: res <= 0;
	1763: res <= 0;
	1764: res <= 0;
	1765: res <= 0;
	1766: res <= 0;
	1767: res <= 0;
	1768: res <= 0;
	1769: res <= 0;
	1770: res <= 0;
	1771: res <= 15;
	1772: res <= 15;
	1773: res <= 15;
	1774: res <= 0;
	1775: res <= 0;
	1776: res <= 0;
	1777: res <= 14;
	1778: res <= 15;
	1779: res <= 15;
	1780: res <= 15;
	1781: res <= 15;
	1782: res <= 3;
	1783: res <= 0;
	1784: res <= 15;
	1785: res <= 15;
	1786: res <= 15;
	1787: res <= 1;
	1788: res <= 0;
	1789: res <= 0;
	1790: res <= 0;
	1791: res <= 0;
	1792: res <= 0;
	1793: res <= 0;
	1794: res <= 0;
	1795: res <= 0;
	1796: res <= 0;
	1797: res <= 0;
	1798: res <= 0;
	1799: res <= 0;
	1800: res <= 0;
	1801: res <= 0;
	1802: res <= 0;
	1803: res <= 0;
	1804: res <= 0;
	1805: res <= 0;
	1806: res <= 0;
	1807: res <= 0;
	1808: res <= 0;
	1809: res <= 0;
	1810: res <= 0;
	1811: res <= 0;
	1812: res <= 0;
	1813: res <= 0;
	1814: res <= 0;
	1815: res <= 8;
	1816: res <= 15;
	1817: res <= 15;
	1818: res <= 1;
	1819: res <= 0;
	1820: res <= 0;
	1821: res <= 0;
	1822: res <= 15;
	1823: res <= 15;
	1824: res <= 15;
	1825: res <= 15;
	1826: res <= 15;
	1827: res <= 1;
	1828: res <= 8;
	1829: res <= 15;
	1830: res <= 15;
	1831: res <= 15;
	1832: res <= 1;
	1833: res <= 0;
	1834: res <= 0;
	1835: res <= 0;
	1836: res <= 0;
	1837: res <= 0;
	1838: res <= 0;
	1839: res <= 0;
	1840: res <= 0;
	1841: res <= 0;
	1842: res <= 0;
	1843: res <= 0;
	1844: res <= 0;
	1845: res <= 0;
	1846: res <= 0;
	1847: res <= 0;
	1848: res <= 0;
	1849: res <= 0;
	1850: res <= 0;
	1851: res <= 0;
	1852: res <= 0;
	1853: res <= 0;
	1854: res <= 0;
	1855: res <= 0;
	1856: res <= 0;
	1857: res <= 0;
	1858: res <= 0;
	1859: res <= 0;
	1860: res <= 14;
	1861: res <= 15;
	1862: res <= 7;
	1863: res <= 0;
	1864: res <= 0;
	1865: res <= 0;
	1866: res <= 0;
	1867: res <= 15;
	1868: res <= 15;
	1869: res <= 15;
	1870: res <= 15;
	1871: res <= 15;
	1872: res <= 1;
	1873: res <= 12;
	1874: res <= 15;
	1875: res <= 15;
	1876: res <= 15;
	1877: res <= 1;
	1878: res <= 0;
	1879: res <= 0;
	1880: res <= 0;
	1881: res <= 0;
	1882: res <= 0;
	1883: res <= 0;
	1884: res <= 0;
	1885: res <= 0;
	1886: res <= 0;
	1887: res <= 0;
	1888: res <= 0;
	1889: res <= 0;
	1890: res <= 0;
	1891: res <= 0;
	1892: res <= 0;
	1893: res <= 0;
	1894: res <= 0;
	1895: res <= 0;
	1896: res <= 0;
	1897: res <= 0;
	1898: res <= 0;
	1899: res <= 0;
	1900: res <= 0;
	1901: res <= 0;
	1902: res <= 0;
	1903: res <= 0;
	1904: res <= 0;
	1905: res <= 15;
	1906: res <= 15;
	1907: res <= 3;
	1908: res <= 0;
	1909: res <= 0;
	1910: res <= 0;
	1911: res <= 0;
	1912: res <= 15;
	1913: res <= 15;
	1914: res <= 15;
	1915: res <= 15;
	1916: res <= 15;
	1917: res <= 0;
	1918: res <= 14;
	1919: res <= 15;
	1920: res <= 15;
	1921: res <= 15;
	1922: res <= 0;
	1923: res <= 0;
	1924: res <= 0;
	1925: res <= 0;
	1926: res <= 0;
	1927: res <= 0;
	1928: res <= 0;
	1929: res <= 0;
	1930: res <= 0;
	1931: res <= 0;
	1932: res <= 0;
	1933: res <= 0;
	1934: res <= 0;
	1935: res <= 0;
	1936: res <= 0;
	1937: res <= 0;
	1938: res <= 0;
	1939: res <= 0;
	1940: res <= 0;
	1941: res <= 0;
	1942: res <= 0;
	1943: res <= 0;
	1944: res <= 0;
	1945: res <= 0;
	1946: res <= 0;
	1947: res <= 0;
	1948: res <= 0;
	1949: res <= 0;
	1950: res <= 15;
	1951: res <= 15;
	1952: res <= 0;
	1953: res <= 0;
	1954: res <= 0;
	1955: res <= 0;
	1956: res <= 8;
	1957: res <= 15;
	1958: res <= 15;
	1959: res <= 15;
	1960: res <= 15;
	1961: res <= 15;
	1962: res <= 0;
	1963: res <= 15;
	1964: res <= 15;
	1965: res <= 15;
	1966: res <= 15;
	1967: res <= 0;
	1968: res <= 0;
	1969: res <= 0;
	1970: res <= 0;
	1971: res <= 12;
	1972: res <= 15;
	1973: res <= 0;
	1974: res <= 0;
	1975: res <= 0;
	1976: res <= 0;
	1977: res <= 0;
	1978: res <= 0;
	1979: res <= 0;
	1980: res <= 0;
	1981: res <= 0;
	1982: res <= 0;
	1983: res <= 0;
	1984: res <= 0;
	1985: res <= 0;
	1986: res <= 0;
	1987: res <= 0;
	1988: res <= 0;
	1989: res <= 0;
	1990: res <= 0;
	1991: res <= 0;
	1992: res <= 0;
	1993: res <= 0;
	1994: res <= 8;
	1995: res <= 15;
	1996: res <= 7;
	1997: res <= 0;
	1998: res <= 0;
	1999: res <= 0;
	2000: res <= 0;
	2001: res <= 8;
	2002: res <= 15;
	2003: res <= 15;
	2004: res <= 15;
	2005: res <= 15;
	2006: res <= 7;
	2007: res <= 12;
	2008: res <= 15;
	2009: res <= 15;
	2010: res <= 15;
	2011: res <= 15;
	2012: res <= 0;
	2013: res <= 0;
	2014: res <= 0;
	2015: res <= 0;
	2016: res <= 12;
	2017: res <= 15;
	2018: res <= 0;
	2019: res <= 0;
	2020: res <= 0;
	2021: res <= 0;
	2022: res <= 0;
	2023: res <= 0;
	2024: res <= 0;
	2025: res <= 0;
	2026: res <= 0;
	2027: res <= 0;
	2028: res <= 0;
	2029: res <= 0;
	2030: res <= 0;
	2031: res <= 0;
	2032: res <= 0;
	2033: res <= 0;
	2034: res <= 0;
	2035: res <= 0;
	2036: res <= 0;
	2037: res <= 0;
	2038: res <= 0;
	2039: res <= 12;
	2040: res <= 15;
	2041: res <= 3;
	2042: res <= 0;
	2043: res <= 0;
	2044: res <= 0;
	2045: res <= 0;
	2046: res <= 12;
	2047: res <= 15;
	2048: res <= 15;
	2049: res <= 15;
	2050: res <= 15;
	2051: res <= 7;
	2052: res <= 14;
	2053: res <= 15;
	2054: res <= 15;
	2055: res <= 15;
	2056: res <= 7;
	2057: res <= 0;
	2058: res <= 0;
	2059: res <= 0;
	2060: res <= 0;
	2061: res <= 12;
	2062: res <= 15;
	2063: res <= 0;
	2064: res <= 0;
	2065: res <= 0;
	2066: res <= 0;
	2067: res <= 0;
	2068: res <= 0;
	2069: res <= 0;
	2070: res <= 0;
	2071: res <= 0;
	2072: res <= 0;
	2073: res <= 0;
	2074: res <= 0;
	2075: res <= 0;
	2076: res <= 0;
	2077: res <= 0;
	2078: res <= 0;
	2079: res <= 0;
	2080: res <= 0;
	2081: res <= 0;
	2082: res <= 0;
	2083: res <= 0;
	2084: res <= 14;
	2085: res <= 15;
	2086: res <= 1;
	2087: res <= 0;
	2088: res <= 0;
	2089: res <= 0;
	2090: res <= 0;
	2091: res <= 12;
	2092: res <= 15;
	2093: res <= 15;
	2094: res <= 15;
	2095: res <= 15;
	2096: res <= 3;
	2097: res <= 15;
	2098: res <= 15;
	2099: res <= 15;
	2100: res <= 15;
	2101: res <= 3;
	2102: res <= 0;
	2103: res <= 0;
	2104: res <= 0;
	2105: res <= 0;
	2106: res <= 12;
	2107: res <= 1;
	2108: res <= 7;
	2109: res <= 0;
	2110: res <= 0;
	2111: res <= 0;
	2112: res <= 0;
	2113: res <= 0;
	2114: res <= 0;
	2115: res <= 0;
	2116: res <= 0;
	2117: res <= 0;
	2118: res <= 0;
	2119: res <= 0;
	2120: res <= 0;
	2121: res <= 0;
	2122: res <= 0;
	2123: res <= 0;
	2124: res <= 0;
	2125: res <= 0;
	2126: res <= 0;
	2127: res <= 0;
	2128: res <= 0;
	2129: res <= 14;
	2130: res <= 15;
	2131: res <= 0;
	2132: res <= 0;
	2133: res <= 0;
	2134: res <= 0;
	2135: res <= 0;
	2136: res <= 14;
	2137: res <= 15;
	2138: res <= 15;
	2139: res <= 15;
	2140: res <= 15;
	2141: res <= 9;
	2142: res <= 15;
	2143: res <= 15;
	2144: res <= 15;
	2145: res <= 15;
	2146: res <= 3;
	2147: res <= 0;
	2148: res <= 0;
	2149: res <= 0;
	2150: res <= 0;
	2151: res <= 12;
	2152: res <= 1;
	2153: res <= 7;
	2154: res <= 0;
	2155: res <= 0;
	2156: res <= 0;
	2157: res <= 0;
	2158: res <= 0;
	2159: res <= 0;
	2160: res <= 0;
	2161: res <= 0;
	2162: res <= 0;
	2163: res <= 0;
	2164: res <= 0;
	2165: res <= 0;
	2166: res <= 0;
	2167: res <= 0;
	2168: res <= 0;
	2169: res <= 0;
	2170: res <= 0;
	2171: res <= 0;
	2172: res <= 0;
	2173: res <= 0;
	2174: res <= 15;
	2175: res <= 7;
	2176: res <= 0;
	2177: res <= 0;
	2178: res <= 0;
	2179: res <= 0;
	2180: res <= 0;
	2181: res <= 14;
	2182: res <= 15;
	2183: res <= 15;
	2184: res <= 15;
	2185: res <= 15;
	2186: res <= 12;
	2187: res <= 15;
	2188: res <= 15;
	2189: res <= 15;
	2190: res <= 15;
	2191: res <= 1;
	2192: res <= 0;
	2193: res <= 0;
	2194: res <= 0;
	2195: res <= 0;
	2196: res <= 12;
	2197: res <= 1;
	2198: res <= 7;
	2199: res <= 0;
	2200: res <= 0;
	2201: res <= 0;
	2202: res <= 0;
	2203: res <= 0;
	2204: res <= 0;
	2205: res <= 0;
	2206: res <= 0;
	2207: res <= 0;
	2208: res <= 0;
	2209: res <= 0;
	2210: res <= 0;
	2211: res <= 0;
	2212: res <= 0;
	2213: res <= 0;
	2214: res <= 0;
	2215: res <= 0;
	2216: res <= 0;
	2217: res <= 0;
	2218: res <= 8;
	2219: res <= 15;
	2220: res <= 3;
	2221: res <= 0;
	2222: res <= 0;
	2223: res <= 0;
	2224: res <= 0;
	2225: res <= 0;
	2226: res <= 14;
	2227: res <= 15;
	2228: res <= 15;
	2229: res <= 15;
	2230: res <= 7;
	2231: res <= 14;
	2232: res <= 15;
	2233: res <= 15;
	2234: res <= 15;
	2235: res <= 15;
	2236: res <= 0;
	2237: res <= 0;
	2238: res <= 0;
	2239: res <= 0;
	2240: res <= 0;
	2241: res <= 12;
	2242: res <= 1;
	2243: res <= 7;
	2244: res <= 0;
	2245: res <= 0;
	2246: res <= 0;
	2247: res <= 0;
	2248: res <= 0;
	2249: res <= 0;
	2250: res <= 0;
	2251: res <= 0;
	2252: res <= 0;
	2253: res <= 0;
	2254: res <= 0;
	2255: res <= 0;
	2256: res <= 0;
	2257: res <= 0;
	2258: res <= 0;
	2259: res <= 0;
	2260: res <= 0;
	2261: res <= 0;
	2262: res <= 0;
	2263: res <= 8;
	2264: res <= 15;
	2265: res <= 3;
	2266: res <= 0;
	2267: res <= 0;
	2268: res <= 0;
	2269: res <= 0;
	2270: res <= 0;
	2271: res <= 15;
	2272: res <= 15;
	2273: res <= 15;
	2274: res <= 15;
	2275: res <= 3;
	2276: res <= 15;
	2277: res <= 15;
	2278: res <= 15;
	2279: res <= 15;
	2280: res <= 7;
	2281: res <= 0;
	2282: res <= 0;
	2283: res <= 0;
	2284: res <= 0;
	2285: res <= 0;
	2286: res <= 12;
	2287: res <= 1;
	2288: res <= 7;
	2289: res <= 0;
	2290: res <= 0;
	2291: res <= 0;
	2292: res <= 0;
	2293: res <= 0;
	2294: res <= 0;
	2295: res <= 0;
	2296: res <= 0;
	2297: res <= 0;
	2298: res <= 0;
	2299: res <= 0;
	2300: res <= 0;
	2301: res <= 0;
	2302: res <= 0;
	2303: res <= 0;
	2304: res <= 0;
	2305: res <= 0;
	2306: res <= 0;
	2307: res <= 0;
	2308: res <= 12;
	2309: res <= 15;
	2310: res <= 1;
	2311: res <= 0;
	2312: res <= 0;
	2313: res <= 0;
	2314: res <= 0;
	2315: res <= 0;
	2316: res <= 15;
	2317: res <= 15;
	2318: res <= 15;
	2319: res <= 15;
	2320: res <= 9;
	2321: res <= 15;
	2322: res <= 15;
	2323: res <= 15;
	2324: res <= 15;
	2325: res <= 7;
	2326: res <= 0;
	2327: res <= 0;
	2328: res <= 0;
	2329: res <= 0;
	2330: res <= 0;
	2331: res <= 12;
	2332: res <= 1;
	2333: res <= 7;
	2334: res <= 0;
	2335: res <= 0;
	2336: res <= 0;
	2337: res <= 0;
	2338: res <= 0;
	2339: res <= 0;
	2340: res <= 0;
	2341: res <= 0;
	2342: res <= 0;
	2343: res <= 0;
	2344: res <= 0;
	2345: res <= 0;
	2346: res <= 0;
	2347: res <= 0;
	2348: res <= 0;
	2349: res <= 0;
	2350: res <= 0;
	2351: res <= 0;
	2352: res <= 0;
	2353: res <= 12;
	2354: res <= 15;
	2355: res <= 0;
	2356: res <= 0;
	2357: res <= 0;
	2358: res <= 0;
	2359: res <= 0;
	2360: res <= 8;
	2361: res <= 15;
	2362: res <= 15;
	2363: res <= 15;
	2364: res <= 15;
	2365: res <= 12;
	2366: res <= 15;
	2367: res <= 15;
	2368: res <= 15;
	2369: res <= 15;
	2370: res <= 3;
	2371: res <= 0;
	2372: res <= 0;
	2373: res <= 0;
	2374: res <= 0;
	2375: res <= 0;
	2376: res <= 12;
	2377: res <= 15;
	2378: res <= 0;
	2379: res <= 0;
	2380: res <= 0;
	2381: res <= 0;
	2382: res <= 0;
	2383: res <= 0;
	2384: res <= 0;
	2385: res <= 0;
	2386: res <= 0;
	2387: res <= 0;
	2388: res <= 0;
	2389: res <= 0;
	2390: res <= 0;
	2391: res <= 0;
	2392: res <= 0;
	2393: res <= 0;
	2394: res <= 0;
	2395: res <= 0;
	2396: res <= 0;
	2397: res <= 0;
	2398: res <= 12;
	2399: res <= 15;
	2400: res <= 0;
	2401: res <= 0;
	2402: res <= 0;
	2403: res <= 0;
	2404: res <= 0;
	2405: res <= 8;
	2406: res <= 15;
	2407: res <= 15;
	2408: res <= 15;
	2409: res <= 7;
	2410: res <= 14;
	2411: res <= 15;
	2412: res <= 15;
	2413: res <= 15;
	2414: res <= 15;
	2415: res <= 1;
	2416: res <= 0;
	2417: res <= 0;
	2418: res <= 0;
	2419: res <= 0;
	2420: res <= 0;
	2421: res <= 12;
	2422: res <= 15;
	2423: res <= 0;
	2424: res <= 0;
	2425: res <= 0;
	2426: res <= 0;
	2427: res <= 0;
	2428: res <= 0;
	2429: res <= 0;
	2430: res <= 0;
	2431: res <= 0;
	2432: res <= 0;
	2433: res <= 0;
	2434: res <= 0;
	2435: res <= 0;
	2436: res <= 0;
	2437: res <= 0;
	2438: res <= 0;
	2439: res <= 0;
	2440: res <= 0;
	2441: res <= 0;
	2442: res <= 0;
	2443: res <= 14;
	2444: res <= 7;
	2445: res <= 0;
	2446: res <= 0;
	2447: res <= 0;
	2448: res <= 0;
	2449: res <= 0;
	2450: res <= 8;
	2451: res <= 15;
	2452: res <= 15;
	2453: res <= 15;
	2454: res <= 3;
	2455: res <= 15;
	2456: res <= 15;
	2457: res <= 15;
	2458: res <= 15;
	2459: res <= 15;
	2460: res <= 0;
	2461: res <= 0;
	2462: res <= 0;
	2463: res <= 0;
	2464: res <= 0;
	2465: res <= 0;
	2466: res <= 12;
	2467: res <= 15;
	2468: res <= 0;
	2469: res <= 0;
	2470: res <= 0;
	2471: res <= 0;
	2472: res <= 0;
	2473: res <= 0;
	2474: res <= 0;
	2475: res <= 0;
	2476: res <= 0;
	2477: res <= 0;
	2478: res <= 0;
	2479: res <= 0;
	2480: res <= 0;
	2481: res <= 0;
	2482: res <= 0;
	2483: res <= 0;
	2484: res <= 0;
	2485: res <= 0;
	2486: res <= 0;
	2487: res <= 0;
	2488: res <= 14;
	2489: res <= 7;
	2490: res <= 0;
	2491: res <= 0;
	2492: res <= 0;
	2493: res <= 0;
	2494: res <= 0;
	2495: res <= 12;
	2496: res <= 15;
	2497: res <= 15;
	2498: res <= 15;
	2499: res <= 9;
	2500: res <= 15;
	2501: res <= 15;
	2502: res <= 15;
	2503: res <= 15;
	2504: res <= 7;
	2505: res <= 0;
	2506: res <= 0;
	2507: res <= 0;
	2508: res <= 0;
	2509: res <= 0;
	2510: res <= 0;
	2511: res <= 12;
	2512: res <= 1;
	2513: res <= 7;
	2514: res <= 0;
	2515: res <= 0;
	2516: res <= 0;
	2517: res <= 0;
	2518: res <= 0;
	2519: res <= 0;
	2520: res <= 0;
	2521: res <= 0;
	2522: res <= 0;
	2523: res <= 0;
	2524: res <= 0;
	2525: res <= 0;
	2526: res <= 0;
	2527: res <= 0;
	2528: res <= 0;
	2529: res <= 0;
	2530: res <= 0;
	2531: res <= 0;
	2532: res <= 0;
	2533: res <= 14;
	2534: res <= 7;
	2535: res <= 0;
	2536: res <= 0;
	2537: res <= 0;
	2538: res <= 0;
	2539: res <= 0;
	2540: res <= 12;
	2541: res <= 15;
	2542: res <= 15;
	2543: res <= 15;
	2544: res <= 12;
	2545: res <= 15;
	2546: res <= 15;
	2547: res <= 15;
	2548: res <= 15;
	2549: res <= 3;
	2550: res <= 0;
	2551: res <= 0;
	2552: res <= 0;
	2553: res <= 0;
	2554: res <= 0;
	2555: res <= 0;
	2556: res <= 12;
	2557: res <= 1;
	2558: res <= 7;
	2559: res <= 0;
	2560: res <= 0;
	2561: res <= 0;
	2562: res <= 0;
	2563: res <= 0;
	2564: res <= 0;
	2565: res <= 0;
	2566: res <= 0;
	2567: res <= 0;
	2568: res <= 0;
	2569: res <= 0;
	2570: res <= 0;
	2571: res <= 0;
	2572: res <= 0;
	2573: res <= 0;
	2574: res <= 0;
	2575: res <= 0;
	2576: res <= 0;
	2577: res <= 0;
	2578: res <= 15;
	2579: res <= 7;
	2580: res <= 0;
	2581: res <= 0;
	2582: res <= 0;
	2583: res <= 0;
	2584: res <= 0;
	2585: res <= 14;
	2586: res <= 15;
	2587: res <= 15;
	2588: res <= 15;
	2589: res <= 14;
	2590: res <= 15;
	2591: res <= 15;
	2592: res <= 15;
	2593: res <= 15;
	2594: res <= 3;
	2595: res <= 0;
	2596: res <= 0;
	2597: res <= 0;
	2598: res <= 0;
	2599: res <= 0;
	2600: res <= 0;
	2601: res <= 12;
	2602: res <= 1;
	2603: res <= 7;
	2604: res <= 0;
	2605: res <= 0;
	2606: res <= 0;
	2607: res <= 0;
	2608: res <= 0;
	2609: res <= 0;
	2610: res <= 0;
	2611: res <= 0;
	2612: res <= 0;
	2613: res <= 0;
	2614: res <= 0;
	2615: res <= 0;
	2616: res <= 0;
	2617: res <= 0;
	2618: res <= 0;
	2619: res <= 0;
	2620: res <= 0;
	2621: res <= 0;
	2622: res <= 0;
	2623: res <= 15;
	2624: res <= 3;
	2625: res <= 0;
	2626: res <= 0;
	2627: res <= 0;
	2628: res <= 0;
	2629: res <= 0;
	2630: res <= 14;
	2631: res <= 15;
	2632: res <= 15;
	2633: res <= 7;
	2634: res <= 15;
	2635: res <= 15;
	2636: res <= 15;
	2637: res <= 15;
	2638: res <= 15;
	2639: res <= 1;
	2640: res <= 0;
	2641: res <= 0;
	2642: res <= 0;
	2643: res <= 0;
	2644: res <= 0;
	2645: res <= 0;
	2646: res <= 12;
	2647: res <= 1;
	2648: res <= 7;
	2649: res <= 0;
	2650: res <= 0;
	2651: res <= 0;
	2652: res <= 0;
	2653: res <= 0;
	2654: res <= 0;
	2655: res <= 0;
	2656: res <= 0;
	2657: res <= 0;
	2658: res <= 0;
	2659: res <= 0;
	2660: res <= 0;
	2661: res <= 0;
	2662: res <= 0;
	2663: res <= 0;
	2664: res <= 0;
	2665: res <= 0;
	2666: res <= 0;
	2667: res <= 0;
	2668: res <= 15;
	2669: res <= 3;
	2670: res <= 0;
	2671: res <= 0;
	2672: res <= 0;
	2673: res <= 0;
	2674: res <= 0;
	2675: res <= 14;
	2676: res <= 15;
	2677: res <= 15;
	2678: res <= 11;
	2679: res <= 15;
	2680: res <= 15;
	2681: res <= 15;
	2682: res <= 15;
	2683: res <= 15;
	2684: res <= 0;
	2685: res <= 0;
	2686: res <= 0;
	2687: res <= 0;
	2688: res <= 0;
	2689: res <= 0;
	2690: res <= 0;
	2691: res <= 12;
	2692: res <= 1;
	2693: res <= 7;
	2694: res <= 0;
	2695: res <= 0;
	2696: res <= 0;
	2697: res <= 0;
	2698: res <= 0;
	2699: res <= 0;
	2700: res <= 0;
	2701: res <= 0;
	2702: res <= 0;
	2703: res <= 0;
	2704: res <= 0;
	2705: res <= 0;
	2706: res <= 0;
	2707: res <= 0;
	2708: res <= 0;
	2709: res <= 0;
	2710: res <= 0;
	2711: res <= 0;
	2712: res <= 0;
	2713: res <= 15;
	2714: res <= 3;
	2715: res <= 0;
	2716: res <= 0;
	2717: res <= 0;
	2718: res <= 0;
	2719: res <= 0;
	2720: res <= 15;
	2721: res <= 15;
	2722: res <= 15;
	2723: res <= 13;
	2724: res <= 15;
	2725: res <= 15;
	2726: res <= 15;
	2727: res <= 15;
	2728: res <= 7;
	2729: res <= 0;
	2730: res <= 0;
	2731: res <= 0;
	2732: res <= 0;
	2733: res <= 0;
	2734: res <= 0;
	2735: res <= 0;
	2736: res <= 12;
	2737: res <= 1;
	2738: res <= 7;
	2739: res <= 0;
	2740: res <= 0;
	2741: res <= 0;
	2742: res <= 0;
	2743: res <= 0;
	2744: res <= 0;
	2745: res <= 0;
	2746: res <= 0;
	2747: res <= 0;
	2748: res <= 0;
	2749: res <= 0;
	2750: res <= 0;
	2751: res <= 0;
	2752: res <= 0;
	2753: res <= 0;
	2754: res <= 0;
	2755: res <= 0;
	2756: res <= 0;
	2757: res <= 0;
	2758: res <= 15;
	2759: res <= 3;
	2760: res <= 0;
	2761: res <= 0;
	2762: res <= 0;
	2763: res <= 0;
	2764: res <= 0;
	2765: res <= 15;
	2766: res <= 15;
	2767: res <= 15;
	2768: res <= 14;
	2769: res <= 15;
	2770: res <= 15;
	2771: res <= 15;
	2772: res <= 15;
	2773: res <= 11;
	2774: res <= 1;
	2775: res <= 0;
	2776: res <= 0;
	2777: res <= 0;
	2778: res <= 0;
	2779: res <= 0;
	2780: res <= 0;
	2781: res <= 12;
	2782: res <= 15;
	2783: res <= 0;
	2784: res <= 0;
	2785: res <= 0;
	2786: res <= 0;
	2787: res <= 0;
	2788: res <= 0;
	2789: res <= 0;
	2790: res <= 0;
	2791: res <= 0;
	2792: res <= 0;
	2793: res <= 0;
	2794: res <= 0;
	2795: res <= 0;
	2796: res <= 0;
	2797: res <= 0;
	2798: res <= 0;
	2799: res <= 0;
	2800: res <= 0;
	2801: res <= 0;
	2802: res <= 0;
	2803: res <= 15;
	2804: res <= 3;
	2805: res <= 0;
	2806: res <= 0;
	2807: res <= 0;
	2808: res <= 0;
	2809: res <= 0;
	2810: res <= 15;
	2811: res <= 15;
	2812: res <= 7;
	2813: res <= 14;
	2814: res <= 15;
	2815: res <= 15;
	2816: res <= 15;
	2817: res <= 15;
	2818: res <= 11;
	2819: res <= 1;
	2820: res <= 0;
	2821: res <= 0;
	2822: res <= 0;
	2823: res <= 0;
	2824: res <= 0;
	2825: res <= 0;
	2826: res <= 12;
	2827: res <= 15;
	2828: res <= 0;
	2829: res <= 0;
	2830: res <= 0;
	2831: res <= 0;
	2832: res <= 0;
	2833: res <= 0;
	2834: res <= 0;
	2835: res <= 0;
	2836: res <= 0;
	2837: res <= 0;
	2838: res <= 0;
	2839: res <= 0;
	2840: res <= 0;
	2841: res <= 0;
	2842: res <= 0;
	2843: res <= 0;
	2844: res <= 0;
	2845: res <= 0;
	2846: res <= 0;
	2847: res <= 8;
	2848: res <= 15;
	2849: res <= 3;
	2850: res <= 0;
	2851: res <= 0;
	2852: res <= 0;
	2853: res <= 0;
	2854: res <= 8;
	2855: res <= 15;
	2856: res <= 15;
	2857: res <= 7;
	2858: res <= 15;
	2859: res <= 15;
	2860: res <= 15;
	2861: res <= 15;
	2862: res <= 15;
	2863: res <= 13;
	2864: res <= 1;
	2865: res <= 0;
	2866: res <= 0;
	2867: res <= 0;
	2868: res <= 0;
	2869: res <= 0;
	2870: res <= 0;
	2871: res <= 12;
	2872: res <= 15;
	2873: res <= 0;
	2874: res <= 0;
	2875: res <= 0;
	2876: res <= 0;
	2877: res <= 0;
	2878: res <= 0;
	2879: res <= 0;
	2880: res <= 0;
	2881: res <= 0;
	2882: res <= 0;
	2883: res <= 0;
	2884: res <= 7;
	2885: res <= 12;
	2886: res <= 1;
	2887: res <= 0;
	2888: res <= 0;
	2889: res <= 0;
	2890: res <= 0;
	2891: res <= 0;
	2892: res <= 8;
	2893: res <= 15;
	2894: res <= 3;
	2895: res <= 0;
	2896: res <= 0;
	2897: res <= 0;
	2898: res <= 0;
	2899: res <= 8;
	2900: res <= 15;
	2901: res <= 15;
	2902: res <= 11;
	2903: res <= 15;
	2904: res <= 15;
	2905: res <= 15;
	2906: res <= 15;
	2907: res <= 15;
	2908: res <= 14;
	2909: res <= 1;
	2910: res <= 0;
	2911: res <= 0;
	2912: res <= 0;
	2913: res <= 0;
	2914: res <= 0;
	2915: res <= 0;
	2916: res <= 0;
	2917: res <= 0;
	2918: res <= 0;
	2919: res <= 0;
	2920: res <= 0;
	2921: res <= 0;
	2922: res <= 0;
	2923: res <= 0;
	2924: res <= 0;
	2925: res <= 0;
	2926: res <= 0;
	2927: res <= 0;
	2928: res <= 0;
	2929: res <= 7;
	2930: res <= 12;
	2931: res <= 1;
	2932: res <= 0;
	2933: res <= 0;
	2934: res <= 0;
	2935: res <= 0;
	2936: res <= 0;
	2937: res <= 8;
	2938: res <= 15;
	2939: res <= 3;
	2940: res <= 0;
	2941: res <= 0;
	2942: res <= 0;
	2943: res <= 0;
	2944: res <= 8;
	2945: res <= 15;
	2946: res <= 15;
	2947: res <= 13;
	2948: res <= 15;
	2949: res <= 15;
	2950: res <= 15;
	2951: res <= 15;
	2952: res <= 7;
	2953: res <= 15;
	2954: res <= 1;
	2955: res <= 0;
	2956: res <= 0;
	2957: res <= 14;
	2958: res <= 0;
	2959: res <= 0;
	2960: res <= 0;
	2961: res <= 0;
	2962: res <= 0;
	2963: res <= 0;
	2964: res <= 0;
	2965: res <= 0;
	2966: res <= 0;
	2967: res <= 0;
	2968: res <= 0;
	2969: res <= 0;
	2970: res <= 0;
	2971: res <= 0;
	2972: res <= 0;
	2973: res <= 0;
	2974: res <= 7;
	2975: res <= 12;
	2976: res <= 1;
	2977: res <= 0;
	2978: res <= 0;
	2979: res <= 0;
	2980: res <= 0;
	2981: res <= 0;
	2982: res <= 8;
	2983: res <= 15;
	2984: res <= 3;
	2985: res <= 0;
	2986: res <= 0;
	2987: res <= 0;
	2988: res <= 0;
	2989: res <= 8;
	2990: res <= 15;
	2991: res <= 15;
	2992: res <= 15;
	2993: res <= 15;
	2994: res <= 15;
	2995: res <= 15;
	2996: res <= 15;
	2997: res <= 11;
	2998: res <= 15;
	2999: res <= 1;
	3000: res <= 0;
	3001: res <= 12;
	3002: res <= 15;
	3003: res <= 0;
	3004: res <= 0;
	3005: res <= 0;
	3006: res <= 0;
	3007: res <= 0;
	3008: res <= 0;
	3009: res <= 0;
	3010: res <= 0;
	3011: res <= 0;
	3012: res <= 0;
	3013: res <= 0;
	3014: res <= 0;
	3015: res <= 0;
	3016: res <= 0;
	3017: res <= 0;
	3018: res <= 0;
	3019: res <= 8;
	3020: res <= 3;
	3021: res <= 0;
	3022: res <= 0;
	3023: res <= 0;
	3024: res <= 0;
	3025: res <= 0;
	3026: res <= 0;
	3027: res <= 0;
	3028: res <= 15;
	3029: res <= 3;
	3030: res <= 0;
	3031: res <= 0;
	3032: res <= 0;
	3033: res <= 0;
	3034: res <= 12;
	3035: res <= 15;
	3036: res <= 15;
	3037: res <= 14;
	3038: res <= 15;
	3039: res <= 15;
	3040: res <= 15;
	3041: res <= 15;
	3042: res <= 13;
	3043: res <= 15;
	3044: res <= 0;
	3045: res <= 14;
	3046: res <= 15;
	3047: res <= 7;
	3048: res <= 0;
	3049: res <= 0;
	3050: res <= 0;
	3051: res <= 0;
	3052: res <= 0;
	3053: res <= 0;
	3054: res <= 0;
	3055: res <= 0;
	3056: res <= 0;
	3057: res <= 0;
	3058: res <= 0;
	3059: res <= 0;
	3060: res <= 0;
	3061: res <= 0;
	3062: res <= 0;
	3063: res <= 0;
	3064: res <= 8;
	3065: res <= 3;
	3066: res <= 0;
	3067: res <= 0;
	3068: res <= 0;
	3069: res <= 0;
	3070: res <= 0;
	3071: res <= 0;
	3072: res <= 0;
	3073: res <= 15;
	3074: res <= 3;
	3075: res <= 0;
	3076: res <= 0;
	3077: res <= 0;
	3078: res <= 0;
	3079: res <= 12;
	3080: res <= 15;
	3081: res <= 7;
	3082: res <= 15;
	3083: res <= 15;
	3084: res <= 15;
	3085: res <= 15;
	3086: res <= 15;
	3087: res <= 13;
	3088: res <= 3;
	3089: res <= 12;
	3090: res <= 15;
	3091: res <= 15;
	3092: res <= 7;
	3093: res <= 0;
	3094: res <= 0;
	3095: res <= 0;
	3096: res <= 0;
	3097: res <= 7;
	3098: res <= 0;
	3099: res <= 0;
	3100: res <= 0;
	3101: res <= 0;
	3102: res <= 0;
	3103: res <= 0;
	3104: res <= 0;
	3105: res <= 0;
	3106: res <= 0;
	3107: res <= 0;
	3108: res <= 0;
	3109: res <= 8;
	3110: res <= 3;
	3111: res <= 0;
	3112: res <= 0;
	3113: res <= 0;
	3114: res <= 0;
	3115: res <= 0;
	3116: res <= 0;
	3117: res <= 0;
	3118: res <= 15;
	3119: res <= 3;
	3120: res <= 0;
	3121: res <= 0;
	3122: res <= 0;
	3123: res <= 0;
	3124: res <= 12;
	3125: res <= 15;
	3126: res <= 11;
	3127: res <= 15;
	3128: res <= 15;
	3129: res <= 15;
	3130: res <= 15;
	3131: res <= 15;
	3132: res <= 0;
	3133: res <= 8;
	3134: res <= 15;
	3135: res <= 15;
	3136: res <= 15;
	3137: res <= 3;
	3138: res <= 0;
	3139: res <= 0;
	3140: res <= 0;
	3141: res <= 0;
	3142: res <= 7;
	3143: res <= 0;
	3144: res <= 0;
	3145: res <= 0;
	3146: res <= 0;
	3147: res <= 0;
	3148: res <= 0;
	3149: res <= 0;
	3150: res <= 0;
	3151: res <= 0;
	3152: res <= 0;
	3153: res <= 0;
	3154: res <= 7;
	3155: res <= 12;
	3156: res <= 1;
	3157: res <= 0;
	3158: res <= 0;
	3159: res <= 0;
	3160: res <= 0;
	3161: res <= 0;
	3162: res <= 0;
	3163: res <= 15;
	3164: res <= 3;
	3165: res <= 0;
	3166: res <= 0;
	3167: res <= 0;
	3168: res <= 0;
	3169: res <= 12;
	3170: res <= 15;
	3171: res <= 15;
	3172: res <= 15;
	3173: res <= 15;
	3174: res <= 15;
	3175: res <= 15;
	3176: res <= 3;
	3177: res <= 0;
	3178: res <= 15;
	3179: res <= 15;
	3180: res <= 15;
	3181: res <= 15;
	3182: res <= 1;
	3183: res <= 0;
	3184: res <= 0;
	3185: res <= 0;
	3186: res <= 0;
	3187: res <= 7;
	3188: res <= 0;
	3189: res <= 0;
	3190: res <= 0;
	3191: res <= 0;
	3192: res <= 0;
	3193: res <= 0;
	3194: res <= 0;
	3195: res <= 0;
	3196: res <= 0;
	3197: res <= 0;
	3198: res <= 0;
	3199: res <= 7;
	3200: res <= 12;
	3201: res <= 1;
	3202: res <= 0;
	3203: res <= 0;
	3204: res <= 0;
	3205: res <= 0;
	3206: res <= 0;
	3207: res <= 0;
	3208: res <= 15;
	3209: res <= 3;
	3210: res <= 0;
	3211: res <= 0;
	3212: res <= 0;
	3213: res <= 0;
	3214: res <= 14;
	3215: res <= 15;
	3216: res <= 13;
	3217: res <= 15;
	3218: res <= 15;
	3219: res <= 15;
	3220: res <= 15;
	3221: res <= 0;
	3222: res <= 14;
	3223: res <= 15;
	3224: res <= 15;
	3225: res <= 15;
	3226: res <= 15;
	3227: res <= 1;
	3228: res <= 0;
	3229: res <= 0;
	3230: res <= 0;
	3231: res <= 14;
	3232: res <= 8;
	3233: res <= 3;
	3234: res <= 0;
	3235: res <= 0;
	3236: res <= 0;
	3237: res <= 0;
	3238: res <= 0;
	3239: res <= 0;
	3240: res <= 0;
	3241: res <= 0;
	3242: res <= 0;
	3243: res <= 0;
	3244: res <= 7;
	3245: res <= 12;
	3246: res <= 1;
	3247: res <= 0;
	3248: res <= 0;
	3249: res <= 0;
	3250: res <= 0;
	3251: res <= 0;
	3252: res <= 0;
	3253: res <= 14;
	3254: res <= 7;
	3255: res <= 0;
	3256: res <= 0;
	3257: res <= 0;
	3258: res <= 0;
	3259: res <= 14;
	3260: res <= 15;
	3261: res <= 14;
	3262: res <= 15;
	3263: res <= 15;
	3264: res <= 15;
	3265: res <= 3;
	3266: res <= 12;
	3267: res <= 15;
	3268: res <= 15;
	3269: res <= 15;
	3270: res <= 15;
	3271: res <= 15;
	3272: res <= 0;
	3273: res <= 0;
	3274: res <= 0;
	3275: res <= 0;
	3276: res <= 14;
	3277: res <= 8;
	3278: res <= 3;
	3279: res <= 0;
	3280: res <= 0;
	3281: res <= 0;
	3282: res <= 0;
	3283: res <= 0;
	3284: res <= 0;
	3285: res <= 0;
	3286: res <= 0;
	3287: res <= 0;
	3288: res <= 0;
	3289: res <= 0;
	3290: res <= 0;
	3291: res <= 0;
	3292: res <= 0;
	3293: res <= 0;
	3294: res <= 0;
	3295: res <= 0;
	3296: res <= 0;
	3297: res <= 0;
	3298: res <= 14;
	3299: res <= 7;
	3300: res <= 0;
	3301: res <= 0;
	3302: res <= 0;
	3303: res <= 0;
	3304: res <= 15;
	3305: res <= 15;
	3306: res <= 14;
	3307: res <= 15;
	3308: res <= 15;
	3309: res <= 15;
	3310: res <= 8;
	3311: res <= 15;
	3312: res <= 15;
	3313: res <= 15;
	3314: res <= 15;
	3315: res <= 15;
	3316: res <= 3;
	3317: res <= 0;
	3318: res <= 0;
	3319: res <= 0;
	3320: res <= 0;
	3321: res <= 14;
	3322: res <= 8;
	3323: res <= 3;
	3324: res <= 0;
	3325: res <= 0;
	3326: res <= 0;
	3327: res <= 0;
	3328: res <= 0;
	3329: res <= 0;
	3330: res <= 0;
	3331: res <= 0;
	3332: res <= 0;
	3333: res <= 0;
	3334: res <= 0;
	3335: res <= 0;
	3336: res <= 0;
	3337: res <= 0;
	3338: res <= 0;
	3339: res <= 0;
	3340: res <= 0;
	3341: res <= 0;
	3342: res <= 0;
	3343: res <= 14;
	3344: res <= 7;
	3345: res <= 0;
	3346: res <= 0;
	3347: res <= 0;
	3348: res <= 0;
	3349: res <= 15;
	3350: res <= 7;
	3351: res <= 15;
	3352: res <= 15;
	3353: res <= 15;
	3354: res <= 3;
	3355: res <= 14;
	3356: res <= 15;
	3357: res <= 15;
	3358: res <= 15;
	3359: res <= 15;
	3360: res <= 15;
	3361: res <= 1;
	3362: res <= 0;
	3363: res <= 0;
	3364: res <= 0;
	3365: res <= 0;
	3366: res <= 14;
	3367: res <= 8;
	3368: res <= 3;
	3369: res <= 0;
	3370: res <= 0;
	3371: res <= 0;
	3372: res <= 0;
	3373: res <= 0;
	3374: res <= 0;
	3375: res <= 0;
	3376: res <= 0;
	3377: res <= 0;
	3378: res <= 0;
	3379: res <= 0;
	3380: res <= 0;
	3381: res <= 0;
	3382: res <= 0;
	3383: res <= 0;
	3384: res <= 0;
	3385: res <= 0;
	3386: res <= 0;
	3387: res <= 0;
	3388: res <= 14;
	3389: res <= 7;
	3390: res <= 0;
	3391: res <= 0;
	3392: res <= 0;
	3393: res <= 0;
	3394: res <= 15;
	3395: res <= 11;
	3396: res <= 15;
	3397: res <= 15;
	3398: res <= 15;
	3399: res <= 9;
	3400: res <= 15;
	3401: res <= 15;
	3402: res <= 15;
	3403: res <= 15;
	3404: res <= 15;
	3405: res <= 15;
	3406: res <= 0;
	3407: res <= 0;
	3408: res <= 0;
	3409: res <= 0;
	3410: res <= 0;
	3411: res <= 14;
	3412: res <= 8;
	3413: res <= 3;
	3414: res <= 0;
	3415: res <= 0;
	3416: res <= 0;
	3417: res <= 0;
	3418: res <= 0;
	3419: res <= 0;
	3420: res <= 0;
	3421: res <= 0;
	3422: res <= 0;
	3423: res <= 0;
	3424: res <= 2;
	3425: res <= 8;
	3426: res <= 0;
	3427: res <= 0;
	3428: res <= 0;
	3429: res <= 0;
	3430: res <= 0;
	3431: res <= 0;
	3432: res <= 0;
	3433: res <= 12;
	3434: res <= 15;
	3435: res <= 0;
	3436: res <= 0;
	3437: res <= 0;
	3438: res <= 0;
	3439: res <= 15;
	3440: res <= 11;
	3441: res <= 15;
	3442: res <= 15;
	3443: res <= 7;
	3444: res <= 12;
	3445: res <= 15;
	3446: res <= 15;
	3447: res <= 15;
	3448: res <= 15;
	3449: res <= 15;
	3450: res <= 3;
	3451: res <= 0;
	3452: res <= 0;
	3453: res <= 0;
	3454: res <= 0;
	3455: res <= 0;
	3456: res <= 14;
	3457: res <= 8;
	3458: res <= 3;
	3459: res <= 0;
	3460: res <= 0;
	3461: res <= 0;
	3462: res <= 0;
	3463: res <= 0;
	3464: res <= 0;
	3465: res <= 0;
	3466: res <= 0;
	3467: res <= 0;
	3468: res <= 0;
	3469: res <= 4;
	3470: res <= 4;
	3471: res <= 0;
	3472: res <= 0;
	3473: res <= 4;
	3474: res <= 5;
	3475: res <= 1;
	3476: res <= 0;
	3477: res <= 0;
	3478: res <= 12;
	3479: res <= 15;
	3480: res <= 1;
	3481: res <= 0;
	3482: res <= 0;
	3483: res <= 8;
	3484: res <= 15;
	3485: res <= 13;
	3486: res <= 15;
	3487: res <= 15;
	3488: res <= 1;
	3489: res <= 15;
	3490: res <= 15;
	3491: res <= 15;
	3492: res <= 15;
	3493: res <= 15;
	3494: res <= 15;
	3495: res <= 1;
	3496: res <= 0;
	3497: res <= 0;
	3498: res <= 0;
	3499: res <= 0;
	3500: res <= 0;
	3501: res <= 0;
	3502: res <= 7;
	3503: res <= 0;
	3504: res <= 0;
	3505: res <= 0;
	3506: res <= 0;
	3507: res <= 0;
	3508: res <= 0;
	3509: res <= 0;
	3510: res <= 0;
	3511: res <= 0;
	3512: res <= 0;
	3513: res <= 0;
	3514: res <= 8;
	3515: res <= 2;
	3516: res <= 0;
	3517: res <= 0;
	3518: res <= 8;
	3519: res <= 10;
	3520: res <= 0;
	3521: res <= 0;
	3522: res <= 0;
	3523: res <= 12;
	3524: res <= 15;
	3525: res <= 1;
	3526: res <= 0;
	3527: res <= 0;
	3528: res <= 8;
	3529: res <= 15;
	3530: res <= 12;
	3531: res <= 15;
	3532: res <= 15;
	3533: res <= 12;
	3534: res <= 15;
	3535: res <= 15;
	3536: res <= 15;
	3537: res <= 15;
	3538: res <= 15;
	3539: res <= 7;
	3540: res <= 0;
	3541: res <= 0;
	3542: res <= 0;
	3543: res <= 0;
	3544: res <= 0;
	3545: res <= 0;
	3546: res <= 0;
	3547: res <= 7;
	3548: res <= 0;
	3549: res <= 0;
	3550: res <= 0;
	3551: res <= 0;
	3552: res <= 0;
	3553: res <= 0;
	3554: res <= 0;
	3555: res <= 0;
	3556: res <= 0;
	3557: res <= 0;
	3558: res <= 0;
	3559: res <= 0;
	3560: res <= 1;
	3561: res <= 0;
	3562: res <= 0;
	3563: res <= 4;
	3564: res <= 5;
	3565: res <= 1;
	3566: res <= 0;
	3567: res <= 0;
	3568: res <= 8;
	3569: res <= 15;
	3570: res <= 3;
	3571: res <= 0;
	3572: res <= 0;
	3573: res <= 8;
	3574: res <= 15;
	3575: res <= 14;
	3576: res <= 15;
	3577: res <= 3;
	3578: res <= 14;
	3579: res <= 15;
	3580: res <= 15;
	3581: res <= 15;
	3582: res <= 15;
	3583: res <= 15;
	3584: res <= 3;
	3585: res <= 0;
	3586: res <= 0;
	3587: res <= 0;
	3588: res <= 0;
	3589: res <= 0;
	3590: res <= 0;
	3591: res <= 0;
	3592: res <= 7;
	3593: res <= 0;
	3594: res <= 0;
	3595: res <= 0;
	3596: res <= 0;
	3597: res <= 0;
	3598: res <= 0;
	3599: res <= 0;
	3600: res <= 0;
	3601: res <= 0;
	3602: res <= 0;
	3603: res <= 0;
	3604: res <= 8;
	3605: res <= 2;
	3606: res <= 0;
	3607: res <= 0;
	3608: res <= 8;
	3609: res <= 10;
	3610: res <= 0;
	3611: res <= 0;
	3612: res <= 0;
	3613: res <= 8;
	3614: res <= 15;
	3615: res <= 3;
	3616: res <= 0;
	3617: res <= 0;
	3618: res <= 8;
	3619: res <= 7;
	3620: res <= 15;
	3621: res <= 15;
	3622: res <= 1;
	3623: res <= 15;
	3624: res <= 15;
	3625: res <= 15;
	3626: res <= 15;
	3627: res <= 15;
	3628: res <= 15;
	3629: res <= 0;
	3630: res <= 0;
	3631: res <= 0;
	3632: res <= 0;
	3633: res <= 0;
	3634: res <= 0;
	3635: res <= 0;
	3636: res <= 0;
	3637: res <= 0;
	3638: res <= 0;
	3639: res <= 0;
	3640: res <= 0;
	3641: res <= 0;
	3642: res <= 0;
	3643: res <= 0;
	3644: res <= 0;
	3645: res <= 0;
	3646: res <= 0;
	3647: res <= 0;
	3648: res <= 0;
	3649: res <= 4;
	3650: res <= 4;
	3651: res <= 0;
	3652: res <= 0;
	3653: res <= 4;
	3654: res <= 5;
	3655: res <= 1;
	3656: res <= 0;
	3657: res <= 0;
	3658: res <= 0;
	3659: res <= 15;
	3660: res <= 7;
	3661: res <= 0;
	3662: res <= 0;
	3663: res <= 8;
	3664: res <= 7;
	3665: res <= 15;
	3666: res <= 7;
	3667: res <= 12;
	3668: res <= 15;
	3669: res <= 15;
	3670: res <= 15;
	3671: res <= 15;
	3672: res <= 15;
	3673: res <= 7;
	3674: res <= 0;
	3675: res <= 0;
	3676: res <= 0;
	3677: res <= 0;
	3678: res <= 0;
	3679: res <= 0;
	3680: res <= 0;
	3681: res <= 0;
	3682: res <= 0;
	3683: res <= 0;
	3684: res <= 0;
	3685: res <= 0;
	3686: res <= 0;
	3687: res <= 0;
	3688: res <= 0;
	3689: res <= 0;
	3690: res <= 0;
	3691: res <= 0;
	3692: res <= 0;
	3693: res <= 0;
	3694: res <= 2;
	3695: res <= 8;
	3696: res <= 0;
	3697: res <= 0;
	3698: res <= 8;
	3699: res <= 10;
	3700: res <= 0;
	3701: res <= 0;
	3702: res <= 0;
	3703: res <= 0;
	3704: res <= 14;
	3705: res <= 15;
	3706: res <= 0;
	3707: res <= 0;
	3708: res <= 12;
	3709: res <= 11;
	3710: res <= 15;
	3711: res <= 3;
	3712: res <= 15;
	3713: res <= 15;
	3714: res <= 15;
	3715: res <= 15;
	3716: res <= 15;
	3717: res <= 15;
	3718: res <= 1;
	3719: res <= 0;
	3720: res <= 0;
	3721: res <= 0;
	3722: res <= 0;
	3723: res <= 0;
	3724: res <= 0;
	3725: res <= 0;
	3726: res <= 0;
	3727: res <= 0;
	3728: res <= 0;
	3729: res <= 0;
	3730: res <= 0;
	3731: res <= 0;
	3732: res <= 0;
	3733: res <= 0;
	3734: res <= 0;
	3735: res <= 0;
	3736: res <= 0;
	3737: res <= 0;
	3738: res <= 0;
	3739: res <= 0;
	3740: res <= 0;
	3741: res <= 0;
	3742: res <= 0;
	3743: res <= 4;
	3744: res <= 5;
	3745: res <= 1;
	3746: res <= 0;
	3747: res <= 0;
	3748: res <= 0;
	3749: res <= 14;
	3750: res <= 15;
	3751: res <= 1;
	3752: res <= 0;
	3753: res <= 12;
	3754: res <= 11;
	3755: res <= 15;
	3756: res <= 8;
	3757: res <= 15;
	3758: res <= 15;
	3759: res <= 15;
	3760: res <= 15;
	3761: res <= 15;
	3762: res <= 7;
	3763: res <= 0;
	3764: res <= 0;
	3765: res <= 0;
	3766: res <= 0;
	3767: res <= 0;
	3768: res <= 0;
	3769: res <= 0;
	3770: res <= 0;
	3771: res <= 0;
	3772: res <= 15;
	3773: res <= 3;
	3774: res <= 0;
	3775: res <= 0;
	3776: res <= 0;
	3777: res <= 0;
	3778: res <= 0;
	3779: res <= 0;
	3780: res <= 0;
	3781: res <= 0;
	3782: res <= 0;
	3783: res <= 0;
	3784: res <= 0;
	3785: res <= 0;
	3786: res <= 0;
	3787: res <= 0;
	3788: res <= 0;
	3789: res <= 0;
	3790: res <= 0;
	3791: res <= 0;
	3792: res <= 0;
	3793: res <= 0;
	3794: res <= 12;
	3795: res <= 15;
	3796: res <= 3;
	3797: res <= 0;
	3798: res <= 12;
	3799: res <= 13;
	3800: res <= 7;
	3801: res <= 12;
	3802: res <= 15;
	3803: res <= 15;
	3804: res <= 15;
	3805: res <= 15;
	3806: res <= 15;
	3807: res <= 1;
	3808: res <= 0;
	3809: res <= 0;
	3810: res <= 0;
	3811: res <= 0;
	3812: res <= 0;
	3813: res <= 0;
	3814: res <= 0;
	3815: res <= 0;
	3816: res <= 0;
	3817: res <= 15;
	3818: res <= 3;
	3819: res <= 0;
	3820: res <= 0;
	3821: res <= 0;
	3822: res <= 0;
	3823: res <= 0;
	3824: res <= 0;
	3825: res <= 0;
	3826: res <= 0;
	3827: res <= 0;
	3828: res <= 0;
	3829: res <= 0;
	3830: res <= 0;
	3831: res <= 0;
	3832: res <= 0;
	3833: res <= 0;
	3834: res <= 0;
	3835: res <= 0;
	3836: res <= 0;
	3837: res <= 0;
	3838: res <= 0;
	3839: res <= 8;
	3840: res <= 15;
	3841: res <= 7;
	3842: res <= 0;
	3843: res <= 12;
	3844: res <= 13;
	3845: res <= 3;
	3846: res <= 15;
	3847: res <= 15;
	3848: res <= 15;
	3849: res <= 15;
	3850: res <= 15;
	3851: res <= 7;
	3852: res <= 0;
	3853: res <= 0;
	3854: res <= 0;
	3855: res <= 0;
	3856: res <= 0;
	3857: res <= 0;
	3858: res <= 0;
	3859: res <= 0;
	3860: res <= 0;
	3861: res <= 0;
	3862: res <= 15;
	3863: res <= 3;
	3864: res <= 0;
	3865: res <= 0;
	3866: res <= 0;
	3867: res <= 0;
	3868: res <= 0;
	3869: res <= 0;
	3870: res <= 0;
	3871: res <= 0;
	3872: res <= 0;
	3873: res <= 0;
	3874: res <= 0;
	3875: res <= 0;
	3876: res <= 0;
	3877: res <= 0;
	3878: res <= 0;
	3879: res <= 0;
	3880: res <= 0;
	3881: res <= 0;
	3882: res <= 0;
	3883: res <= 0;
	3884: res <= 0;
	3885: res <= 15;
	3886: res <= 15;
	3887: res <= 0;
	3888: res <= 12;
	3889: res <= 14;
	3890: res <= 13;
	3891: res <= 15;
	3892: res <= 15;
	3893: res <= 15;
	3894: res <= 15;
	3895: res <= 15;
	3896: res <= 1;
	3897: res <= 0;
	3898: res <= 0;
	3899: res <= 0;
	3900: res <= 0;
	3901: res <= 0;
	3902: res <= 0;
	3903: res <= 0;
	3904: res <= 0;
	3905: res <= 0;
	3906: res <= 14;
	3907: res <= 0;
	3908: res <= 0;
	3909: res <= 0;
	3910: res <= 0;
	3911: res <= 0;
	3912: res <= 0;
	3913: res <= 0;
	3914: res <= 0;
	3915: res <= 0;
	3916: res <= 0;
	3917: res <= 0;
	3918: res <= 0;
	3919: res <= 5;
	3920: res <= 5;
	3921: res <= 0;
	3922: res <= 0;
	3923: res <= 14;
	3924: res <= 15;
	3925: res <= 0;
	3926: res <= 0;
	3927: res <= 0;
	3928: res <= 0;
	3929: res <= 0;
	3930: res <= 14;
	3931: res <= 15;
	3932: res <= 3;
	3933: res <= 14;
	3934: res <= 6;
	3935: res <= 14;
	3936: res <= 15;
	3937: res <= 15;
	3938: res <= 15;
	3939: res <= 15;
	3940: res <= 3;
	3941: res <= 6;
	3942: res <= 0;
	3943: res <= 0;
	3944: res <= 0;
	3945: res <= 0;
	3946: res <= 0;
	3947: res <= 0;
	3948: res <= 0;
	3949: res <= 0;
	3950: res <= 0;
	3951: res <= 14;
	3952: res <= 0;
	3953: res <= 0;
	3954: res <= 0;
	3955: res <= 0;
	3956: res <= 0;
	3957: res <= 0;
	3958: res <= 0;
	3959: res <= 0;
	3960: res <= 0;
	3961: res <= 0;
	3962: res <= 0;
	3963: res <= 0;
	3964: res <= 5;
	3965: res <= 5;
	3966: res <= 0;
	3967: res <= 0;
	3968: res <= 0;
	3969: res <= 0;
	3970: res <= 0;
	3971: res <= 0;
	3972: res <= 0;
	3973: res <= 0;
	3974: res <= 0;
	3975: res <= 12;
	3976: res <= 15;
	3977: res <= 7;
	3978: res <= 6;
	3979: res <= 3;
	3980: res <= 15;
	3981: res <= 15;
	3982: res <= 15;
	3983: res <= 15;
	3984: res <= 15;
	3985: res <= 12;
	3986: res <= 3;
	3987: res <= 0;
	3988: res <= 0;
	3989: res <= 0;
	3990: res <= 0;
	3991: res <= 0;
	3992: res <= 0;
	3993: res <= 0;
	3994: res <= 0;
	3995: res <= 0;
	3996: res <= 14;
	3997: res <= 0;
	3998: res <= 0;
	3999: res <= 0;
	4000: res <= 0;
	4001: res <= 0;
	4002: res <= 0;
	4003: res <= 0;
	4004: res <= 0;
	4005: res <= 0;
	4006: res <= 0;
	4007: res <= 0;
	4008: res <= 0;
	4009: res <= 5;
	4010: res <= 5;
	4011: res <= 0;
	4012: res <= 0;
	4013: res <= 14;
	4014: res <= 15;
	4015: res <= 0;
	4016: res <= 0;
	4017: res <= 0;
	4018: res <= 0;
	4019: res <= 0;
	4020: res <= 8;
	4021: res <= 15;
	4022: res <= 15;
	4023: res <= 6;
	4024: res <= 12;
	4025: res <= 15;
	4026: res <= 15;
	4027: res <= 15;
	4028: res <= 15;
	4029: res <= 9;
	4030: res <= 15;
	4031: res <= 1;
	4032: res <= 0;
	4033: res <= 0;
	4034: res <= 0;
	4035: res <= 0;
	4036: res <= 0;
	4037: res <= 0;
	4038: res <= 0;
	4039: res <= 0;
	4040: res <= 0;
	4041: res <= 14;
	4042: res <= 0;
	4043: res <= 0;
	4044: res <= 0;
	4045: res <= 0;
	4046: res <= 0;
	4047: res <= 0;
	4048: res <= 0;
	4049: res <= 0;
	4050: res <= 0;
	4051: res <= 0;
	4052: res <= 0;
	4053: res <= 0;
	4054: res <= 5;
	4055: res <= 5;
	4056: res <= 0;
	4057: res <= 0;
	4058: res <= 0;
	4059: res <= 0;
	4060: res <= 0;
	4061: res <= 0;
	4062: res <= 0;
	4063: res <= 0;
	4064: res <= 0;
	4065: res <= 0;
	4066: res <= 15;
	4067: res <= 7;
	4068: res <= 2;
	4069: res <= 14;
	4070: res <= 3;
	4071: res <= 0;
	4072: res <= 0;
	4073: res <= 15;
	4074: res <= 15;
	4075: res <= 15;
	4076: res <= 0;
	4077: res <= 0;
	4078: res <= 0;
	4079: res <= 0;
	4080: res <= 0;
	4081: res <= 0;
	4082: res <= 0;
	4083: res <= 0;
	4084: res <= 0;
	4085: res <= 0;
	4086: res <= 14;
	4087: res <= 0;
	4088: res <= 0;
	4089: res <= 0;
	4090: res <= 0;
	4091: res <= 0;
	4092: res <= 0;
	4093: res <= 0;
	4094: res <= 0;
	4095: res <= 0;
	4096: res <= 0;
	4097: res <= 0;
	4098: res <= 0;
	4099: res <= 5;
	4100: res <= 5;
	4101: res <= 0;
	4102: res <= 0;
	4103: res <= 14;
	4104: res <= 15;
	4105: res <= 0;
	4106: res <= 0;
	4107: res <= 0;
	4108: res <= 0;
	4109: res <= 0;
	4110: res <= 0;
	4111: res <= 14;
	4112: res <= 7;
	4113: res <= 3;
	4114: res <= 15;
	4115: res <= 0;
	4116: res <= 0;
	4117: res <= 15;
	4118: res <= 15;
	4119: res <= 15;
	4120: res <= 7;
	4121: res <= 0;
	4122: res <= 0;
	4123: res <= 0;
	4124: res <= 0;
	4125: res <= 0;
	4126: res <= 0;
	4127: res <= 0;
	4128: res <= 0;
	4129: res <= 0;
	4130: res <= 0;
	4131: res <= 14;
	4132: res <= 0;
	4133: res <= 0;
	4134: res <= 0;
	4135: res <= 0;
	4136: res <= 0;
	4137: res <= 0;
	4138: res <= 0;
	4139: res <= 0;
	4140: res <= 0;
	4141: res <= 0;
	4142: res <= 0;
	4143: res <= 0;
	4144: res <= 5;
	4145: res <= 5;
	4146: res <= 0;
	4147: res <= 0;
	4148: res <= 0;
	4149: res <= 0;
	4150: res <= 0;
	4151: res <= 0;
	4152: res <= 0;
	4153: res <= 0;
	4154: res <= 0;
	4155: res <= 0;
	4156: res <= 8;
	4157: res <= 7;
	4158: res <= 8;
	4159: res <= 3;
	4160: res <= 15;
	4161: res <= 15;
	4162: res <= 15;
	4163: res <= 15;
	4164: res <= 15;
	4165: res <= 1;
	4166: res <= 0;
	4167: res <= 0;
	4168: res <= 0;
	4169: res <= 0;
	4170: res <= 0;
	4171: res <= 0;
	4172: res <= 0;
	4173: res <= 0;
	4174: res <= 0;
	4175: res <= 0;
	4176: res <= 14;
	4177: res <= 0;
	4178: res <= 0;
	4179: res <= 0;
	4180: res <= 0;
	4181: res <= 0;
	4182: res <= 0;
	4183: res <= 0;
	4184: res <= 0;
	4185: res <= 0;
	4186: res <= 0;
	4187: res <= 0;
	4188: res <= 0;
	4189: res <= 0;
	4190: res <= 0;
	4191: res <= 0;
	4192: res <= 0;
	4193: res <= 14;
	4194: res <= 15;
	4195: res <= 0;
	4196: res <= 0;
	4197: res <= 0;
	4198: res <= 0;
	4199: res <= 0;
	4200: res <= 0;
	4201: res <= 0;
	4202: res <= 7;
	4203: res <= 12;
	4204: res <= 9;
	4205: res <= 15;
	4206: res <= 15;
	4207: res <= 15;
	4208: res <= 15;
	4209: res <= 15;
	4210: res <= 0;
	4211: res <= 0;
	4212: res <= 0;
	4213: res <= 0;
	4214: res <= 0;
	4215: res <= 0;
	4216: res <= 0;
	4217: res <= 0;
	4218: res <= 0;
	4219: res <= 0;
	4220: res <= 0;
	4221: res <= 14;
	4222: res <= 0;
	4223: res <= 0;
	4224: res <= 0;
	4225: res <= 0;
	4226: res <= 0;
	4227: res <= 0;
	4228: res <= 0;
	4229: res <= 0;
	4230: res <= 0;
	4231: res <= 0;
	4232: res <= 0;
	4233: res <= 0;
	4234: res <= 0;
	4235: res <= 0;
	4236: res <= 0;
	4237: res <= 0;
	4238: res <= 0;
	4239: res <= 0;
	4240: res <= 0;
	4241: res <= 0;
	4242: res <= 0;
	4243: res <= 0;
	4244: res <= 0;
	4245: res <= 0;
	4246: res <= 0;
	4247: res <= 0;
	4248: res <= 12;
	4249: res <= 14;
	4250: res <= 15;
	4251: res <= 15;
	4252: res <= 15;
	4253: res <= 15;
	4254: res <= 3;
	4255: res <= 0;
	4256: res <= 0;
	4257: res <= 0;
	4258: res <= 0;
	4259: res <= 0;
	4260: res <= 0;
	4261: res <= 0;
	4262: res <= 0;
	4263: res <= 0;
	4264: res <= 0;
	4265: res <= 0;
	4266: res <= 14;
	4267: res <= 0;
	4268: res <= 0;
	4269: res <= 0;
	4270: res <= 0;
	4271: res <= 0;
	4272: res <= 0;
	4273: res <= 0;
	4274: res <= 0;
	4275: res <= 0;
	4276: res <= 0;
	4277: res <= 0;
	4278: res <= 0;
	4279: res <= 0;
	4280: res <= 0;
	4281: res <= 0;
	4282: res <= 0;
	4283: res <= 0;
	4284: res <= 0;
	4285: res <= 0;
	4286: res <= 0;
	4287: res <= 0;
	4288: res <= 0;
	4289: res <= 0;
	4290: res <= 0;
	4291: res <= 0;
	4292: res <= 0;
	4293: res <= 0;
	4294: res <= 15;
	4295: res <= 15;
	4296: res <= 15;
	4297: res <= 15;
	4298: res <= 15;
	4299: res <= 0;
	4300: res <= 0;
	4301: res <= 0;
	4302: res <= 0;
	4303: res <= 0;
	4304: res <= 0;
	4305: res <= 0;
	4306: res <= 0;
	4307: res <= 0;
	4308: res <= 0;
	4309: res <= 0;
	4310: res <= 0;
	4311: res <= 0;
	4312: res <= 15;
	4313: res <= 3;
	4314: res <= 0;
	4315: res <= 0;
	4316: res <= 0;
	4317: res <= 0;
	4318: res <= 0;
	4319: res <= 0;
	4320: res <= 0;
	4321: res <= 0;
	4322: res <= 0;
	4323: res <= 0;
	4324: res <= 0;
	4325: res <= 0;
	4326: res <= 0;
	4327: res <= 0;
	4328: res <= 0;
	4329: res <= 0;
	4330: res <= 0;
	4331: res <= 0;
	4332: res <= 0;
	4333: res <= 0;
	4334: res <= 0;
	4335: res <= 0;
	4336: res <= 0;
	4337: res <= 0;
	4338: res <= 0;
	4339: res <= 15;
	4340: res <= 15;
	4341: res <= 15;
	4342: res <= 15;
	4343: res <= 0;
	4344: res <= 0;
	4345: res <= 0;
	4346: res <= 0;
	4347: res <= 0;
	4348: res <= 0;
	4349: res <= 0;
	4350: res <= 0;
	4351: res <= 0;
	4352: res <= 0;
	4353: res <= 0;
	4354: res <= 0;
	4355: res <= 0;
	4356: res <= 0;
	4357: res <= 15;
	4358: res <= 3;
	4359: res <= 0;
	4360: res <= 0;
	4361: res <= 0;
	4362: res <= 0;
	4363: res <= 0;
	4364: res <= 0;
	4365: res <= 0;
	4366: res <= 0;
	4367: res <= 0;
	4368: res <= 0;
	4369: res <= 0;
	4370: res <= 0;
	4371: res <= 0;
	4372: res <= 0;
	4373: res <= 0;
	4374: res <= 0;
	4375: res <= 0;
	4376: res <= 0;
	4377: res <= 0;
	4378: res <= 0;
	4379: res <= 0;
	4380: res <= 0;
	4381: res <= 0;
	4382: res <= 0;
	4383: res <= 0;
	4384: res <= 0;
	4385: res <= 0;
	4386: res <= 0;
	4387: res <= 0;
	4388: res <= 0;
	4389: res <= 0;
	4390: res <= 0;
	4391: res <= 0;
	4392: res <= 0;
	4393: res <= 0;
	4394: res <= 0;
	4395: res <= 0;
	4396: res <= 0;
	4397: res <= 0;
	4398: res <= 0;
	4399: res <= 0;
	4400: res <= 0;
	4401: res <= 0;
	4402: res <= 15;
	4403: res <= 3;
	4404: res <= 0;
	4405: res <= 0;
	4406: res <= 0;
	4407: res <= 0;
	4408: res <= 0;
	4409: res <= 0;
	4410: res <= 0;
	4411: res <= 0;
	4412: res <= 0;
	4413: res <= 0;
	4414: res <= 0;
	4415: res <= 0;
	4416: res <= 0;
	4417: res <= 0;
	4418: res <= 0;
	4419: res <= 0;
	4420: res <= 0;
	4421: res <= 0;
	4422: res <= 0;
	4423: res <= 0;
	4424: res <= 0;
	4425: res <= 0;
	4426: res <= 0;
	4427: res <= 0;
	4428: res <= 0;
	4429: res <= 0;
	4430: res <= 0;
	4431: res <= 0;
	4432: res <= 0;
	4433: res <= 0;
	4434: res <= 0;
	4435: res <= 0;
	4436: res <= 0;
	4437: res <= 0;
	4438: res <= 0;
	4439: res <= 0;
	4440: res <= 0;
	4441: res <= 0;
	4442: res <= 0;
	4443: res <= 0;
	4444: res <= 0;
	4445: res <= 0;
	4446: res <= 0;
	4447: res <= 0;
	4448: res <= 0;
	4449: res <= 0;
	4450: res <= 0;
	4451: res <= 0;
	4452: res <= 0;
	4453: res <= 0;
	4454: res <= 0;
	4455: res <= 0;
	4456: res <= 0;
	4457: res <= 0;
	4458: res <= 0;
	4459: res <= 0;
	4460: res <= 0;
	4461: res <= 0;
	4462: res <= 0;
	4463: res <= 0;
	4464: res <= 0;
	4465: res <= 0;
	4466: res <= 0;
	4467: res <= 0;
	4468: res <= 0;
	4469: res <= 0;
	4470: res <= 0;
	4471: res <= 0;
	4472: res <= 0;
	4473: res <= 0;
	4474: res <= 0;
	4475: res <= 0;
	4476: res <= 0;
	4477: res <= 0;
	4478: res <= 0;
	4479: res <= 0;
	4480: res <= 0;
	4481: res <= 0;
	4482: res <= 0;
	4483: res <= 0;
	4484: res <= 0;
	4485: res <= 0;
	4486: res <= 0;
	4487: res <= 0;
	4488: res <= 0;
	4489: res <= 0;
	4490: res <= 0;
	4491: res <= 0;
	4492: res <= 0;
	4493: res <= 0;
	4494: res <= 0;
	4495: res <= 0;
	4496: res <= 0;
	4497: res <= 0;
	4498: res <= 0;
	4499: res <= 0;
endcase
end

endmodule
