magic
tech sky130B
magscale 1 2
timestamp 1683541462
<< viali >>
rect 5825 37281 5859 37315
rect 9689 37281 9723 37315
rect 1961 37213 1995 37247
rect 6653 37213 6687 37247
rect 8493 37213 8527 37247
rect 11897 37213 11931 37247
rect 15209 37213 15243 37247
rect 18245 37213 18279 37247
rect 19625 37213 19659 37247
rect 20177 37213 20211 37247
rect 22109 37213 22143 37247
rect 25053 37213 25087 37247
rect 27169 37213 27203 37247
rect 27353 37213 27387 37247
rect 28457 37213 28491 37247
rect 32505 37213 32539 37247
rect 36921 37213 36955 37247
rect 38209 37213 38243 37247
rect 2513 37145 2547 37179
rect 5549 37145 5583 37179
rect 7021 37145 7055 37179
rect 7941 37145 7975 37179
rect 9505 37145 9539 37179
rect 12265 37145 12299 37179
rect 15761 37145 15795 37179
rect 18797 37145 18831 37179
rect 20453 37145 20487 37179
rect 22845 37145 22879 37179
rect 25881 37145 25915 37179
rect 32321 37145 32355 37179
rect 36645 37145 36679 37179
rect 37657 37145 37691 37179
rect 5181 37077 5215 37111
rect 5641 37077 5675 37111
rect 9137 37077 9171 37111
rect 9597 37077 9631 37111
rect 19533 37077 19567 37111
rect 27169 37077 27203 37111
rect 28549 37077 28583 37111
rect 6009 36873 6043 36907
rect 9597 36873 9631 36907
rect 24133 36873 24167 36907
rect 26525 36873 26559 36907
rect 4896 36805 4930 36839
rect 8484 36805 8518 36839
rect 13194 36737 13228 36771
rect 13461 36737 13495 36771
rect 14289 36737 14323 36771
rect 17049 36737 17083 36771
rect 17785 36737 17819 36771
rect 21005 36737 21039 36771
rect 22109 36737 22143 36771
rect 22376 36737 22410 36771
rect 26341 36737 26375 36771
rect 26617 36737 26651 36771
rect 27537 36737 27571 36771
rect 27804 36737 27838 36771
rect 30777 36737 30811 36771
rect 31033 36737 31067 36771
rect 32321 36737 32355 36771
rect 32577 36737 32611 36771
rect 34601 36737 34635 36771
rect 36461 36737 36495 36771
rect 37841 36737 37875 36771
rect 4629 36669 4663 36703
rect 8217 36669 8251 36703
rect 14565 36669 14599 36703
rect 18061 36669 18095 36703
rect 19993 36669 20027 36703
rect 25605 36669 25639 36703
rect 25881 36669 25915 36703
rect 34345 36669 34379 36703
rect 36645 36669 36679 36703
rect 38117 36669 38151 36703
rect 12081 36533 12115 36567
rect 16037 36533 16071 36567
rect 16957 36533 16991 36567
rect 19533 36533 19567 36567
rect 23489 36533 23523 36567
rect 26341 36533 26375 36567
rect 28917 36533 28951 36567
rect 29653 36533 29687 36567
rect 33701 36533 33735 36567
rect 35725 36533 35759 36567
rect 13461 36329 13495 36363
rect 15209 36329 15243 36363
rect 25605 36329 25639 36363
rect 27537 36329 27571 36363
rect 28273 36329 28307 36363
rect 30113 36329 30147 36363
rect 31861 36329 31895 36363
rect 33977 36329 34011 36363
rect 9229 36261 9263 36295
rect 5733 36193 5767 36227
rect 5917 36193 5951 36227
rect 9597 36193 9631 36227
rect 12909 36193 12943 36227
rect 15761 36193 15795 36227
rect 21465 36193 21499 36227
rect 26157 36193 26191 36227
rect 26433 36193 26467 36227
rect 31493 36193 31527 36227
rect 33609 36193 33643 36227
rect 34897 36193 34931 36227
rect 6469 36125 6503 36159
rect 10517 36125 10551 36159
rect 13001 36125 13035 36159
rect 15117 36125 15151 36159
rect 16129 36125 16163 36159
rect 18061 36125 18095 36159
rect 19901 36125 19935 36159
rect 20453 36125 20487 36159
rect 20729 36125 20763 36159
rect 24593 36125 24627 36159
rect 25697 36125 25731 36159
rect 28457 36125 28491 36159
rect 28733 36125 28767 36159
rect 30205 36125 30239 36159
rect 30481 36125 30515 36159
rect 31585 36125 31619 36159
rect 32965 36125 32999 36159
rect 33793 36125 33827 36159
rect 36829 36125 36863 36159
rect 5641 36057 5675 36091
rect 6736 36057 6770 36091
rect 9689 36057 9723 36091
rect 9781 36057 9815 36091
rect 10784 36057 10818 36091
rect 18337 36057 18371 36091
rect 19625 36057 19659 36091
rect 24869 36057 24903 36091
rect 32781 36057 32815 36091
rect 33149 36057 33183 36091
rect 35142 36057 35176 36091
rect 37096 36057 37130 36091
rect 5273 35989 5307 36023
rect 7849 35989 7883 36023
rect 11897 35989 11931 36023
rect 13093 35989 13127 36023
rect 17555 35989 17589 36023
rect 20453 35989 20487 36023
rect 22477 35989 22511 36023
rect 28641 35989 28675 36023
rect 29929 35989 29963 36023
rect 36277 35989 36311 36023
rect 38209 35989 38243 36023
rect 7113 35785 7147 35819
rect 7573 35785 7607 35819
rect 11713 35785 11747 35819
rect 22109 35785 22143 35819
rect 22569 35785 22603 35819
rect 32689 35785 32723 35819
rect 33425 35785 33459 35819
rect 36829 35785 36863 35819
rect 37473 35785 37507 35819
rect 7481 35649 7515 35683
rect 9873 35649 9907 35683
rect 12081 35649 12115 35683
rect 14933 35649 14967 35683
rect 17049 35649 17083 35683
rect 18245 35649 18279 35683
rect 18613 35649 18647 35683
rect 18981 35649 19015 35683
rect 19625 35649 19659 35683
rect 20545 35649 20579 35683
rect 22477 35649 22511 35683
rect 23673 35649 23707 35683
rect 23857 35649 23891 35683
rect 25421 35649 25455 35683
rect 26065 35649 26099 35683
rect 27261 35649 27295 35683
rect 28825 35649 28859 35683
rect 29092 35649 29126 35683
rect 32505 35649 32539 35683
rect 32689 35649 32723 35683
rect 33333 35649 33367 35683
rect 33517 35649 33551 35683
rect 36737 35649 36771 35683
rect 37841 35649 37875 35683
rect 7757 35581 7791 35615
rect 9965 35581 9999 35615
rect 10149 35581 10183 35615
rect 12173 35581 12207 35615
rect 12357 35581 12391 35615
rect 20821 35581 20855 35615
rect 22753 35581 22787 35615
rect 23305 35581 23339 35615
rect 24961 35581 24995 35615
rect 25513 35581 25547 35615
rect 26249 35581 26283 35615
rect 27721 35581 27755 35615
rect 37933 35581 37967 35615
rect 38025 35581 38059 35615
rect 24869 35513 24903 35547
rect 9505 35445 9539 35479
rect 14841 35445 14875 35479
rect 16957 35445 16991 35479
rect 18245 35445 18279 35479
rect 25053 35445 25087 35479
rect 30205 35445 30239 35479
rect 29101 35241 29135 35275
rect 31493 35241 31527 35275
rect 32689 35241 32723 35275
rect 11345 35173 11379 35207
rect 23489 35173 23523 35207
rect 25329 35173 25363 35207
rect 26893 35173 26927 35207
rect 5825 35105 5859 35139
rect 11805 35105 11839 35139
rect 13369 35105 13403 35139
rect 15577 35105 15611 35139
rect 17325 35105 17359 35139
rect 23397 35105 23431 35139
rect 25421 35105 25455 35139
rect 29193 35105 29227 35139
rect 36369 35105 36403 35139
rect 9137 35037 9171 35071
rect 9404 35037 9438 35071
rect 11897 35037 11931 35071
rect 13093 35037 13127 35071
rect 13277 35037 13311 35071
rect 18245 35037 18279 35071
rect 18521 35037 18555 35071
rect 19441 35037 19475 35071
rect 19717 35037 19751 35071
rect 20453 35037 20487 35071
rect 20637 35037 20671 35071
rect 22109 35037 22143 35071
rect 23857 35037 23891 35071
rect 23949 35037 23983 35071
rect 24869 35037 24903 35071
rect 24961 35037 24995 35071
rect 26617 35037 26651 35071
rect 27353 35037 27387 35071
rect 27446 35037 27480 35071
rect 28917 35037 28951 35071
rect 29009 35037 29043 35071
rect 30849 35037 30883 35071
rect 30942 35037 30976 35071
rect 31355 35037 31389 35071
rect 32965 35037 32999 35071
rect 5549 34969 5583 35003
rect 11805 34969 11839 35003
rect 12633 34969 12667 35003
rect 15853 34969 15887 35003
rect 18730 34969 18764 35003
rect 20545 34969 20579 35003
rect 21097 34969 21131 35003
rect 22385 34969 22419 35003
rect 23029 34969 23063 35003
rect 26709 34969 26743 35003
rect 26893 34969 26927 35003
rect 31125 34969 31159 35003
rect 31217 34969 31251 35003
rect 32689 34969 32723 35003
rect 36636 34969 36670 35003
rect 5181 34901 5215 34935
rect 5641 34901 5675 34935
rect 10517 34901 10551 34935
rect 18613 34901 18647 34935
rect 18889 34901 18923 34935
rect 25697 34901 25731 34935
rect 27721 34901 27755 34935
rect 32873 34901 32907 34935
rect 37749 34901 37783 34935
rect 5733 34697 5767 34731
rect 9505 34697 9539 34731
rect 9873 34697 9907 34731
rect 9965 34697 9999 34731
rect 19809 34697 19843 34731
rect 20913 34697 20947 34731
rect 25329 34697 25363 34731
rect 30113 34697 30147 34731
rect 31309 34697 31343 34731
rect 32689 34697 32723 34731
rect 37473 34697 37507 34731
rect 20315 34629 20349 34663
rect 26433 34629 26467 34663
rect 32321 34629 32355 34663
rect 32521 34629 32555 34663
rect 4353 34561 4387 34595
rect 4620 34561 4654 34595
rect 7573 34561 7607 34595
rect 7757 34561 7791 34595
rect 13369 34561 13403 34595
rect 19993 34561 20027 34595
rect 20085 34561 20119 34595
rect 20177 34561 20211 34595
rect 21097 34561 21131 34595
rect 21281 34561 21315 34595
rect 23673 34561 23707 34595
rect 24869 34561 24903 34595
rect 25145 34561 25179 34595
rect 26249 34561 26283 34595
rect 26617 34561 26651 34595
rect 27169 34561 27203 34595
rect 29469 34561 29503 34595
rect 30205 34561 30239 34595
rect 30665 34561 30699 34595
rect 30758 34561 30792 34595
rect 30941 34561 30975 34595
rect 31033 34561 31067 34595
rect 31171 34561 31205 34595
rect 33333 34561 33367 34595
rect 34253 34561 34287 34595
rect 34509 34561 34543 34595
rect 37841 34561 37875 34595
rect 7481 34493 7515 34527
rect 8217 34493 8251 34527
rect 10149 34493 10183 34527
rect 13645 34493 13679 34527
rect 15117 34493 15151 34527
rect 20453 34493 20487 34527
rect 22661 34493 22695 34527
rect 23857 34493 23891 34527
rect 24961 34493 24995 34527
rect 27629 34493 27663 34527
rect 33241 34493 33275 34527
rect 33701 34493 33735 34527
rect 37933 34493 37967 34527
rect 38025 34493 38059 34527
rect 23213 34425 23247 34459
rect 22569 34357 22603 34391
rect 22753 34357 22787 34391
rect 22845 34357 22879 34391
rect 25145 34357 25179 34391
rect 29193 34357 29227 34391
rect 32505 34357 32539 34391
rect 35633 34357 35667 34391
rect 10425 34153 10459 34187
rect 10885 34153 10919 34187
rect 20453 34153 20487 34187
rect 30389 34153 30423 34187
rect 31861 34153 31895 34187
rect 19625 34085 19659 34119
rect 28733 34085 28767 34119
rect 5549 34017 5583 34051
rect 5641 34017 5675 34051
rect 10609 34017 10643 34051
rect 21189 34017 21223 34051
rect 22109 34017 22143 34051
rect 27077 34017 27111 34051
rect 38117 34017 38151 34051
rect 7665 33949 7699 33983
rect 7849 33949 7883 33983
rect 8493 33949 8527 33983
rect 9321 33949 9355 33983
rect 9413 33949 9447 33983
rect 10701 33949 10735 33983
rect 11989 33949 12023 33983
rect 12173 33949 12207 33983
rect 15393 33949 15427 33983
rect 15577 33949 15611 33983
rect 16865 33949 16899 33983
rect 17049 33949 17083 33983
rect 17509 33949 17543 33983
rect 18429 33949 18463 33983
rect 18613 33949 18647 33983
rect 19441 33949 19475 33983
rect 19625 33949 19659 33983
rect 20269 33949 20303 33983
rect 20453 33949 20487 33983
rect 21281 33949 21315 33983
rect 22385 33949 22419 33983
rect 22477 33949 22511 33983
rect 22569 33949 22603 33983
rect 22753 33949 22787 33983
rect 23305 33949 23339 33983
rect 23581 33949 23615 33983
rect 24685 33949 24719 33983
rect 25053 33949 25087 33983
rect 25421 33949 25455 33983
rect 26157 33949 26191 33983
rect 26433 33949 26467 33983
rect 28641 33949 28675 33983
rect 28917 33949 28951 33983
rect 29745 33949 29779 33983
rect 29838 33949 29872 33983
rect 30251 33949 30285 33983
rect 31217 33949 31251 33983
rect 31365 33949 31399 33983
rect 31682 33949 31716 33983
rect 37841 33949 37875 33983
rect 5733 33881 5767 33915
rect 10425 33881 10459 33915
rect 17785 33881 17819 33915
rect 21557 33881 21591 33915
rect 21649 33881 21683 33915
rect 23213 33881 23247 33915
rect 26525 33881 26559 33915
rect 27905 33881 27939 33915
rect 30021 33881 30055 33915
rect 30113 33881 30147 33915
rect 31493 33881 31527 33915
rect 31585 33881 31619 33915
rect 6101 33813 6135 33847
rect 9137 33813 9171 33847
rect 12081 33813 12115 33847
rect 15485 33813 15519 33847
rect 17049 33813 17083 33847
rect 18521 33813 18555 33847
rect 21005 33813 21039 33847
rect 29101 33813 29135 33847
rect 13645 33609 13679 33643
rect 14749 33609 14783 33643
rect 16037 33609 16071 33643
rect 17417 33609 17451 33643
rect 20269 33609 20303 33643
rect 21373 33609 21407 33643
rect 31677 33609 31711 33643
rect 36185 33609 36219 33643
rect 7113 33541 7147 33575
rect 19165 33541 19199 33575
rect 24869 33541 24903 33575
rect 31309 33541 31343 33575
rect 33425 33541 33459 33575
rect 5917 33473 5951 33507
rect 8585 33473 8619 33507
rect 8769 33473 8803 33507
rect 9689 33473 9723 33507
rect 10149 33473 10183 33507
rect 10609 33473 10643 33507
rect 12173 33473 12207 33507
rect 12357 33473 12391 33507
rect 13277 33473 13311 33507
rect 13369 33473 13403 33507
rect 13461 33473 13495 33507
rect 14105 33473 14139 33507
rect 14565 33473 14599 33507
rect 15393 33473 15427 33507
rect 15853 33473 15887 33507
rect 18153 33473 18187 33507
rect 19349 33473 19383 33507
rect 19441 33473 19475 33507
rect 19625 33473 19659 33507
rect 19717 33473 19751 33507
rect 20177 33473 20211 33507
rect 20453 33473 20487 33507
rect 21465 33473 21499 33507
rect 22477 33473 22511 33507
rect 23121 33473 23155 33507
rect 26157 33473 26191 33507
rect 27445 33473 27479 33507
rect 28641 33473 28675 33507
rect 29837 33473 29871 33507
rect 31033 33473 31067 33507
rect 31126 33473 31160 33507
rect 31401 33473 31435 33507
rect 31539 33473 31573 33507
rect 33057 33473 33091 33507
rect 33150 33473 33184 33507
rect 33333 33473 33367 33507
rect 33563 33473 33597 33507
rect 34529 33473 34563 33507
rect 34713 33473 34747 33507
rect 34805 33473 34839 33507
rect 34897 33473 34931 33507
rect 35541 33473 35575 33507
rect 35634 33473 35668 33507
rect 35817 33473 35851 33507
rect 35909 33473 35943 33507
rect 36047 33473 36081 33507
rect 37841 33473 37875 33507
rect 6009 33405 6043 33439
rect 8217 33405 8251 33439
rect 9413 33405 9447 33439
rect 10517 33405 10551 33439
rect 14473 33405 14507 33439
rect 15669 33405 15703 33439
rect 17693 33405 17727 33439
rect 18245 33405 18279 33439
rect 22385 33405 22419 33439
rect 23213 33405 23247 33439
rect 23305 33405 23339 33439
rect 23673 33405 23707 33439
rect 25237 33405 25271 33439
rect 25605 33405 25639 33439
rect 26433 33405 26467 33439
rect 27721 33405 27755 33439
rect 29009 33405 29043 33439
rect 30297 33405 30331 33439
rect 37933 33405 37967 33439
rect 38025 33405 38059 33439
rect 12357 33337 12391 33371
rect 33701 33337 33735 33371
rect 35081 33337 35115 33371
rect 5733 33269 5767 33303
rect 7205 33269 7239 33303
rect 14197 33269 14231 33303
rect 15485 33269 15519 33303
rect 17785 33269 17819 33303
rect 20637 33269 20671 33303
rect 22109 33269 22143 33303
rect 22477 33269 22511 33303
rect 25007 33269 25041 33303
rect 25145 33269 25179 33303
rect 26249 33269 26283 33303
rect 37473 33269 37507 33303
rect 5457 33065 5491 33099
rect 7573 33065 7607 33099
rect 10793 33065 10827 33099
rect 11253 33065 11287 33099
rect 14381 33065 14415 33099
rect 15301 33065 15335 33099
rect 15669 33065 15703 33099
rect 17601 33065 17635 33099
rect 17785 33065 17819 33099
rect 18337 33065 18371 33099
rect 25237 33065 25271 33099
rect 30389 33065 30423 33099
rect 30849 33065 30883 33099
rect 32505 33065 32539 33099
rect 38209 33065 38243 33099
rect 6929 32997 6963 33031
rect 10333 32997 10367 33031
rect 12357 32997 12391 33031
rect 25421 32997 25455 33031
rect 7757 32929 7791 32963
rect 10885 32929 10919 32963
rect 14565 32929 14599 32963
rect 17417 32929 17451 32963
rect 18521 32929 18555 32963
rect 20913 32929 20947 32963
rect 23121 32929 23155 32963
rect 24777 32929 24811 32963
rect 36829 32929 36863 32963
rect 5181 32861 5215 32895
rect 5273 32861 5307 32895
rect 6837 32861 6871 32895
rect 7021 32861 7055 32895
rect 7481 32861 7515 32895
rect 8401 32861 8435 32895
rect 9873 32861 9907 32895
rect 10149 32861 10183 32895
rect 11069 32861 11103 32895
rect 12265 32861 12299 32895
rect 12449 32861 12483 32895
rect 12541 32861 12575 32895
rect 12725 32861 12759 32895
rect 13553 32861 13587 32895
rect 13737 32861 13771 32895
rect 14657 32861 14691 32895
rect 14749 32861 14783 32895
rect 15301 32861 15335 32895
rect 15393 32861 15427 32895
rect 17325 32861 17359 32895
rect 17601 32861 17635 32895
rect 18245 32861 18279 32895
rect 19625 32861 19659 32895
rect 19809 32861 19843 32895
rect 20453 32861 20487 32895
rect 20545 32861 20579 32895
rect 22937 32861 22971 32895
rect 23213 32861 23247 32895
rect 24869 32861 24903 32895
rect 25237 32861 25271 32895
rect 26249 32861 26283 32895
rect 26709 32861 26743 32895
rect 27813 32861 27847 32895
rect 28181 32861 28215 32895
rect 28733 32861 28767 32895
rect 29745 32861 29779 32895
rect 29838 32861 29872 32895
rect 30113 32861 30147 32895
rect 30251 32861 30285 32895
rect 30987 32861 31021 32895
rect 31345 32861 31379 32895
rect 31493 32861 31527 32895
rect 31953 32861 31987 32895
rect 32229 32861 32263 32895
rect 32321 32861 32355 32895
rect 35725 32861 35759 32895
rect 35863 32861 35897 32895
rect 36093 32861 36127 32895
rect 36231 32861 36265 32895
rect 37096 32861 37130 32895
rect 8217 32793 8251 32827
rect 8585 32793 8619 32827
rect 10793 32793 10827 32827
rect 20821 32793 20855 32827
rect 28917 32793 28951 32827
rect 30021 32793 30055 32827
rect 31125 32793 31159 32827
rect 31217 32793 31251 32827
rect 32137 32793 32171 32827
rect 36001 32793 36035 32827
rect 7757 32725 7791 32759
rect 9965 32725 9999 32759
rect 13737 32725 13771 32759
rect 18521 32725 18555 32759
rect 19717 32725 19751 32759
rect 20269 32725 20303 32759
rect 22753 32725 22787 32759
rect 26249 32725 26283 32759
rect 36369 32725 36403 32759
rect 12449 32521 12483 32555
rect 14749 32521 14783 32555
rect 25881 32521 25915 32555
rect 28743 32521 28777 32555
rect 30757 32521 30791 32555
rect 35449 32521 35483 32555
rect 6929 32453 6963 32487
rect 8033 32453 8067 32487
rect 10517 32453 10551 32487
rect 12265 32453 12299 32487
rect 14289 32453 14323 32487
rect 30389 32453 30423 32487
rect 35081 32453 35115 32487
rect 35173 32453 35207 32487
rect 38117 32453 38151 32487
rect 4537 32385 4571 32419
rect 4629 32385 4663 32419
rect 5273 32385 5307 32419
rect 6009 32385 6043 32419
rect 6561 32385 6595 32419
rect 6837 32385 6871 32419
rect 8769 32385 8803 32419
rect 9781 32385 9815 32419
rect 9965 32385 9999 32419
rect 10149 32385 10183 32419
rect 10333 32385 10367 32419
rect 12081 32385 12115 32419
rect 12173 32385 12207 32419
rect 14473 32385 14507 32419
rect 14565 32385 14599 32419
rect 15209 32385 15243 32419
rect 15393 32385 15427 32419
rect 16313 32385 16347 32419
rect 16865 32385 16899 32419
rect 17233 32385 17267 32419
rect 17325 32385 17359 32419
rect 20453 32385 20487 32419
rect 22201 32385 22235 32419
rect 22293 32385 22327 32419
rect 23489 32385 23523 32419
rect 23857 32385 23891 32419
rect 24409 32385 24443 32419
rect 24501 32385 24535 32419
rect 24685 32385 24719 32419
rect 25789 32385 25823 32419
rect 26249 32385 26283 32419
rect 27629 32385 27663 32419
rect 27997 32385 28031 32419
rect 28641 32385 28675 32419
rect 30113 32385 30147 32419
rect 30206 32385 30240 32419
rect 30481 32385 30515 32419
rect 30578 32385 30612 32419
rect 33037 32385 33071 32419
rect 34897 32385 34931 32419
rect 35265 32385 35299 32419
rect 37841 32385 37875 32419
rect 10057 32317 10091 32351
rect 20637 32317 20671 32351
rect 25145 32317 25179 32351
rect 32781 32317 32815 32351
rect 11897 32249 11931 32283
rect 17509 32249 17543 32283
rect 4813 32181 4847 32215
rect 5917 32181 5951 32215
rect 14289 32181 14323 32215
rect 15301 32181 15335 32215
rect 15577 32181 15611 32215
rect 16129 32181 16163 32215
rect 16957 32181 16991 32215
rect 20269 32181 20303 32215
rect 22293 32181 22327 32215
rect 23857 32181 23891 32215
rect 34161 32181 34195 32215
rect 9321 31977 9355 32011
rect 9965 31977 9999 32011
rect 10425 31977 10459 32011
rect 12173 31977 12207 32011
rect 12725 31977 12759 32011
rect 14841 31977 14875 32011
rect 15209 31977 15243 32011
rect 15853 31977 15887 32011
rect 17233 31977 17267 32011
rect 19625 31977 19659 32011
rect 23765 31977 23799 32011
rect 32781 31977 32815 32011
rect 37749 31977 37783 32011
rect 6837 31909 6871 31943
rect 6929 31909 6963 31943
rect 7205 31909 7239 31943
rect 10793 31909 10827 31943
rect 13001 31909 13035 31943
rect 13737 31909 13771 31943
rect 15669 31909 15703 31943
rect 16681 31909 16715 31943
rect 19809 31909 19843 31943
rect 22937 31909 22971 31943
rect 32321 31909 32355 31943
rect 5365 31841 5399 31875
rect 6193 31841 6227 31875
rect 14841 31841 14875 31875
rect 15945 31841 15979 31875
rect 17049 31841 17083 31875
rect 18521 31841 18555 31875
rect 19533 31841 19567 31875
rect 21557 31841 21591 31875
rect 22845 31841 22879 31875
rect 27905 31841 27939 31875
rect 28273 31841 28307 31875
rect 29837 31841 29871 31875
rect 36369 31841 36403 31875
rect 4169 31773 4203 31807
rect 4353 31773 4387 31807
rect 4813 31773 4847 31807
rect 4905 31773 4939 31807
rect 5825 31773 5859 31807
rect 6745 31773 6779 31807
rect 7021 31773 7055 31807
rect 7941 31773 7975 31807
rect 8033 31773 8067 31807
rect 8217 31773 8251 31807
rect 8309 31773 8343 31807
rect 9229 31773 9263 31807
rect 9505 31773 9539 31807
rect 9689 31773 9723 31807
rect 10425 31773 10459 31807
rect 10517 31773 10551 31807
rect 11621 31773 11655 31807
rect 11713 31773 11747 31807
rect 11897 31773 11931 31807
rect 11989 31773 12023 31807
rect 12633 31773 12667 31807
rect 12817 31773 12851 31807
rect 13461 31773 13495 31807
rect 14749 31773 14783 31807
rect 15025 31773 15059 31807
rect 16037 31773 16071 31807
rect 16865 31773 16899 31807
rect 17325 31773 17359 31807
rect 18705 31773 18739 31807
rect 19441 31773 19475 31807
rect 21189 31773 21223 31807
rect 21373 31773 21407 31807
rect 22937 31773 22971 31807
rect 23857 31773 23891 31807
rect 24593 31773 24627 31807
rect 24777 31773 24811 31807
rect 25513 31773 25547 31807
rect 25881 31773 25915 31807
rect 27169 31773 27203 31807
rect 27261 31773 27295 31807
rect 27997 31773 28031 31807
rect 28365 31773 28399 31807
rect 29745 31773 29779 31807
rect 29923 31773 29957 31807
rect 32045 31773 32079 31807
rect 32781 31773 32815 31807
rect 32965 31773 32999 31807
rect 35265 31773 35299 31807
rect 35358 31773 35392 31807
rect 35541 31773 35575 31807
rect 35633 31773 35667 31807
rect 35771 31773 35805 31807
rect 6009 31705 6043 31739
rect 13737 31705 13771 31739
rect 18889 31705 18923 31739
rect 22661 31705 22695 31739
rect 24041 31705 24075 31739
rect 26985 31705 27019 31739
rect 29009 31705 29043 31739
rect 32321 31705 32355 31739
rect 36636 31705 36670 31739
rect 4077 31637 4111 31671
rect 7757 31637 7791 31671
rect 9597 31637 9631 31671
rect 13553 31637 13587 31671
rect 21189 31637 21223 31671
rect 24685 31637 24719 31671
rect 32137 31637 32171 31671
rect 35909 31637 35943 31671
rect 10241 31433 10275 31467
rect 12265 31433 12299 31467
rect 18889 31433 18923 31467
rect 22109 31433 22143 31467
rect 25053 31433 25087 31467
rect 28457 31433 28491 31467
rect 31309 31433 31343 31467
rect 32505 31433 32539 31467
rect 32689 31433 32723 31467
rect 34897 31433 34931 31467
rect 36553 31433 36587 31467
rect 36921 31433 36955 31467
rect 7389 31365 7423 31399
rect 8217 31365 8251 31399
rect 11897 31365 11931 31399
rect 12081 31365 12115 31399
rect 13461 31365 13495 31399
rect 15393 31365 15427 31399
rect 15761 31365 15795 31399
rect 30941 31365 30975 31399
rect 31033 31365 31067 31399
rect 32321 31365 32355 31399
rect 38117 31365 38151 31399
rect 4813 31297 4847 31331
rect 4997 31297 5031 31331
rect 5825 31297 5859 31331
rect 6009 31297 6043 31331
rect 6561 31297 6595 31331
rect 6745 31297 6779 31331
rect 8861 31297 8895 31331
rect 9965 31297 9999 31331
rect 10149 31297 10183 31331
rect 12725 31297 12759 31331
rect 12909 31297 12943 31331
rect 14289 31297 14323 31331
rect 16957 31297 16991 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 18705 31297 18739 31331
rect 19625 31297 19659 31331
rect 19809 31297 19843 31331
rect 21281 31297 21315 31331
rect 21465 31297 21499 31331
rect 22109 31297 22143 31331
rect 22477 31297 22511 31331
rect 23397 31297 23431 31331
rect 23673 31297 23707 31331
rect 24593 31297 24627 31331
rect 24869 31297 24903 31331
rect 26065 31297 26099 31331
rect 26157 31297 26191 31331
rect 26249 31297 26283 31331
rect 26433 31297 26467 31331
rect 27261 31297 27295 31331
rect 27813 31297 27847 31331
rect 28365 31297 28399 31331
rect 28641 31297 28675 31331
rect 29193 31297 29227 31331
rect 29377 31297 29411 31331
rect 30665 31297 30699 31331
rect 30758 31297 30792 31331
rect 31130 31297 31164 31331
rect 34345 31297 34379 31331
rect 34529 31297 34563 31331
rect 34621 31297 34655 31331
rect 34713 31297 34747 31331
rect 36461 31297 36495 31331
rect 37841 31297 37875 31331
rect 6653 31229 6687 31263
rect 9045 31229 9079 31263
rect 9137 31229 9171 31263
rect 17325 31229 17359 31263
rect 17417 31229 17451 31263
rect 19441 31229 19475 31263
rect 19717 31229 19751 31263
rect 19901 31229 19935 31263
rect 23489 31229 23523 31263
rect 23857 31229 23891 31263
rect 36369 31229 36403 31263
rect 24685 31161 24719 31195
rect 5181 31093 5215 31127
rect 5733 31093 5767 31127
rect 8677 31093 8711 31127
rect 12725 31093 12759 31127
rect 18337 31093 18371 31127
rect 21465 31093 21499 31127
rect 25789 31093 25823 31127
rect 29193 31093 29227 31127
rect 32505 31093 32539 31127
rect 6745 30889 6779 30923
rect 7021 30889 7055 30923
rect 8217 30889 8251 30923
rect 12449 30889 12483 30923
rect 14565 30889 14599 30923
rect 14749 30889 14783 30923
rect 18061 30889 18095 30923
rect 19901 30889 19935 30923
rect 20453 30889 20487 30923
rect 21097 30889 21131 30923
rect 24041 30889 24075 30923
rect 25145 30889 25179 30923
rect 25973 30889 26007 30923
rect 26341 30889 26375 30923
rect 28457 30889 28491 30923
rect 4905 30821 4939 30855
rect 6101 30821 6135 30855
rect 7849 30821 7883 30855
rect 7941 30821 7975 30855
rect 9413 30821 9447 30855
rect 19441 30821 19475 30855
rect 26801 30821 26835 30855
rect 30021 30821 30055 30855
rect 31401 30821 31435 30855
rect 6653 30753 6687 30787
rect 11713 30753 11747 30787
rect 13553 30753 13587 30787
rect 13737 30753 13771 30787
rect 14473 30753 14507 30787
rect 15669 30753 15703 30787
rect 19717 30753 19751 30787
rect 20637 30753 20671 30787
rect 25053 30753 25087 30787
rect 32229 30753 32263 30787
rect 32689 30753 32723 30787
rect 5733 30685 5767 30719
rect 6837 30685 6871 30719
rect 7757 30685 7791 30719
rect 8033 30685 8067 30719
rect 9413 30685 9447 30719
rect 10425 30685 10459 30719
rect 11805 30685 11839 30719
rect 11989 30685 12023 30719
rect 12173 30685 12207 30719
rect 13461 30685 13495 30719
rect 14289 30685 14323 30719
rect 14565 30685 14599 30719
rect 15393 30685 15427 30719
rect 15577 30685 15611 30719
rect 15761 30685 15795 30719
rect 15945 30685 15979 30719
rect 16497 30685 16531 30719
rect 16681 30685 16715 30719
rect 16865 30685 16899 30719
rect 17785 30685 17819 30719
rect 17877 30685 17911 30719
rect 19625 30685 19659 30719
rect 20361 30685 20395 30719
rect 21097 30685 21131 30719
rect 22477 30685 22511 30719
rect 22661 30685 22695 30719
rect 23857 30685 23891 30719
rect 24041 30685 24075 30719
rect 25329 30685 25363 30719
rect 25973 30685 26007 30719
rect 26065 30685 26099 30719
rect 27169 30685 27203 30719
rect 27629 30685 27663 30719
rect 27813 30685 27847 30719
rect 28273 30685 28307 30719
rect 28457 30685 28491 30719
rect 29837 30685 29871 30719
rect 29929 30685 29963 30719
rect 30757 30685 30791 30719
rect 30850 30685 30884 30719
rect 31033 30685 31067 30719
rect 31222 30685 31256 30719
rect 32321 30685 32355 30719
rect 37841 30685 37875 30719
rect 5089 30617 5123 30651
rect 5273 30617 5307 30651
rect 5917 30617 5951 30651
rect 6561 30617 6595 30651
rect 18061 30617 18095 30651
rect 19901 30617 19935 30651
rect 26985 30617 27019 30651
rect 31125 30617 31159 30651
rect 38117 30617 38151 30651
rect 12081 30549 12115 30583
rect 13737 30549 13771 30583
rect 15209 30549 15243 30583
rect 17601 30549 17635 30583
rect 20637 30549 20671 30583
rect 22845 30549 22879 30583
rect 25513 30549 25547 30583
rect 27721 30549 27755 30583
rect 28641 30549 28675 30583
rect 13185 30345 13219 30379
rect 16129 30345 16163 30379
rect 30389 30345 30423 30379
rect 34989 30345 35023 30379
rect 9873 30277 9907 30311
rect 10333 30277 10367 30311
rect 15117 30277 15151 30311
rect 24593 30277 24627 30311
rect 24777 30277 24811 30311
rect 30021 30277 30055 30311
rect 33876 30277 33910 30311
rect 37841 30277 37875 30311
rect 2789 30209 2823 30243
rect 3056 30209 3090 30243
rect 4813 30209 4847 30243
rect 4997 30209 5031 30243
rect 5549 30209 5583 30243
rect 5825 30209 5859 30243
rect 7205 30209 7239 30243
rect 7757 30209 7791 30243
rect 8585 30209 8619 30243
rect 8769 30209 8803 30243
rect 9689 30209 9723 30243
rect 10517 30209 10551 30243
rect 10609 30209 10643 30243
rect 11713 30209 11747 30243
rect 11805 30209 11839 30243
rect 13093 30209 13127 30243
rect 13277 30209 13311 30243
rect 14565 30209 14599 30243
rect 15393 30209 15427 30243
rect 16221 30209 16255 30243
rect 17785 30209 17819 30243
rect 17877 30209 17911 30243
rect 18337 30209 18371 30243
rect 18521 30209 18555 30243
rect 20177 30209 20211 30243
rect 20361 30209 20395 30243
rect 22661 30209 22695 30243
rect 23397 30209 23431 30243
rect 23857 30209 23891 30243
rect 24041 30209 24075 30243
rect 24961 30209 24995 30243
rect 25421 30209 25455 30243
rect 25605 30209 25639 30243
rect 25973 30209 26007 30243
rect 27629 30209 27663 30243
rect 29009 30209 29043 30243
rect 29193 30209 29227 30243
rect 29745 30209 29779 30243
rect 29838 30209 29872 30243
rect 30113 30209 30147 30243
rect 30251 30209 30285 30243
rect 32505 30209 32539 30243
rect 32689 30209 32723 30243
rect 35633 30209 35667 30243
rect 35726 30209 35760 30243
rect 35909 30209 35943 30243
rect 36001 30209 36035 30243
rect 36139 30209 36173 30243
rect 5641 30141 5675 30175
rect 5733 30141 5767 30175
rect 8401 30141 8435 30175
rect 9413 30141 9447 30175
rect 15209 30141 15243 30175
rect 23029 30141 23063 30175
rect 26065 30141 26099 30175
rect 27905 30141 27939 30175
rect 33609 30141 33643 30175
rect 37933 30141 37967 30175
rect 38025 30141 38059 30175
rect 10793 30073 10827 30107
rect 12081 30073 12115 30107
rect 15577 30073 15611 30107
rect 17509 30073 17543 30107
rect 22826 30073 22860 30107
rect 22937 30073 22971 30107
rect 24041 30073 24075 30107
rect 36277 30073 36311 30107
rect 4169 30005 4203 30039
rect 4813 30005 4847 30039
rect 6009 30005 6043 30039
rect 9505 30005 9539 30039
rect 10333 30005 10367 30039
rect 11713 30005 11747 30039
rect 14473 30005 14507 30039
rect 15117 30005 15151 30039
rect 17693 30005 17727 30039
rect 18521 30005 18555 30039
rect 19993 30005 20027 30039
rect 26525 30005 26559 30039
rect 29009 30005 29043 30039
rect 32505 30005 32539 30039
rect 37473 30005 37507 30039
rect 3985 29801 4019 29835
rect 11897 29801 11931 29835
rect 12081 29801 12115 29835
rect 17233 29801 17267 29835
rect 17417 29801 17451 29835
rect 20729 29801 20763 29835
rect 22293 29801 22327 29835
rect 23397 29801 23431 29835
rect 26065 29801 26099 29835
rect 28622 29801 28656 29835
rect 30389 29801 30423 29835
rect 32137 29801 32171 29835
rect 34253 29801 34287 29835
rect 35449 29801 35483 29835
rect 36277 29801 36311 29835
rect 38209 29801 38243 29835
rect 11529 29733 11563 29767
rect 21557 29733 21591 29767
rect 22845 29733 22879 29767
rect 26249 29733 26283 29767
rect 28733 29733 28767 29767
rect 3433 29665 3467 29699
rect 4629 29665 4663 29699
rect 17509 29665 17543 29699
rect 21465 29665 21499 29699
rect 21649 29665 21683 29699
rect 28825 29665 28859 29699
rect 36829 29665 36863 29699
rect 3157 29597 3191 29631
rect 3341 29597 3375 29631
rect 6009 29597 6043 29631
rect 7205 29597 7239 29631
rect 7297 29597 7331 29631
rect 7573 29597 7607 29631
rect 7757 29597 7791 29631
rect 9321 29597 9355 29631
rect 15025 29597 15059 29631
rect 16497 29597 16531 29631
rect 16681 29597 16715 29631
rect 17417 29597 17451 29631
rect 20361 29597 20395 29631
rect 20453 29597 20487 29631
rect 20821 29597 20855 29631
rect 21741 29597 21775 29631
rect 22477 29597 22511 29631
rect 22661 29597 22695 29631
rect 23305 29597 23339 29631
rect 23489 29597 23523 29631
rect 26985 29597 27019 29631
rect 27445 29597 27479 29631
rect 28457 29597 28491 29631
rect 29745 29597 29779 29631
rect 29893 29597 29927 29631
rect 30021 29597 30055 29631
rect 30251 29597 30285 29631
rect 31033 29597 31067 29631
rect 31126 29597 31160 29631
rect 31498 29597 31532 29631
rect 32413 29597 32447 29631
rect 32873 29597 32907 29631
rect 34897 29597 34931 29631
rect 35265 29597 35299 29631
rect 36093 29597 36127 29631
rect 37096 29597 37130 29631
rect 26111 29563 26145 29597
rect 2973 29529 3007 29563
rect 4445 29529 4479 29563
rect 5733 29529 5767 29563
rect 10885 29529 10919 29563
rect 11897 29529 11931 29563
rect 12633 29529 12667 29563
rect 13461 29529 13495 29563
rect 14289 29529 14323 29563
rect 17693 29529 17727 29563
rect 22201 29529 22235 29563
rect 25881 29529 25915 29563
rect 29193 29529 29227 29563
rect 30113 29529 30147 29563
rect 31309 29529 31343 29563
rect 31401 29529 31435 29563
rect 32137 29529 32171 29563
rect 33140 29529 33174 29563
rect 35081 29529 35115 29563
rect 35173 29529 35207 29563
rect 4353 29461 4387 29495
rect 7573 29461 7607 29495
rect 16589 29461 16623 29495
rect 21005 29461 21039 29495
rect 27077 29461 27111 29495
rect 31677 29461 31711 29495
rect 32321 29461 32355 29495
rect 9413 29257 9447 29291
rect 11161 29257 11195 29291
rect 14657 29257 14691 29291
rect 16313 29257 16347 29291
rect 19257 29257 19291 29291
rect 23397 29257 23431 29291
rect 24961 29257 24995 29291
rect 32505 29257 32539 29291
rect 32689 29257 32723 29291
rect 4353 29189 4387 29223
rect 4445 29189 4479 29223
rect 6745 29189 6779 29223
rect 6929 29189 6963 29223
rect 8953 29189 8987 29223
rect 11713 29189 11747 29223
rect 11897 29189 11931 29223
rect 14289 29189 14323 29223
rect 14381 29189 14415 29223
rect 17417 29189 17451 29223
rect 28457 29189 28491 29223
rect 28549 29189 28583 29223
rect 31677 29189 31711 29223
rect 32321 29189 32355 29223
rect 35081 29189 35115 29223
rect 37933 29189 37967 29223
rect 4261 29121 4295 29155
rect 4629 29121 4663 29155
rect 5273 29121 5307 29155
rect 5549 29121 5583 29155
rect 8125 29121 8159 29155
rect 8401 29121 8435 29155
rect 9229 29121 9263 29155
rect 9965 29121 9999 29155
rect 10057 29121 10091 29155
rect 10977 29121 11011 29155
rect 11161 29121 11195 29155
rect 12173 29121 12207 29155
rect 12633 29121 12667 29155
rect 12817 29121 12851 29155
rect 13277 29121 13311 29155
rect 13461 29121 13495 29155
rect 14105 29121 14139 29155
rect 14473 29121 14507 29155
rect 16129 29121 16163 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17877 29121 17911 29155
rect 18797 29121 18831 29155
rect 19533 29121 19567 29155
rect 19625 29121 19659 29155
rect 19717 29121 19751 29155
rect 19901 29121 19935 29155
rect 20361 29121 20395 29155
rect 22569 29121 22603 29155
rect 22753 29121 22787 29155
rect 23581 29121 23615 29155
rect 23673 29121 23707 29155
rect 23765 29121 23799 29155
rect 23857 29121 23891 29155
rect 25973 29121 26007 29155
rect 27169 29121 27203 29155
rect 27537 29121 27571 29155
rect 28365 29121 28399 29155
rect 28733 29121 28767 29155
rect 29193 29121 29227 29155
rect 30389 29121 30423 29155
rect 30757 29121 30791 29155
rect 31309 29121 31343 29155
rect 31493 29121 31527 29155
rect 34897 29121 34931 29155
rect 35173 29121 35207 29155
rect 35265 29121 35299 29155
rect 36461 29121 36495 29155
rect 37565 29121 37599 29155
rect 5457 29053 5491 29087
rect 9045 29053 9079 29087
rect 15853 29053 15887 29087
rect 15945 29053 15979 29087
rect 18245 29053 18279 29087
rect 20637 29053 20671 29087
rect 20821 29053 20855 29087
rect 25145 29053 25179 29087
rect 25237 29053 25271 29087
rect 25329 29053 25363 29087
rect 25421 29053 25455 29087
rect 26065 29053 26099 29087
rect 27353 29053 27387 29087
rect 29377 29053 29411 29087
rect 36737 29053 36771 29087
rect 4077 28985 4111 29019
rect 5089 28985 5123 29019
rect 8125 28985 8159 29019
rect 13645 28985 13679 29019
rect 18337 28985 18371 29019
rect 20453 28985 20487 29019
rect 22937 28985 22971 29019
rect 26341 28985 26375 29019
rect 28181 28985 28215 29019
rect 5365 28917 5399 28951
rect 6653 28917 6687 28951
rect 8953 28917 8987 28951
rect 9965 28917 9999 28951
rect 11897 28917 11931 28951
rect 12633 28917 12667 28951
rect 13461 28917 13495 28951
rect 18429 28917 18463 28951
rect 25973 28917 26007 28951
rect 27261 28917 27295 28951
rect 32505 28917 32539 28951
rect 35449 28917 35483 28951
rect 4629 28713 4663 28747
rect 10333 28713 10367 28747
rect 11897 28713 11931 28747
rect 12541 28713 12575 28747
rect 15117 28713 15151 28747
rect 17693 28713 17727 28747
rect 19809 28713 19843 28747
rect 27077 28713 27111 28747
rect 31125 28713 31159 28747
rect 32321 28713 32355 28747
rect 7481 28645 7515 28679
rect 16405 28645 16439 28679
rect 24961 28645 24995 28679
rect 25053 28645 25087 28679
rect 10425 28577 10459 28611
rect 15025 28577 15059 28611
rect 16129 28577 16163 28611
rect 16497 28577 16531 28611
rect 21465 28577 21499 28611
rect 25145 28577 25179 28611
rect 32965 28577 32999 28611
rect 33425 28577 33459 28611
rect 36645 28577 36679 28611
rect 4721 28509 4755 28543
rect 5457 28509 5491 28543
rect 6653 28509 6687 28543
rect 6929 28509 6963 28543
rect 7389 28509 7423 28543
rect 7573 28509 7607 28543
rect 9137 28509 9171 28543
rect 9597 28509 9631 28543
rect 10609 28509 10643 28543
rect 12541 28509 12575 28543
rect 12725 28509 12759 28543
rect 14749 28509 14783 28543
rect 14887 28509 14921 28543
rect 15209 28509 15243 28543
rect 16313 28509 16347 28543
rect 16589 28509 16623 28543
rect 16773 28509 16807 28543
rect 17601 28509 17635 28543
rect 17785 28509 17819 28543
rect 19441 28509 19475 28543
rect 21189 28509 21223 28543
rect 23121 28509 23155 28543
rect 23213 28509 23247 28543
rect 23489 28509 23523 28543
rect 23765 28509 23799 28543
rect 24041 28509 24075 28543
rect 24593 28509 24627 28543
rect 27353 28509 27387 28543
rect 28273 28509 28307 28543
rect 28641 28509 28675 28543
rect 30665 28509 30699 28543
rect 31217 28509 31251 28543
rect 31677 28509 31711 28543
rect 31770 28509 31804 28543
rect 31953 28509 31987 28543
rect 32142 28509 32176 28543
rect 33057 28509 33091 28543
rect 35541 28509 35575 28543
rect 35634 28509 35668 28543
rect 35817 28509 35851 28543
rect 35909 28509 35943 28543
rect 36047 28509 36081 28543
rect 5641 28441 5675 28475
rect 6561 28441 6595 28475
rect 10333 28441 10367 28475
rect 12081 28441 12115 28475
rect 19625 28441 19659 28475
rect 21557 28441 21591 28475
rect 21674 28441 21708 28475
rect 22569 28441 22603 28475
rect 27169 28441 27203 28475
rect 28365 28441 28399 28475
rect 28457 28441 28491 28475
rect 32045 28441 32079 28475
rect 36912 28441 36946 28475
rect 5273 28373 5307 28407
rect 9229 28373 9263 28407
rect 10793 28373 10827 28407
rect 11713 28373 11747 28407
rect 11897 28373 11931 28407
rect 21833 28373 21867 28407
rect 25421 28373 25455 28407
rect 28089 28373 28123 28407
rect 36185 28373 36219 28407
rect 38025 28373 38059 28407
rect 14657 28169 14691 28203
rect 16957 28169 16991 28203
rect 25973 28169 26007 28203
rect 28549 28169 28583 28203
rect 30389 28169 30423 28203
rect 37473 28169 37507 28203
rect 37841 28169 37875 28203
rect 6837 28101 6871 28135
rect 25145 28101 25179 28135
rect 27813 28101 27847 28135
rect 30021 28101 30055 28135
rect 31033 28101 31067 28135
rect 34406 28101 34440 28135
rect 37933 28101 37967 28135
rect 4997 28033 5031 28067
rect 5089 28033 5123 28067
rect 5181 28033 5215 28067
rect 5365 28033 5399 28067
rect 9321 28033 9355 28067
rect 9505 28033 9539 28067
rect 10241 28033 10275 28067
rect 10517 28033 10551 28067
rect 12633 28033 12667 28067
rect 13461 28033 13495 28067
rect 14105 28033 14139 28067
rect 14473 28033 14507 28067
rect 16865 28033 16899 28067
rect 17049 28033 17083 28067
rect 20177 28033 20211 28067
rect 22385 28033 22419 28067
rect 22661 28033 22695 28067
rect 23213 28033 23247 28067
rect 24041 28033 24075 28067
rect 25421 28033 25455 28067
rect 25973 28033 26007 28067
rect 26249 28033 26283 28067
rect 27353 28033 27387 28067
rect 28365 28033 28399 28067
rect 29745 28033 29779 28067
rect 29838 28033 29872 28067
rect 30113 28033 30147 28067
rect 30251 28033 30285 28067
rect 31769 28033 31803 28067
rect 32321 28033 32355 28067
rect 32413 28033 32447 28067
rect 32597 28033 32631 28067
rect 32689 28033 32723 28067
rect 32873 28033 32907 28067
rect 7205 27965 7239 27999
rect 10425 27965 10459 27999
rect 13369 27965 13403 27999
rect 20269 27965 20303 27999
rect 27445 27965 27479 27999
rect 34161 27965 34195 27999
rect 38025 27965 38059 27999
rect 10701 27897 10735 27931
rect 22385 27897 22419 27931
rect 24501 27897 24535 27931
rect 4813 27829 4847 27863
rect 6653 27829 6687 27863
rect 6837 27829 6871 27863
rect 9413 27829 9447 27863
rect 10241 27829 10275 27863
rect 14197 27829 14231 27863
rect 20177 27829 20211 27863
rect 20545 27829 20579 27863
rect 23397 27829 23431 27863
rect 27169 27829 27203 27863
rect 27537 27829 27571 27863
rect 35541 27829 35575 27863
rect 18705 27625 18739 27659
rect 31125 27625 31159 27659
rect 31493 27625 31527 27659
rect 4261 27557 4295 27591
rect 10701 27557 10735 27591
rect 16957 27557 16991 27591
rect 18521 27557 18555 27591
rect 23581 27557 23615 27591
rect 23765 27557 23799 27591
rect 30481 27557 30515 27591
rect 33517 27557 33551 27591
rect 4353 27489 4387 27523
rect 5365 27489 5399 27523
rect 7297 27489 7331 27523
rect 7933 27489 7967 27523
rect 16865 27489 16899 27523
rect 18705 27489 18739 27523
rect 18797 27489 18831 27523
rect 19441 27489 19475 27523
rect 26985 27489 27019 27523
rect 31125 27489 31159 27523
rect 32689 27489 32723 27523
rect 37197 27489 37231 27523
rect 4169 27421 4203 27455
rect 4445 27421 4479 27455
rect 4629 27421 4663 27455
rect 5089 27421 5123 27455
rect 5273 27421 5307 27455
rect 5457 27421 5491 27455
rect 5641 27421 5675 27455
rect 7113 27421 7147 27455
rect 8022 27421 8056 27455
rect 8125 27421 8159 27455
rect 8217 27421 8251 27455
rect 9137 27421 9171 27455
rect 9321 27421 9355 27455
rect 10517 27421 10551 27455
rect 12357 27421 12391 27455
rect 16773 27421 16807 27455
rect 17049 27421 17083 27455
rect 18889 27421 18923 27455
rect 20177 27421 20211 27455
rect 21557 27421 21591 27455
rect 22201 27421 22235 27455
rect 22661 27421 22695 27455
rect 26341 27421 26375 27455
rect 26525 27421 26559 27455
rect 26617 27421 26651 27455
rect 26709 27421 26743 27455
rect 27445 27421 27479 27455
rect 27629 27421 27663 27455
rect 27721 27421 27755 27455
rect 27813 27421 27847 27455
rect 29837 27421 29871 27455
rect 29930 27421 29964 27455
rect 30113 27421 30147 27455
rect 30343 27421 30377 27455
rect 31033 27421 31067 27455
rect 31309 27421 31343 27455
rect 32965 27421 32999 27455
rect 33701 27421 33735 27455
rect 34069 27421 34103 27455
rect 34897 27421 34931 27455
rect 34989 27421 35023 27455
rect 35173 27421 35207 27455
rect 36921 27421 36955 27455
rect 37841 27421 37875 27455
rect 10333 27353 10367 27387
rect 12624 27353 12658 27387
rect 19993 27353 20027 27387
rect 21097 27353 21131 27387
rect 24041 27353 24075 27387
rect 25237 27353 25271 27387
rect 25421 27353 25455 27387
rect 30205 27353 30239 27387
rect 33793 27353 33827 27387
rect 33885 27353 33919 27387
rect 35357 27353 35391 27387
rect 38117 27353 38151 27387
rect 3985 27285 4019 27319
rect 5825 27285 5859 27319
rect 6929 27285 6963 27319
rect 7757 27285 7791 27319
rect 9229 27285 9263 27319
rect 13737 27285 13771 27319
rect 16589 27285 16623 27319
rect 19625 27285 19659 27319
rect 20085 27285 20119 27319
rect 22385 27285 22419 27319
rect 25053 27285 25087 27319
rect 28089 27285 28123 27319
rect 4169 27081 4203 27115
rect 6745 27081 6779 27115
rect 7297 27081 7331 27115
rect 12817 27081 12851 27115
rect 15945 27081 15979 27115
rect 20177 27081 20211 27115
rect 22477 27081 22511 27115
rect 24593 27081 24627 27115
rect 26341 27081 26375 27115
rect 37933 27081 37967 27115
rect 3056 27013 3090 27047
rect 5549 27013 5583 27047
rect 13185 27013 13219 27047
rect 22017 27013 22051 27047
rect 24041 27013 24075 27047
rect 26157 27013 26191 27047
rect 30389 27013 30423 27047
rect 31401 27013 31435 27047
rect 34805 27013 34839 27047
rect 35633 27013 35667 27047
rect 2789 26945 2823 26979
rect 5089 26945 5123 26979
rect 5273 26945 5307 26979
rect 6561 26945 6595 26979
rect 6837 26945 6871 26979
rect 7297 26945 7331 26979
rect 7481 26945 7515 26979
rect 8033 26945 8067 26979
rect 8309 26945 8343 26979
rect 8907 26945 8941 26979
rect 9045 26945 9079 26979
rect 9137 26945 9171 26979
rect 9229 26945 9263 26979
rect 10241 26945 10275 26979
rect 10425 26945 10459 26979
rect 13001 26945 13035 26979
rect 13093 26945 13127 26979
rect 13369 26945 13403 26979
rect 14832 26945 14866 26979
rect 17417 26945 17451 26979
rect 18061 26945 18095 26979
rect 18981 26945 19015 26979
rect 19257 26945 19291 26979
rect 20085 26945 20119 26979
rect 20269 26945 20303 26979
rect 20821 26945 20855 26979
rect 22293 26945 22327 26979
rect 22937 26945 22971 26979
rect 23213 26945 23247 26979
rect 23949 26945 23983 26979
rect 24133 26945 24167 26979
rect 24777 26945 24811 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 25237 26945 25271 26979
rect 27629 26945 27663 26979
rect 28089 26945 28123 26979
rect 29101 26945 29135 26979
rect 29745 26945 29779 26979
rect 30849 26945 30883 26979
rect 31217 26945 31251 26979
rect 32597 26945 32631 26979
rect 34161 26945 34195 26979
rect 34345 26945 34379 26979
rect 37841 26945 37875 26979
rect 8769 26877 8803 26911
rect 14565 26877 14599 26911
rect 17141 26877 17175 26911
rect 18153 26877 18187 26911
rect 20913 26877 20947 26911
rect 22109 26877 22143 26911
rect 23029 26877 23063 26911
rect 28365 26877 28399 26911
rect 33333 26877 33367 26911
rect 38025 26877 38059 26911
rect 8033 26809 8067 26843
rect 9413 26809 9447 26843
rect 17049 26809 17083 26843
rect 18981 26809 19015 26843
rect 21189 26809 21223 26843
rect 23397 26809 23431 26843
rect 24961 26809 24995 26843
rect 26525 26809 26559 26843
rect 4905 26741 4939 26775
rect 5457 26741 5491 26775
rect 6561 26741 6595 26775
rect 10241 26741 10275 26775
rect 21005 26741 21039 26775
rect 22293 26741 22327 26775
rect 23029 26741 23063 26775
rect 26341 26741 26375 26775
rect 34345 26741 34379 26775
rect 37473 26741 37507 26775
rect 9321 26537 9355 26571
rect 14749 26537 14783 26571
rect 22845 26537 22879 26571
rect 23489 26537 23523 26571
rect 35541 26537 35575 26571
rect 37933 26537 37967 26571
rect 21557 26469 21591 26503
rect 28273 26469 28307 26503
rect 30941 26469 30975 26503
rect 34069 26469 34103 26503
rect 5089 26401 5123 26435
rect 6009 26401 6043 26435
rect 11069 26401 11103 26435
rect 15209 26401 15243 26435
rect 15301 26401 15335 26435
rect 16037 26401 16071 26435
rect 20637 26401 20671 26435
rect 22661 26401 22695 26435
rect 30297 26401 30331 26435
rect 32321 26401 32355 26435
rect 33241 26401 33275 26435
rect 33425 26401 33459 26435
rect 36553 26401 36587 26435
rect 5181 26333 5215 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 5917 26333 5951 26367
rect 6101 26333 6135 26367
rect 8309 26333 8343 26367
rect 8585 26333 8619 26367
rect 10609 26333 10643 26367
rect 15117 26333 15151 26367
rect 16221 26333 16255 26367
rect 17049 26333 17083 26367
rect 17601 26333 17635 26367
rect 17693 26333 17727 26367
rect 18245 26333 18279 26367
rect 19625 26333 19659 26367
rect 19717 26333 19751 26367
rect 20913 26333 20947 26367
rect 21097 26333 21131 26367
rect 21760 26333 21794 26367
rect 22017 26333 22051 26367
rect 22845 26333 22879 26367
rect 23489 26333 23523 26367
rect 23673 26333 23707 26367
rect 24777 26333 24811 26367
rect 24961 26333 24995 26367
rect 25053 26333 25087 26367
rect 25145 26333 25179 26367
rect 25329 26333 25363 26367
rect 27721 26333 27755 26367
rect 27905 26333 27939 26367
rect 27997 26333 28031 26367
rect 28089 26333 28123 26367
rect 29745 26333 29779 26367
rect 29929 26333 29963 26367
rect 33149 26333 33183 26367
rect 34069 26333 34103 26367
rect 34253 26333 34287 26367
rect 34989 26333 35023 26367
rect 35081 26333 35115 26367
rect 35265 26333 35299 26367
rect 35357 26333 35391 26367
rect 36820 26333 36854 26367
rect 8217 26265 8251 26299
rect 9505 26265 9539 26299
rect 11314 26265 11348 26299
rect 16405 26265 16439 26299
rect 19441 26265 19475 26299
rect 22569 26265 22603 26299
rect 24593 26265 24627 26299
rect 32076 26265 32110 26299
rect 4905 26197 4939 26231
rect 9137 26197 9171 26231
rect 9305 26197 9339 26231
rect 10425 26197 10459 26231
rect 12449 26197 12483 26231
rect 18061 26197 18095 26231
rect 21925 26197 21959 26231
rect 23029 26197 23063 26231
rect 30205 26197 30239 26231
rect 32781 26197 32815 26231
rect 5641 25993 5675 26027
rect 11161 25993 11195 26027
rect 12817 25993 12851 26027
rect 17325 25993 17359 26027
rect 20453 25993 20487 26027
rect 31217 25993 31251 26027
rect 34529 25993 34563 26027
rect 6745 25925 6779 25959
rect 9689 25925 9723 25959
rect 17049 25925 17083 25959
rect 17417 25925 17451 25959
rect 27905 25925 27939 25959
rect 29009 25925 29043 25959
rect 34253 25925 34287 25959
rect 36378 25925 36412 25959
rect 5457 25857 5491 25891
rect 5733 25857 5767 25891
rect 6653 25857 6687 25891
rect 6837 25857 6871 25891
rect 8125 25857 8159 25891
rect 8585 25857 8619 25891
rect 9965 25857 9999 25891
rect 10609 25857 10643 25891
rect 10793 25857 10827 25891
rect 10885 25857 10919 25891
rect 10977 25857 11011 25891
rect 12725 25857 12759 25891
rect 13001 25857 13035 25891
rect 14105 25857 14139 25891
rect 14381 25857 14415 25891
rect 17233 25857 17267 25891
rect 18153 25857 18187 25891
rect 18613 25857 18647 25891
rect 20637 25857 20671 25891
rect 22017 25857 22051 25891
rect 22201 25857 22235 25891
rect 23305 25857 23339 25891
rect 23581 25857 23615 25891
rect 27721 25857 27755 25891
rect 27813 25857 27847 25891
rect 28089 25857 28123 25891
rect 30205 25857 30239 25891
rect 30665 25857 30699 25891
rect 30757 25857 30791 25891
rect 30941 25857 30975 25891
rect 31033 25857 31067 25891
rect 33977 25857 34011 25891
rect 34161 25857 34195 25891
rect 34345 25857 34379 25891
rect 37841 25857 37875 25891
rect 5273 25789 5307 25823
rect 5365 25789 5399 25823
rect 8217 25789 8251 25823
rect 9781 25789 9815 25823
rect 18521 25789 18555 25823
rect 20085 25789 20119 25823
rect 20177 25789 20211 25823
rect 22569 25789 22603 25823
rect 36645 25789 36679 25823
rect 38117 25789 38151 25823
rect 23305 25721 23339 25755
rect 4997 25653 5031 25687
rect 9965 25653 9999 25687
rect 10149 25653 10183 25687
rect 13185 25653 13219 25687
rect 17601 25653 17635 25687
rect 27537 25653 27571 25687
rect 35265 25653 35299 25687
rect 6561 25449 6595 25483
rect 9505 25449 9539 25483
rect 14289 25449 14323 25483
rect 25237 25449 25271 25483
rect 4353 25381 4387 25415
rect 18613 25381 18647 25415
rect 28733 25381 28767 25415
rect 32597 25381 32631 25415
rect 4905 25313 4939 25347
rect 5273 25313 5307 25347
rect 5365 25313 5399 25347
rect 6837 25313 6871 25347
rect 7573 25313 7607 25347
rect 16681 25313 16715 25347
rect 19441 25313 19475 25347
rect 27445 25313 27479 25347
rect 28641 25313 28675 25347
rect 29929 25313 29963 25347
rect 30389 25313 30423 25347
rect 33057 25313 33091 25347
rect 4169 25245 4203 25279
rect 4445 25245 4479 25279
rect 6745 25245 6779 25279
rect 6929 25245 6963 25279
rect 7021 25245 7055 25279
rect 9781 25245 9815 25279
rect 12357 25245 12391 25279
rect 12624 25245 12658 25279
rect 14473 25245 14507 25279
rect 14749 25245 14783 25279
rect 16129 25245 16163 25279
rect 16221 25245 16255 25279
rect 16589 25245 16623 25279
rect 18245 25245 18279 25279
rect 18429 25245 18463 25279
rect 18521 25245 18555 25279
rect 18705 25245 18739 25279
rect 19625 25245 19659 25279
rect 19993 25245 20027 25279
rect 20545 25245 20579 25279
rect 21005 25245 21039 25279
rect 23121 25245 23155 25279
rect 23581 25245 23615 25279
rect 25145 25245 25179 25279
rect 26157 25245 26191 25279
rect 26249 25245 26283 25279
rect 26525 25245 26559 25279
rect 27077 25245 27111 25279
rect 27261 25245 27295 25279
rect 28549 25245 28583 25279
rect 28825 25245 28859 25279
rect 30021 25245 30055 25279
rect 31953 25245 31987 25279
rect 32046 25245 32080 25279
rect 32418 25245 32452 25279
rect 33425 25245 33459 25279
rect 33609 25245 33643 25279
rect 34989 25245 35023 25279
rect 35817 25245 35851 25279
rect 36645 25245 36679 25279
rect 7757 25177 7791 25211
rect 7941 25177 7975 25211
rect 9321 25177 9355 25211
rect 14657 25177 14691 25211
rect 17233 25177 17267 25211
rect 19901 25177 19935 25211
rect 24961 25177 24995 25211
rect 26341 25177 26375 25211
rect 30297 25177 30331 25211
rect 32229 25177 32263 25211
rect 32321 25177 32355 25211
rect 36912 25177 36946 25211
rect 3985 25109 4019 25143
rect 5549 25109 5583 25143
rect 9505 25109 9539 25143
rect 13737 25109 13771 25143
rect 18889 25109 18923 25143
rect 20729 25109 20763 25143
rect 22661 25109 22695 25143
rect 25973 25109 26007 25143
rect 29009 25109 29043 25143
rect 29745 25109 29779 25143
rect 33425 25109 33459 25143
rect 38025 25109 38059 25143
rect 19257 24905 19291 24939
rect 24317 24905 24351 24939
rect 37473 24905 37507 24939
rect 3056 24837 3090 24871
rect 7021 24837 7055 24871
rect 8401 24837 8435 24871
rect 8601 24837 8635 24871
rect 10425 24837 10459 24871
rect 13461 24837 13495 24871
rect 21281 24837 21315 24871
rect 25053 24837 25087 24871
rect 37841 24837 37875 24871
rect 2789 24769 2823 24803
rect 5089 24769 5123 24803
rect 6837 24769 6871 24803
rect 7113 24769 7147 24803
rect 9413 24769 9447 24803
rect 10241 24769 10275 24803
rect 10517 24769 10551 24803
rect 10609 24769 10643 24803
rect 13277 24769 13311 24803
rect 13553 24769 13587 24803
rect 13645 24769 13679 24803
rect 14565 24769 14599 24803
rect 16865 24769 16899 24803
rect 17693 24769 17727 24803
rect 18061 24769 18095 24803
rect 18521 24769 18555 24803
rect 19073 24769 19107 24803
rect 19257 24769 19291 24803
rect 20269 24769 20303 24803
rect 23121 24769 23155 24803
rect 23305 24769 23339 24803
rect 23489 24769 23523 24803
rect 23765 24769 23799 24803
rect 24317 24769 24351 24803
rect 24593 24769 24627 24803
rect 25237 24769 25271 24803
rect 25789 24769 25823 24803
rect 27629 24769 27663 24803
rect 27905 24769 27939 24803
rect 29009 24769 29043 24803
rect 29469 24769 29503 24803
rect 29561 24769 29595 24803
rect 30113 24769 30147 24803
rect 30389 24769 30423 24803
rect 33793 24769 33827 24803
rect 34969 24769 35003 24803
rect 5181 24701 5215 24735
rect 5273 24701 5307 24735
rect 5365 24701 5399 24735
rect 5549 24701 5583 24735
rect 9229 24701 9263 24735
rect 14289 24701 14323 24735
rect 22937 24701 22971 24735
rect 28089 24701 28123 24735
rect 28825 24701 28859 24735
rect 30849 24701 30883 24735
rect 33885 24701 33919 24735
rect 34161 24701 34195 24735
rect 34713 24701 34747 24735
rect 37933 24701 37967 24735
rect 38117 24701 38151 24735
rect 6837 24633 6871 24667
rect 13829 24633 13863 24667
rect 15853 24633 15887 24667
rect 30205 24633 30239 24667
rect 4169 24565 4203 24599
rect 8585 24565 8619 24599
rect 8769 24565 8803 24599
rect 9597 24565 9631 24599
rect 10793 24565 10827 24599
rect 18429 24565 18463 24599
rect 27721 24565 27755 24599
rect 36093 24565 36127 24599
rect 11989 24361 12023 24395
rect 23213 24361 23247 24395
rect 34161 24361 34195 24395
rect 34897 24361 34931 24395
rect 27077 24293 27111 24327
rect 9321 24225 9355 24259
rect 9413 24225 9447 24259
rect 9597 24225 9631 24259
rect 20821 24225 20855 24259
rect 23305 24225 23339 24259
rect 24593 24225 24627 24259
rect 26341 24225 26375 24259
rect 30573 24225 30607 24259
rect 32413 24225 32447 24259
rect 35265 24225 35299 24259
rect 5733 24157 5767 24191
rect 5825 24157 5859 24191
rect 6009 24157 6043 24191
rect 6837 24157 6871 24191
rect 7113 24157 7147 24191
rect 7665 24157 7699 24191
rect 9505 24157 9539 24191
rect 10609 24157 10643 24191
rect 17233 24157 17267 24191
rect 17417 24157 17451 24191
rect 17785 24157 17819 24191
rect 17969 24157 18003 24191
rect 18245 24157 18279 24191
rect 19625 24157 19659 24191
rect 21465 24157 21499 24191
rect 21833 24157 21867 24191
rect 22017 24157 22051 24191
rect 23029 24157 23063 24191
rect 23857 24157 23891 24191
rect 24041 24157 24075 24191
rect 24869 24157 24903 24191
rect 26801 24157 26835 24191
rect 27261 24157 27295 24191
rect 28043 24157 28077 24191
rect 28456 24157 28490 24191
rect 28549 24157 28583 24191
rect 29837 24157 29871 24191
rect 29929 24157 29963 24191
rect 30113 24157 30147 24191
rect 31217 24157 31251 24191
rect 31365 24157 31399 24191
rect 31585 24157 31619 24191
rect 31682 24157 31716 24191
rect 32321 24157 32355 24191
rect 32597 24157 32631 24191
rect 32689 24157 32723 24191
rect 33793 24157 33827 24191
rect 33977 24157 34011 24191
rect 35081 24157 35115 24191
rect 37841 24157 37875 24191
rect 10876 24089 10910 24123
rect 18705 24089 18739 24123
rect 19717 24089 19751 24123
rect 20729 24089 20763 24123
rect 24961 24089 24995 24123
rect 25329 24089 25363 24123
rect 28181 24089 28215 24123
rect 28273 24089 28307 24123
rect 31493 24089 31527 24123
rect 38117 24089 38151 24123
rect 6193 24021 6227 24055
rect 6653 24021 6687 24055
rect 7021 24021 7055 24055
rect 7757 24021 7791 24055
rect 9137 24021 9171 24055
rect 20269 24021 20303 24055
rect 20637 24021 20671 24055
rect 22845 24021 22879 24055
rect 23949 24021 23983 24055
rect 24777 24021 24811 24055
rect 27905 24021 27939 24055
rect 31861 24021 31895 24055
rect 32873 24021 32907 24055
rect 4169 23817 4203 23851
rect 33333 23817 33367 23851
rect 33891 23817 33925 23851
rect 35541 23817 35575 23851
rect 8668 23749 8702 23783
rect 27813 23749 27847 23783
rect 27997 23749 28031 23783
rect 30205 23749 30239 23783
rect 32965 23749 32999 23783
rect 33793 23749 33827 23783
rect 33977 23749 34011 23783
rect 35173 23749 35207 23783
rect 36553 23749 36587 23783
rect 37933 23749 37967 23783
rect 2789 23681 2823 23715
rect 3056 23681 3090 23715
rect 4813 23681 4847 23715
rect 4905 23681 4939 23715
rect 5089 23681 5123 23715
rect 5181 23681 5215 23715
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 6745 23681 6779 23715
rect 8401 23681 8435 23715
rect 12725 23681 12759 23715
rect 12981 23681 13015 23715
rect 16865 23681 16899 23715
rect 17049 23681 17083 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 20545 23681 20579 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 24225 23681 24259 23715
rect 24777 23681 24811 23715
rect 25605 23681 25639 23715
rect 27721 23681 27755 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 28825 23681 28859 23715
rect 29009 23681 29043 23715
rect 29469 23681 29503 23715
rect 29745 23681 29779 23715
rect 31033 23681 31067 23715
rect 31585 23681 31619 23715
rect 32689 23681 32723 23715
rect 32837 23681 32871 23715
rect 33057 23681 33091 23715
rect 33195 23681 33229 23715
rect 34069 23681 34103 23715
rect 34897 23681 34931 23715
rect 34990 23681 35024 23715
rect 35265 23681 35299 23715
rect 35362 23681 35396 23715
rect 36001 23681 36035 23715
rect 36277 23681 36311 23715
rect 36369 23681 36403 23715
rect 37841 23681 37875 23715
rect 5733 23613 5767 23647
rect 17417 23613 17451 23647
rect 25789 23613 25823 23647
rect 26065 23613 26099 23647
rect 26157 23613 26191 23647
rect 29561 23613 29595 23647
rect 30849 23613 30883 23647
rect 38117 23613 38151 23647
rect 20361 23545 20395 23579
rect 23489 23545 23523 23579
rect 27997 23545 28031 23579
rect 31585 23545 31619 23579
rect 36093 23545 36127 23579
rect 4629 23477 4663 23511
rect 6837 23477 6871 23511
rect 9781 23477 9815 23511
rect 14105 23477 14139 23511
rect 20729 23477 20763 23511
rect 25053 23477 25087 23511
rect 28457 23477 28491 23511
rect 37473 23477 37507 23511
rect 3985 23273 4019 23307
rect 5181 23273 5215 23307
rect 5549 23273 5583 23307
rect 22753 23273 22787 23307
rect 22937 23273 22971 23307
rect 26249 23273 26283 23307
rect 35909 23273 35943 23307
rect 38209 23273 38243 23307
rect 6469 23205 6503 23239
rect 10701 23205 10735 23239
rect 12541 23205 12575 23239
rect 14933 23205 14967 23239
rect 27353 23205 27387 23239
rect 4537 23137 4571 23171
rect 5641 23137 5675 23171
rect 16589 23137 16623 23171
rect 20361 23137 20395 23171
rect 20453 23137 20487 23171
rect 23029 23137 23063 23171
rect 25513 23137 25547 23171
rect 35725 23137 35759 23171
rect 4445 23069 4479 23103
rect 5365 23069 5399 23103
rect 6377 23069 6411 23103
rect 6561 23069 6595 23103
rect 6653 23069 6687 23103
rect 10149 23069 10183 23103
rect 10517 23069 10551 23103
rect 11161 23069 11195 23103
rect 14289 23069 14323 23103
rect 15209 23069 15243 23103
rect 15853 23069 15887 23103
rect 22937 23069 22971 23103
rect 25329 23069 25363 23103
rect 26709 23069 26743 23103
rect 27537 23069 27571 23103
rect 29745 23069 29779 23103
rect 30205 23069 30239 23103
rect 30573 23069 30607 23103
rect 35357 23069 35391 23103
rect 35633 23069 35667 23103
rect 36829 23069 36863 23103
rect 37096 23069 37130 23103
rect 4353 23001 4387 23035
rect 10333 23001 10367 23035
rect 10425 23001 10459 23035
rect 11406 23001 11440 23035
rect 14933 23001 14967 23035
rect 16834 23001 16868 23035
rect 20269 23001 20303 23035
rect 21097 23001 21131 23035
rect 21281 23001 21315 23035
rect 23397 23001 23431 23035
rect 25145 23001 25179 23035
rect 35265 23001 35299 23035
rect 6837 22933 6871 22967
rect 14381 22933 14415 22967
rect 15117 22933 15151 22967
rect 15761 22933 15795 22967
rect 17969 22933 18003 22967
rect 19901 22933 19935 22967
rect 21465 22933 21499 22967
rect 30849 22933 30883 22967
rect 5825 22729 5859 22763
rect 8585 22729 8619 22763
rect 8861 22729 8895 22763
rect 20085 22729 20119 22763
rect 20545 22729 20579 22763
rect 24593 22729 24627 22763
rect 7757 22661 7791 22695
rect 8493 22661 8527 22695
rect 11980 22661 12014 22695
rect 27997 22661 28031 22695
rect 33241 22661 33275 22695
rect 5917 22593 5951 22627
rect 7481 22593 7515 22627
rect 7573 22593 7607 22627
rect 8677 22593 8711 22627
rect 11713 22593 11747 22627
rect 14473 22593 14507 22627
rect 14657 22593 14691 22627
rect 15209 22593 15243 22627
rect 15393 22593 15427 22627
rect 15485 22593 15519 22627
rect 15577 22593 15611 22627
rect 15715 22593 15749 22627
rect 18521 22593 18555 22627
rect 18889 22593 18923 22627
rect 20177 22593 20211 22627
rect 22241 22593 22275 22627
rect 22385 22593 22419 22627
rect 22477 22593 22511 22627
rect 22661 22593 22695 22627
rect 24501 22593 24535 22627
rect 24685 22593 24719 22627
rect 25697 22593 25731 22627
rect 25789 22593 25823 22627
rect 26157 22593 26191 22627
rect 27859 22593 27893 22627
rect 28089 22593 28123 22627
rect 28272 22593 28306 22627
rect 28365 22593 28399 22627
rect 30573 22593 30607 22627
rect 30941 22593 30975 22627
rect 31033 22593 31067 22627
rect 31585 22593 31619 22627
rect 33425 22593 33459 22627
rect 37841 22593 37875 22627
rect 14289 22525 14323 22559
rect 15853 22525 15887 22559
rect 19349 22525 19383 22559
rect 19993 22525 20027 22559
rect 31125 22525 31159 22559
rect 33609 22525 33643 22559
rect 38117 22525 38151 22559
rect 8309 22457 8343 22491
rect 26341 22457 26375 22491
rect 7297 22389 7331 22423
rect 7481 22389 7515 22423
rect 13093 22389 13127 22423
rect 22109 22389 22143 22423
rect 27721 22389 27755 22423
rect 7205 22185 7239 22219
rect 27997 22185 28031 22219
rect 31677 22185 31711 22219
rect 15945 22117 15979 22151
rect 23489 22117 23523 22151
rect 29193 22117 29227 22151
rect 4629 22049 4663 22083
rect 14749 22049 14783 22083
rect 23029 22049 23063 22083
rect 25053 22049 25087 22083
rect 33609 22049 33643 22083
rect 34069 22049 34103 22083
rect 35633 22049 35667 22083
rect 4445 21981 4479 22015
rect 6285 21981 6319 22015
rect 6561 21981 6595 22015
rect 7481 21981 7515 22015
rect 7573 21981 7607 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 9597 21981 9631 22015
rect 14907 21981 14941 22015
rect 15025 21981 15059 22015
rect 15209 21981 15243 22015
rect 16037 21981 16071 22015
rect 20729 21981 20763 22015
rect 20996 21981 21030 22015
rect 23121 21981 23155 22015
rect 25237 21981 25271 22015
rect 25881 21981 25915 22015
rect 26985 21981 27019 22015
rect 27077 21981 27111 22015
rect 27353 21981 27387 22015
rect 27813 21981 27847 22015
rect 27997 21981 28031 22015
rect 28549 21981 28583 22015
rect 28642 21981 28676 22015
rect 28825 21981 28859 22015
rect 28914 21981 28948 22015
rect 29055 21981 29089 22015
rect 29929 21981 29963 22015
rect 30021 21981 30055 22015
rect 30297 21981 30331 22015
rect 31125 21981 31159 22015
rect 31401 21981 31435 22015
rect 31493 21981 31527 22015
rect 32551 21981 32585 22015
rect 32781 21981 32815 22015
rect 32964 21981 32998 22015
rect 33057 21981 33091 22015
rect 33701 21981 33735 22015
rect 35541 21981 35575 22015
rect 35817 21981 35851 22015
rect 35909 21981 35943 22015
rect 36829 21981 36863 22015
rect 6377 21913 6411 21947
rect 9864 21913 9898 21947
rect 15117 21913 15151 21947
rect 27169 21913 27203 21947
rect 30113 21913 30147 21947
rect 31033 21913 31067 21947
rect 32689 21913 32723 21947
rect 37096 21913 37130 21947
rect 3985 21845 4019 21879
rect 4353 21845 4387 21879
rect 6745 21845 6779 21879
rect 10977 21845 11011 21879
rect 15393 21845 15427 21879
rect 22109 21845 22143 21879
rect 25789 21845 25823 21879
rect 26801 21845 26835 21879
rect 29745 21845 29779 21879
rect 32413 21845 32447 21879
rect 36093 21845 36127 21879
rect 38209 21845 38243 21879
rect 4445 21641 4479 21675
rect 9965 21641 9999 21675
rect 14473 21641 14507 21675
rect 18889 21641 18923 21675
rect 32781 21641 32815 21675
rect 35081 21641 35115 21675
rect 36277 21641 36311 21675
rect 37473 21641 37507 21675
rect 37933 21641 37967 21675
rect 3332 21573 3366 21607
rect 10333 21573 10367 21607
rect 17601 21573 17635 21607
rect 17969 21573 18003 21607
rect 18705 21573 18739 21607
rect 23152 21573 23186 21607
rect 32597 21573 32631 21607
rect 33968 21573 34002 21607
rect 35909 21573 35943 21607
rect 36001 21573 36035 21607
rect 37841 21573 37875 21607
rect 5641 21505 5675 21539
rect 6561 21505 6595 21539
rect 6745 21505 6779 21539
rect 6837 21505 6871 21539
rect 6929 21505 6963 21539
rect 7941 21505 7975 21539
rect 8033 21505 8067 21539
rect 8217 21505 8251 21539
rect 8953 21505 8987 21539
rect 9045 21505 9079 21539
rect 10149 21505 10183 21539
rect 10425 21505 10459 21539
rect 11161 21505 11195 21539
rect 14473 21505 14507 21539
rect 14657 21505 14691 21539
rect 15853 21505 15887 21539
rect 15945 21505 15979 21539
rect 17877 21505 17911 21539
rect 18337 21505 18371 21539
rect 23397 21505 23431 21539
rect 24317 21505 24351 21539
rect 27169 21505 27203 21539
rect 27353 21505 27387 21539
rect 28733 21505 28767 21539
rect 28825 21505 28859 21539
rect 29009 21505 29043 21539
rect 29101 21505 29135 21539
rect 29745 21505 29779 21539
rect 29837 21505 29871 21539
rect 32873 21505 32907 21539
rect 35633 21505 35667 21539
rect 35726 21505 35760 21539
rect 36098 21505 36132 21539
rect 3065 21437 3099 21471
rect 5457 21437 5491 21471
rect 5825 21437 5859 21471
rect 8125 21437 8159 21471
rect 10885 21437 10919 21471
rect 16221 21437 16255 21471
rect 16313 21437 16347 21471
rect 24501 21437 24535 21471
rect 24593 21437 24627 21471
rect 24685 21437 24719 21471
rect 24777 21437 24811 21471
rect 30113 21437 30147 21471
rect 30205 21437 30239 21471
rect 33701 21437 33735 21471
rect 38025 21437 38059 21471
rect 11069 21369 11103 21403
rect 29561 21369 29595 21403
rect 32597 21369 32631 21403
rect 7113 21301 7147 21335
rect 8401 21301 8435 21335
rect 8953 21301 8987 21335
rect 10977 21301 11011 21335
rect 15669 21301 15703 21335
rect 22017 21301 22051 21335
rect 24961 21301 24995 21335
rect 27353 21301 27387 21335
rect 28549 21301 28583 21335
rect 6009 21097 6043 21131
rect 9689 21097 9723 21131
rect 15945 21097 15979 21131
rect 16681 21097 16715 21131
rect 28273 21097 28307 21131
rect 31290 21097 31324 21131
rect 31769 21097 31803 21131
rect 36093 21097 36127 21131
rect 12725 21029 12759 21063
rect 20913 21029 20947 21063
rect 31401 21029 31435 21063
rect 14933 20961 14967 20995
rect 15485 20961 15519 20995
rect 26157 20961 26191 20995
rect 31493 20961 31527 20995
rect 35449 20961 35483 20995
rect 35541 20961 35575 20995
rect 4629 20893 4663 20927
rect 10333 20893 10367 20927
rect 10517 20893 10551 20927
rect 10609 20893 10643 20927
rect 10701 20893 10735 20927
rect 11345 20893 11379 20927
rect 15669 20893 15703 20927
rect 15761 20893 15795 20927
rect 16037 20893 16071 20927
rect 16773 20893 16807 20927
rect 16865 20893 16899 20927
rect 22385 20893 22419 20927
rect 23069 20893 23103 20927
rect 23213 20893 23247 20927
rect 23305 20893 23339 20927
rect 23489 20893 23523 20927
rect 24593 20893 24627 20927
rect 24777 20893 24811 20927
rect 25053 20893 25087 20927
rect 26433 20893 26467 20927
rect 27169 20893 27203 20927
rect 27629 20893 27663 20927
rect 27722 20893 27756 20927
rect 27905 20893 27939 20927
rect 27997 20893 28031 20927
rect 28094 20893 28128 20927
rect 35817 20893 35851 20927
rect 35909 20893 35943 20927
rect 37841 20893 37875 20927
rect 4896 20825 4930 20859
rect 9505 20825 9539 20859
rect 9721 20825 9755 20859
rect 11590 20825 11624 20859
rect 14657 20825 14691 20859
rect 22920 20825 22954 20859
rect 31125 20825 31159 20859
rect 38117 20825 38151 20859
rect 9873 20757 9907 20791
rect 10885 20757 10919 20791
rect 14289 20757 14323 20791
rect 14749 20757 14783 20791
rect 16497 20757 16531 20791
rect 24961 20757 24995 20791
rect 27077 20757 27111 20791
rect 7941 20553 7975 20587
rect 14381 20553 14415 20587
rect 14933 20553 14967 20587
rect 20821 20553 20855 20587
rect 33517 20553 33551 20587
rect 13268 20485 13302 20519
rect 27445 20485 27479 20519
rect 35817 20485 35851 20519
rect 37933 20485 37967 20519
rect 6561 20417 6595 20451
rect 6828 20417 6862 20451
rect 15301 20417 15335 20451
rect 17417 20417 17451 20451
rect 18521 20417 18555 20451
rect 19441 20417 19475 20451
rect 19697 20417 19731 20451
rect 22385 20417 22419 20451
rect 24593 20417 24627 20451
rect 25513 20417 25547 20451
rect 25605 20417 25639 20451
rect 25697 20417 25731 20451
rect 27169 20417 27203 20451
rect 27353 20417 27387 20451
rect 27537 20417 27571 20451
rect 29561 20417 29595 20451
rect 30665 20417 30699 20451
rect 30757 20417 30791 20451
rect 31067 20417 31101 20451
rect 33149 20417 33183 20451
rect 33333 20417 33367 20451
rect 35265 20417 35299 20451
rect 35541 20417 35575 20451
rect 35633 20417 35667 20451
rect 37841 20417 37875 20451
rect 13001 20349 13035 20383
rect 15393 20349 15427 20383
rect 15577 20349 15611 20383
rect 17141 20349 17175 20383
rect 18337 20349 18371 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 24777 20349 24811 20383
rect 29285 20349 29319 20383
rect 38025 20349 38059 20383
rect 22017 20281 22051 20315
rect 29377 20281 29411 20315
rect 31309 20281 31343 20315
rect 17233 20213 17267 20247
rect 17601 20213 17635 20247
rect 27721 20213 27755 20247
rect 29745 20213 29779 20247
rect 35357 20213 35391 20247
rect 37473 20213 37507 20247
rect 7113 20009 7147 20043
rect 15301 20009 15335 20043
rect 17141 20009 17175 20043
rect 17601 20009 17635 20043
rect 19441 20009 19475 20043
rect 25053 20009 25087 20043
rect 26525 20009 26559 20043
rect 29837 20009 29871 20043
rect 35541 20009 35575 20043
rect 18521 19941 18555 19975
rect 21465 19941 21499 19975
rect 26636 19941 26670 19975
rect 31493 19941 31527 19975
rect 4629 19873 4663 19907
rect 9137 19873 9171 19907
rect 15945 19873 15979 19907
rect 17233 19873 17267 19907
rect 19993 19873 20027 19907
rect 23213 19873 23247 19907
rect 24685 19873 24719 19907
rect 26433 19873 26467 19907
rect 30941 19873 30975 19907
rect 33517 19873 33551 19907
rect 33977 19873 34011 19907
rect 4537 19805 4571 19839
rect 6561 19805 6595 19839
rect 6837 19805 6871 19839
rect 6929 19805 6963 19839
rect 8125 19805 8159 19839
rect 8309 19805 8343 19839
rect 11713 19805 11747 19839
rect 14749 19805 14783 19839
rect 15761 19805 15795 19839
rect 17417 19805 17451 19839
rect 18245 19805 18279 19839
rect 18337 19805 18371 19839
rect 18613 19805 18647 19839
rect 19901 19805 19935 19839
rect 21644 19805 21678 19839
rect 21741 19805 21775 19839
rect 22017 19805 22051 19839
rect 22477 19805 22511 19839
rect 22845 19805 22879 19839
rect 23397 19805 23431 19839
rect 24777 19805 24811 19839
rect 26801 19805 26835 19839
rect 27261 19805 27295 19839
rect 27445 19805 27479 19839
rect 28549 19805 28583 19839
rect 28642 19805 28676 19839
rect 28917 19805 28951 19839
rect 29014 19805 29048 19839
rect 29745 19805 29779 19839
rect 29837 19805 29871 19839
rect 32321 19805 32355 19839
rect 32414 19805 32448 19839
rect 32686 19805 32720 19839
rect 32827 19805 32861 19839
rect 33609 19805 33643 19839
rect 34897 19805 34931 19839
rect 34990 19805 35024 19839
rect 35265 19805 35299 19839
rect 35362 19805 35396 19839
rect 36737 19805 36771 19839
rect 37004 19805 37038 19839
rect 6745 19737 6779 19771
rect 9382 19737 9416 19771
rect 11437 19737 11471 19771
rect 17141 19737 17175 19771
rect 19809 19737 19843 19771
rect 21833 19737 21867 19771
rect 27813 19737 27847 19771
rect 28825 19737 28859 19771
rect 31033 19737 31067 19771
rect 31217 19737 31251 19771
rect 32597 19737 32631 19771
rect 35173 19737 35207 19771
rect 4077 19669 4111 19703
rect 4445 19669 4479 19703
rect 8217 19669 8251 19703
rect 10517 19669 10551 19703
rect 14657 19669 14691 19703
rect 15669 19669 15703 19703
rect 18061 19669 18095 19703
rect 26157 19669 26191 19703
rect 29193 19669 29227 19703
rect 30113 19669 30147 19703
rect 32965 19669 32999 19703
rect 38117 19669 38151 19703
rect 5641 19465 5675 19499
rect 5733 19465 5767 19499
rect 9137 19465 9171 19499
rect 13093 19465 13127 19499
rect 15117 19465 15151 19499
rect 15577 19465 15611 19499
rect 25145 19465 25179 19499
rect 32682 19465 32716 19499
rect 35725 19465 35759 19499
rect 3700 19397 3734 19431
rect 9413 19397 9447 19431
rect 10793 19397 10827 19431
rect 10885 19397 10919 19431
rect 11958 19397 11992 19431
rect 14657 19397 14691 19431
rect 21281 19397 21315 19431
rect 29561 19397 29595 19431
rect 32597 19397 32631 19431
rect 32781 19397 32815 19431
rect 3433 19329 3467 19363
rect 6837 19329 6871 19363
rect 7021 19329 7055 19363
rect 9321 19329 9355 19363
rect 9505 19329 9539 19363
rect 9689 19329 9723 19363
rect 10609 19329 10643 19363
rect 10977 19329 11011 19363
rect 11713 19329 11747 19363
rect 14841 19329 14875 19363
rect 14933 19329 14967 19363
rect 15945 19329 15979 19363
rect 17325 19329 17359 19363
rect 17417 19329 17451 19363
rect 17601 19329 17635 19363
rect 17693 19329 17727 19363
rect 19441 19329 19475 19363
rect 20170 19329 20204 19363
rect 20453 19329 20487 19363
rect 20637 19329 20671 19363
rect 21465 19329 21499 19363
rect 22293 19329 22327 19363
rect 22753 19329 22787 19363
rect 23029 19329 23063 19363
rect 23121 19329 23155 19363
rect 23397 19329 23431 19363
rect 23581 19329 23615 19363
rect 24593 19329 24627 19363
rect 27169 19329 27203 19363
rect 27629 19329 27663 19363
rect 28641 19329 28675 19363
rect 28825 19329 28859 19363
rect 29285 19329 29319 19363
rect 29433 19329 29467 19363
rect 29653 19329 29687 19363
rect 29750 19329 29784 19363
rect 32505 19329 32539 19363
rect 33241 19329 33275 19363
rect 33333 19329 33367 19363
rect 33517 19329 33551 19363
rect 34345 19329 34379 19363
rect 34601 19329 34635 19363
rect 37841 19329 37875 19363
rect 38117 19329 38151 19363
rect 5917 19261 5951 19295
rect 16037 19261 16071 19295
rect 16221 19261 16255 19295
rect 19073 19261 19107 19295
rect 21097 19261 21131 19295
rect 24869 19261 24903 19295
rect 27905 19261 27939 19295
rect 4813 19193 4847 19227
rect 11161 19193 11195 19227
rect 28825 19193 28859 19227
rect 5273 19125 5307 19159
rect 6929 19125 6963 19159
rect 14933 19125 14967 19159
rect 17141 19125 17175 19159
rect 19993 19125 20027 19159
rect 24777 19125 24811 19159
rect 29929 19125 29963 19159
rect 33517 19125 33551 19159
rect 5825 18921 5859 18955
rect 15577 18921 15611 18955
rect 17785 18921 17819 18955
rect 19993 18921 20027 18955
rect 24593 18921 24627 18955
rect 24777 18921 24811 18955
rect 33425 18921 33459 18955
rect 18153 18853 18187 18887
rect 6745 18785 6779 18819
rect 7113 18785 7147 18819
rect 7205 18785 7239 18819
rect 13645 18785 13679 18819
rect 14841 18785 14875 18819
rect 19441 18785 19475 18819
rect 37749 18785 37783 18819
rect 4445 18717 4479 18751
rect 6837 18717 6871 18751
rect 9321 18717 9355 18751
rect 9689 18717 9723 18751
rect 12357 18717 12391 18751
rect 15485 18717 15519 18751
rect 17969 18717 18003 18751
rect 18245 18717 18279 18751
rect 19809 18717 19843 18751
rect 21281 18717 21315 18751
rect 21465 18717 21499 18751
rect 24777 18717 24811 18751
rect 24961 18717 24995 18751
rect 26157 18717 26191 18751
rect 26433 18717 26467 18751
rect 26525 18717 26559 18751
rect 28181 18717 28215 18751
rect 28549 18717 28583 18751
rect 30849 18717 30883 18751
rect 31309 18717 31343 18751
rect 31861 18717 31895 18751
rect 32045 18717 32079 18751
rect 32781 18717 32815 18751
rect 32929 18717 32963 18751
rect 33057 18717 33091 18751
rect 33246 18717 33280 18751
rect 4712 18649 4746 18683
rect 9413 18649 9447 18683
rect 9505 18649 9539 18683
rect 12449 18649 12483 18683
rect 14657 18649 14691 18683
rect 21373 18649 21407 18683
rect 26341 18649 26375 18683
rect 28273 18649 28307 18683
rect 28365 18649 28399 18683
rect 32321 18649 32355 18683
rect 33149 18649 33183 18683
rect 37473 18649 37507 18683
rect 6561 18581 6595 18615
rect 9137 18581 9171 18615
rect 13001 18581 13035 18615
rect 13369 18581 13403 18615
rect 13461 18581 13495 18615
rect 14289 18581 14323 18615
rect 14749 18581 14783 18615
rect 19625 18581 19659 18615
rect 26709 18581 26743 18615
rect 27997 18581 28031 18615
rect 37105 18581 37139 18615
rect 37565 18581 37599 18615
rect 18981 18377 19015 18411
rect 19073 18377 19107 18411
rect 19809 18377 19843 18411
rect 21465 18377 21499 18411
rect 22017 18377 22051 18411
rect 24869 18377 24903 18411
rect 29653 18377 29687 18411
rect 33241 18377 33275 18411
rect 36645 18377 36679 18411
rect 12081 18309 12115 18343
rect 16865 18309 16899 18343
rect 20269 18309 20303 18343
rect 21005 18309 21039 18343
rect 33609 18309 33643 18343
rect 35265 18309 35299 18343
rect 35357 18309 35391 18343
rect 8309 18241 8343 18275
rect 8576 18241 8610 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 10425 18241 10459 18275
rect 10517 18241 10551 18275
rect 12357 18241 12391 18275
rect 13185 18241 13219 18275
rect 14749 18241 14783 18275
rect 14933 18241 14967 18275
rect 20177 18241 20211 18275
rect 21281 18241 21315 18275
rect 22201 18241 22235 18275
rect 22293 18241 22327 18275
rect 22477 18241 22511 18275
rect 23305 18241 23339 18275
rect 23397 18241 23431 18275
rect 23581 18241 23615 18275
rect 23765 18241 23799 18275
rect 24593 18241 24627 18275
rect 25329 18241 25363 18275
rect 25513 18241 25547 18275
rect 25605 18241 25639 18275
rect 28181 18241 28215 18275
rect 29193 18241 29227 18275
rect 29655 18241 29689 18275
rect 33425 18241 33459 18275
rect 34989 18241 35023 18275
rect 35082 18241 35116 18275
rect 35454 18241 35488 18275
rect 36093 18241 36127 18275
rect 36369 18241 36403 18275
rect 36461 18241 36495 18275
rect 37841 18241 37875 18275
rect 12173 18173 12207 18207
rect 13461 18173 13495 18207
rect 17601 18173 17635 18207
rect 19257 18173 19291 18207
rect 20361 18173 20395 18207
rect 21097 18173 21131 18207
rect 24225 18173 24259 18207
rect 24685 18173 24719 18207
rect 28089 18173 28123 18207
rect 38117 18173 38151 18207
rect 9689 18105 9723 18139
rect 12541 18105 12575 18139
rect 13369 18105 13403 18139
rect 29285 18105 29319 18139
rect 35633 18105 35667 18139
rect 10701 18037 10735 18071
rect 12357 18037 12391 18071
rect 13001 18037 13035 18071
rect 14749 18037 14783 18071
rect 18613 18037 18647 18071
rect 21005 18037 21039 18071
rect 22385 18037 22419 18071
rect 25329 18037 25363 18071
rect 27813 18037 27847 18071
rect 29837 18037 29871 18071
rect 36185 18037 36219 18071
rect 7389 17833 7423 17867
rect 10149 17833 10183 17867
rect 17141 17833 17175 17867
rect 23121 17833 23155 17867
rect 29101 17833 29135 17867
rect 38117 17833 38151 17867
rect 17049 17765 17083 17799
rect 21557 17765 21591 17799
rect 31677 17765 31711 17799
rect 12725 17697 12759 17731
rect 12909 17697 12943 17731
rect 15669 17697 15703 17731
rect 16681 17697 16715 17731
rect 18613 17697 18647 17731
rect 18705 17697 18739 17731
rect 24041 17697 24075 17731
rect 24869 17697 24903 17731
rect 24961 17697 24995 17731
rect 30665 17697 30699 17731
rect 31217 17697 31251 17731
rect 6009 17629 6043 17663
rect 11262 17629 11296 17663
rect 11529 17629 11563 17663
rect 14381 17629 14415 17663
rect 14474 17629 14508 17663
rect 14657 17629 14691 17663
rect 14749 17629 14783 17663
rect 14887 17629 14921 17663
rect 16957 17629 16991 17663
rect 17233 17629 17267 17663
rect 17417 17629 17451 17663
rect 21689 17629 21723 17663
rect 21833 17629 21867 17663
rect 22109 17629 22143 17663
rect 23029 17629 23063 17663
rect 23213 17629 23247 17663
rect 23673 17629 23707 17663
rect 23857 17629 23891 17663
rect 24685 17629 24719 17663
rect 24777 17629 24811 17663
rect 27465 17629 27499 17663
rect 27721 17629 27755 17663
rect 28733 17629 28767 17663
rect 30849 17629 30883 17663
rect 31861 17629 31895 17663
rect 32229 17629 32263 17663
rect 36737 17629 36771 17663
rect 37004 17629 37038 17663
rect 6276 17561 6310 17595
rect 15853 17561 15887 17595
rect 18521 17561 18555 17595
rect 21925 17561 21959 17595
rect 28917 17561 28951 17595
rect 31953 17561 31987 17595
rect 32045 17561 32079 17595
rect 12265 17493 12299 17527
rect 12633 17493 12667 17527
rect 15025 17493 15059 17527
rect 15761 17493 15795 17527
rect 16221 17493 16255 17527
rect 18153 17493 18187 17527
rect 25145 17493 25179 17527
rect 26341 17493 26375 17527
rect 30849 17493 30883 17527
rect 12265 17289 12299 17323
rect 16037 17289 16071 17323
rect 30297 17289 30331 17323
rect 31769 17289 31803 17323
rect 33308 17289 33342 17323
rect 8493 17221 8527 17255
rect 8585 17221 8619 17255
rect 11897 17221 11931 17255
rect 11989 17221 12023 17255
rect 12970 17221 13004 17255
rect 22569 17221 22603 17255
rect 22785 17221 22819 17255
rect 23765 17221 23799 17255
rect 28641 17221 28675 17255
rect 28733 17221 28767 17255
rect 30021 17221 30055 17255
rect 31401 17221 31435 17255
rect 31493 17221 31527 17255
rect 35173 17221 35207 17255
rect 8309 17153 8343 17187
rect 8677 17153 8711 17187
rect 11713 17153 11747 17187
rect 12081 17153 12115 17187
rect 15853 17153 15887 17187
rect 17969 17153 18003 17187
rect 18236 17153 18270 17187
rect 19993 17153 20027 17187
rect 20177 17153 20211 17187
rect 23397 17153 23431 17187
rect 23581 17153 23615 17187
rect 24593 17153 24627 17187
rect 24685 17153 24719 17187
rect 25145 17153 25179 17187
rect 25329 17153 25363 17187
rect 28365 17153 28399 17187
rect 28458 17153 28492 17187
rect 28830 17153 28864 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30113 17153 30147 17187
rect 31217 17153 31251 17187
rect 31585 17153 31619 17187
rect 32873 17153 32907 17187
rect 33425 17153 33459 17187
rect 33701 17153 33735 17187
rect 34621 17153 34655 17187
rect 34897 17153 34931 17187
rect 34989 17153 35023 17187
rect 35725 17153 35759 17187
rect 36001 17153 36035 17187
rect 36093 17153 36127 17187
rect 37841 17153 37875 17187
rect 12725 17085 12759 17119
rect 15577 17085 15611 17119
rect 38117 17085 38151 17119
rect 15669 17017 15703 17051
rect 19349 17017 19383 17051
rect 22937 17017 22971 17051
rect 34713 17017 34747 17051
rect 35817 17017 35851 17051
rect 36277 17017 36311 17051
rect 8861 16949 8895 16983
rect 14105 16949 14139 16983
rect 19809 16949 19843 16983
rect 22753 16949 22787 16983
rect 25605 16949 25639 16983
rect 29009 16949 29043 16983
rect 34897 16745 34931 16779
rect 12909 16677 12943 16711
rect 17233 16677 17267 16711
rect 26709 16677 26743 16711
rect 5641 16609 5675 16643
rect 7665 16609 7699 16643
rect 9137 16609 9171 16643
rect 11529 16609 11563 16643
rect 15853 16609 15887 16643
rect 21281 16609 21315 16643
rect 23489 16609 23523 16643
rect 29837 16609 29871 16643
rect 30297 16609 30331 16643
rect 33609 16609 33643 16643
rect 33885 16609 33919 16643
rect 36737 16609 36771 16643
rect 9393 16541 9427 16575
rect 16120 16541 16154 16575
rect 21465 16541 21499 16575
rect 21925 16541 21959 16575
rect 22017 16541 22051 16575
rect 22385 16541 22419 16575
rect 23213 16541 23247 16575
rect 26157 16541 26191 16575
rect 26341 16541 26375 16575
rect 26525 16541 26559 16575
rect 27353 16541 27387 16575
rect 27445 16541 27479 16575
rect 27721 16541 27755 16575
rect 28181 16541 28215 16575
rect 28365 16541 28399 16575
rect 28549 16541 28583 16575
rect 29745 16541 29779 16575
rect 30021 16541 30055 16575
rect 30113 16541 30147 16575
rect 30941 16541 30975 16575
rect 31125 16541 31159 16575
rect 31309 16541 31343 16575
rect 32045 16541 32079 16575
rect 32193 16541 32227 16575
rect 32321 16541 32355 16575
rect 32413 16541 32447 16575
rect 32510 16541 32544 16575
rect 33517 16541 33551 16575
rect 35076 16541 35110 16575
rect 35393 16541 35427 16575
rect 35541 16541 35575 16575
rect 5908 16473 5942 16507
rect 8401 16473 8435 16507
rect 11796 16473 11830 16507
rect 23397 16473 23431 16507
rect 26433 16473 26467 16507
rect 27537 16473 27571 16507
rect 28457 16473 28491 16507
rect 31217 16473 31251 16507
rect 35173 16473 35207 16507
rect 35265 16473 35299 16507
rect 37004 16473 37038 16507
rect 7021 16405 7055 16439
rect 10517 16405 10551 16439
rect 27169 16405 27203 16439
rect 28733 16405 28767 16439
rect 31493 16405 31527 16439
rect 32689 16405 32723 16439
rect 38117 16405 38151 16439
rect 6561 16201 6595 16235
rect 6929 16201 6963 16235
rect 7021 16201 7055 16235
rect 7941 16201 7975 16235
rect 8953 16201 8987 16235
rect 31033 16201 31067 16235
rect 33517 16201 33551 16235
rect 35817 16201 35851 16235
rect 37473 16201 37507 16235
rect 37933 16201 37967 16235
rect 15945 16133 15979 16167
rect 22661 16133 22695 16167
rect 22877 16133 22911 16167
rect 24317 16133 24351 16167
rect 25973 16133 26007 16167
rect 30481 16133 30515 16167
rect 35541 16133 35575 16167
rect 7882 16065 7916 16099
rect 8309 16065 8343 16099
rect 8861 16065 8895 16099
rect 9045 16065 9079 16099
rect 9781 16065 9815 16099
rect 10048 16065 10082 16099
rect 14289 16065 14323 16099
rect 17233 16065 17267 16099
rect 17325 16065 17359 16099
rect 17509 16065 17543 16099
rect 19717 16065 19751 16099
rect 19984 16065 20018 16099
rect 25697 16065 25731 16099
rect 25789 16065 25823 16099
rect 27261 16065 27295 16099
rect 27353 16065 27387 16099
rect 27445 16065 27479 16099
rect 27537 16065 27571 16099
rect 28825 16065 28859 16099
rect 28917 16065 28951 16099
rect 29009 16065 29043 16099
rect 29101 16065 29135 16099
rect 30389 16065 30423 16099
rect 30757 16065 30791 16099
rect 32321 16065 32355 16099
rect 32413 16065 32447 16099
rect 32597 16065 32631 16099
rect 32689 16065 32723 16099
rect 33333 16065 33367 16099
rect 33701 16065 33735 16099
rect 35173 16065 35207 16099
rect 35266 16065 35300 16099
rect 35403 16065 35437 16099
rect 35638 16065 35672 16099
rect 37841 16065 37875 16099
rect 7205 15997 7239 16031
rect 8401 15997 8435 16031
rect 14565 15997 14599 16031
rect 24225 15997 24259 16031
rect 24409 15997 24443 16031
rect 30849 15997 30883 16031
rect 38025 15997 38059 16031
rect 7757 15861 7791 15895
rect 11161 15861 11195 15895
rect 17693 15861 17727 15895
rect 21097 15861 21131 15895
rect 22845 15861 22879 15895
rect 23029 15861 23063 15895
rect 24777 15861 24811 15895
rect 25973 15861 26007 15895
rect 27721 15861 27755 15895
rect 29285 15861 29319 15895
rect 32873 15861 32907 15895
rect 33701 15861 33735 15895
rect 6469 15657 6503 15691
rect 10425 15657 10459 15691
rect 10793 15657 10827 15691
rect 27169 15657 27203 15691
rect 29101 15657 29135 15691
rect 35633 15657 35667 15691
rect 11805 15589 11839 15623
rect 16865 15589 16899 15623
rect 18521 15589 18555 15623
rect 21465 15589 21499 15623
rect 10885 15521 10919 15555
rect 13001 15521 13035 15555
rect 17601 15521 17635 15555
rect 19625 15521 19659 15555
rect 30389 15521 30423 15555
rect 31493 15521 31527 15555
rect 31677 15521 31711 15555
rect 35449 15521 35483 15555
rect 37841 15521 37875 15555
rect 37933 15521 37967 15555
rect 7593 15453 7627 15487
rect 7849 15453 7883 15487
rect 10609 15453 10643 15487
rect 11805 15453 11839 15487
rect 11897 15453 11931 15487
rect 13737 15453 13771 15487
rect 16129 15453 16163 15487
rect 16221 15453 16255 15487
rect 16957 15453 16991 15487
rect 17877 15453 17911 15487
rect 18613 15453 18647 15487
rect 19441 15453 19475 15487
rect 19717 15453 19751 15487
rect 20545 15453 20579 15487
rect 21644 15453 21678 15487
rect 21741 15453 21775 15487
rect 22017 15453 22051 15487
rect 23029 15453 23063 15487
rect 23305 15453 23339 15487
rect 24869 15453 24903 15487
rect 25053 15453 25087 15487
rect 27077 15453 27111 15487
rect 27261 15453 27295 15487
rect 29009 15453 29043 15487
rect 29193 15453 29227 15487
rect 30573 15453 30607 15487
rect 35357 15453 35391 15487
rect 21833 15385 21867 15419
rect 23397 15385 23431 15419
rect 31401 15385 31435 15419
rect 34989 15385 35023 15419
rect 35081 15385 35115 15419
rect 37749 15385 37783 15419
rect 24961 15317 24995 15351
rect 31033 15317 31067 15351
rect 37381 15317 37415 15351
rect 9965 15113 9999 15147
rect 13921 15113 13955 15147
rect 22092 15113 22126 15147
rect 23949 15113 23983 15147
rect 31769 15113 31803 15147
rect 8953 15045 8987 15079
rect 11989 15045 12023 15079
rect 19257 15045 19291 15079
rect 22477 15045 22511 15079
rect 25697 15045 25731 15079
rect 30656 15045 30690 15079
rect 33241 15045 33275 15079
rect 34866 15045 34900 15079
rect 38117 15045 38151 15079
rect 8125 14977 8159 15011
rect 9873 14977 9907 15011
rect 13553 14977 13587 15011
rect 15945 14977 15979 15011
rect 17141 14977 17175 15011
rect 17233 14977 17267 15011
rect 17325 14977 17359 15011
rect 17509 14977 17543 15011
rect 18889 14977 18923 15011
rect 22241 14977 22275 15011
rect 22385 14977 22419 15011
rect 22661 14977 22695 15011
rect 24133 14977 24167 15011
rect 24409 14977 24443 15011
rect 25421 14977 25455 15011
rect 25605 14977 25639 15011
rect 25841 14977 25875 15011
rect 27353 14977 27387 15011
rect 28365 14977 28399 15011
rect 28549 14977 28583 15011
rect 28641 14977 28675 15011
rect 33609 14977 33643 15011
rect 37841 14977 37875 15011
rect 10057 14909 10091 14943
rect 12725 14909 12759 14943
rect 13461 14909 13495 14943
rect 16129 14909 16163 14943
rect 18429 14909 18463 14943
rect 20361 14909 20395 14943
rect 27169 14909 27203 14943
rect 27721 14909 27755 14943
rect 28181 14909 28215 14943
rect 30389 14909 30423 14943
rect 33333 14909 33367 14943
rect 33701 14909 33735 14943
rect 34621 14909 34655 14943
rect 18061 14841 18095 14875
rect 19993 14841 20027 14875
rect 27629 14841 27663 14875
rect 33885 14841 33919 14875
rect 9505 14773 9539 14807
rect 15761 14773 15795 14807
rect 16865 14773 16899 14807
rect 17969 14773 18003 14807
rect 19901 14773 19935 14807
rect 24317 14773 24351 14807
rect 25973 14773 26007 14807
rect 36001 14773 36035 14807
rect 12725 14569 12759 14603
rect 13277 14569 13311 14603
rect 17233 14569 17267 14603
rect 18705 14569 18739 14603
rect 24869 14569 24903 14603
rect 25237 14569 25271 14603
rect 27169 14569 27203 14603
rect 36093 14569 36127 14603
rect 38301 14569 38335 14603
rect 13369 14501 13403 14535
rect 21465 14501 21499 14535
rect 32965 14501 32999 14535
rect 11529 14433 11563 14467
rect 17877 14433 17911 14467
rect 20177 14433 20211 14467
rect 24961 14433 24995 14467
rect 32689 14433 32723 14467
rect 35449 14433 35483 14467
rect 36921 14433 36955 14467
rect 11621 14365 11655 14399
rect 12633 14365 12667 14399
rect 12817 14365 12851 14399
rect 15301 14365 15335 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 21644 14365 21678 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 23949 14365 23983 14399
rect 24869 14365 24903 14399
rect 27077 14365 27111 14399
rect 35817 14365 35851 14399
rect 35909 14365 35943 14399
rect 37188 14365 37222 14399
rect 12081 14297 12115 14331
rect 13737 14297 13771 14331
rect 15117 14297 15151 14331
rect 15485 14297 15519 14331
rect 17693 14297 17727 14331
rect 23765 14297 23799 14331
rect 35541 14297 35575 14331
rect 17601 14229 17635 14263
rect 19625 14229 19659 14263
rect 19993 14229 20027 14263
rect 20085 14229 20119 14263
rect 23581 14229 23615 14263
rect 33149 14229 33183 14263
rect 9229 14025 9263 14059
rect 12173 14025 12207 14059
rect 17509 14025 17543 14059
rect 23489 14025 23523 14059
rect 25237 14025 25271 14059
rect 8116 13957 8150 13991
rect 13093 13957 13127 13991
rect 16865 13957 16899 13991
rect 19349 13957 19383 13991
rect 22753 13957 22787 13991
rect 25881 13957 25915 13991
rect 26065 13957 26099 13991
rect 27997 13957 28031 13991
rect 28457 13957 28491 13991
rect 7849 13889 7883 13923
rect 10425 13889 10459 13923
rect 11989 13889 12023 13923
rect 13001 13889 13035 13923
rect 13461 13889 13495 13923
rect 14749 13889 14783 13923
rect 15209 13889 15243 13923
rect 15301 13889 15335 13923
rect 17325 13889 17359 13923
rect 18521 13889 18555 13923
rect 18613 13889 18647 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 19625 13889 19659 13923
rect 22661 13889 22695 13923
rect 22937 13889 22971 13923
rect 23765 13889 23799 13923
rect 24041 13889 24075 13923
rect 25053 13889 25087 13923
rect 25789 13889 25823 13923
rect 27721 13889 27755 13923
rect 27813 13889 27847 13923
rect 28825 13889 28859 13923
rect 29009 13889 29043 13923
rect 29469 13889 29503 13923
rect 30021 13889 30055 13923
rect 30113 13889 30147 13923
rect 31125 13889 31159 13923
rect 31309 13889 31343 13923
rect 33241 13889 33275 13923
rect 10517 13821 10551 13855
rect 11805 13821 11839 13855
rect 12909 13821 12943 13855
rect 14381 13821 14415 13855
rect 15025 13821 15059 13855
rect 17233 13821 17267 13855
rect 18245 13821 18279 13855
rect 19533 13821 19567 13855
rect 19993 13821 20027 13855
rect 23627 13821 23661 13855
rect 24133 13821 24167 13855
rect 24593 13821 24627 13855
rect 24961 13821 24995 13855
rect 31033 13821 31067 13855
rect 31769 13821 31803 13855
rect 33333 13821 33367 13855
rect 38301 13821 38335 13855
rect 10793 13753 10827 13787
rect 13921 13753 13955 13787
rect 22937 13753 22971 13787
rect 28825 13753 28859 13787
rect 29929 13753 29963 13787
rect 26065 13685 26099 13719
rect 27997 13685 28031 13719
rect 33517 13685 33551 13719
rect 15485 13481 15519 13515
rect 23489 13481 23523 13515
rect 31217 13481 31251 13515
rect 33057 13481 33091 13515
rect 10517 13413 10551 13447
rect 28641 13413 28675 13447
rect 30297 13413 30331 13447
rect 32965 13413 32999 13447
rect 10241 13345 10275 13379
rect 14381 13345 14415 13379
rect 14933 13345 14967 13379
rect 21741 13345 21775 13379
rect 23673 13345 23707 13379
rect 23765 13345 23799 13379
rect 25053 13345 25087 13379
rect 25605 13345 25639 13379
rect 26065 13345 26099 13379
rect 28457 13345 28491 13379
rect 29837 13345 29871 13379
rect 30849 13345 30883 13379
rect 32597 13345 32631 13379
rect 35725 13345 35759 13379
rect 10149 13277 10183 13311
rect 14565 13277 14599 13311
rect 15853 13277 15887 13311
rect 16129 13277 16163 13311
rect 16221 13277 16255 13311
rect 16497 13277 16531 13311
rect 16773 13277 16807 13311
rect 17325 13277 17359 13311
rect 17509 13277 17543 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 17877 13277 17911 13311
rect 20821 13277 20855 13311
rect 21005 13277 21039 13311
rect 21465 13277 21499 13311
rect 21557 13277 21591 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 25881 13277 25915 13311
rect 27169 13277 27203 13311
rect 27261 13277 27295 13311
rect 27537 13277 27571 13311
rect 27629 13277 27663 13311
rect 28733 13277 28767 13311
rect 29929 13277 29963 13311
rect 30941 13277 30975 13311
rect 33517 13277 33551 13311
rect 33701 13277 33735 13311
rect 35981 13277 36015 13311
rect 20913 13209 20947 13243
rect 26525 13209 26559 13243
rect 14565 13141 14599 13175
rect 21741 13141 21775 13175
rect 28273 13141 28307 13175
rect 33609 13141 33643 13175
rect 37105 13141 37139 13175
rect 12265 12937 12299 12971
rect 13461 12937 13495 12971
rect 23581 12937 23615 12971
rect 28549 12937 28583 12971
rect 35081 12937 35115 12971
rect 15485 12869 15519 12903
rect 15577 12869 15611 12903
rect 22017 12869 22051 12903
rect 7389 12801 7423 12835
rect 7656 12801 7690 12835
rect 9413 12801 9447 12835
rect 12081 12801 12115 12835
rect 12357 12801 12391 12835
rect 13369 12801 13403 12835
rect 13553 12801 13587 12835
rect 15301 12801 15335 12835
rect 17417 12801 17451 12835
rect 21097 12801 21131 12835
rect 21189 12801 21223 12835
rect 21465 12801 21499 12835
rect 22201 12801 22235 12835
rect 22385 12801 22419 12835
rect 22477 12801 22511 12835
rect 23489 12801 23523 12835
rect 23673 12801 23707 12835
rect 25605 12801 25639 12835
rect 25881 12801 25915 12835
rect 27905 12801 27939 12835
rect 27997 12801 28031 12835
rect 28457 12801 28491 12835
rect 28641 12801 28675 12835
rect 33701 12801 33735 12835
rect 33957 12801 33991 12835
rect 9321 12733 9355 12767
rect 9781 12733 9815 12767
rect 17233 12733 17267 12767
rect 25789 12733 25823 12767
rect 27721 12733 27755 12767
rect 8769 12665 8803 12699
rect 15025 12665 15059 12699
rect 21373 12665 21407 12699
rect 12081 12597 12115 12631
rect 17601 12597 17635 12631
rect 20913 12597 20947 12631
rect 25421 12597 25455 12631
rect 27537 12597 27571 12631
rect 38301 12597 38335 12631
rect 10977 12393 11011 12427
rect 14841 12393 14875 12427
rect 16865 12393 16899 12427
rect 18061 12393 18095 12427
rect 20913 12393 20947 12427
rect 25973 12393 26007 12427
rect 27721 12393 27755 12427
rect 13553 12325 13587 12359
rect 14289 12325 14323 12359
rect 16129 12325 16163 12359
rect 19717 12325 19751 12359
rect 9413 12257 9447 12291
rect 14933 12257 14967 12291
rect 15669 12257 15703 12291
rect 17049 12257 17083 12291
rect 17141 12257 17175 12291
rect 17877 12257 17911 12291
rect 21925 12257 21959 12291
rect 25421 12257 25455 12291
rect 31309 12257 31343 12291
rect 32965 12257 32999 12291
rect 35725 12257 35759 12291
rect 9689 12189 9723 12223
rect 11989 12189 12023 12223
rect 12633 12189 12667 12223
rect 13277 12189 13311 12223
rect 14414 12189 14448 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 16405 12189 16439 12223
rect 17233 12189 17267 12223
rect 17325 12189 17359 12223
rect 18153 12189 18187 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 21097 12189 21131 12223
rect 21281 12189 21315 12223
rect 21373 12189 21407 12223
rect 21833 12189 21867 12223
rect 22017 12189 22051 12223
rect 27445 12189 27479 12223
rect 27721 12189 27755 12223
rect 31217 12189 31251 12223
rect 36921 12189 36955 12223
rect 11713 12121 11747 12155
rect 12817 12121 12851 12155
rect 13369 12121 13403 12155
rect 13553 12121 13587 12155
rect 16129 12121 16163 12155
rect 17877 12121 17911 12155
rect 19717 12121 19751 12155
rect 25697 12121 25731 12155
rect 31125 12121 31159 12155
rect 35541 12121 35575 12155
rect 37188 12121 37222 12155
rect 12449 12053 12483 12087
rect 14473 12053 14507 12087
rect 15669 12053 15703 12087
rect 16313 12053 16347 12087
rect 25513 12053 25547 12087
rect 27537 12053 27571 12087
rect 30757 12053 30791 12087
rect 32321 12053 32355 12087
rect 32689 12053 32723 12087
rect 32781 12053 32815 12087
rect 35081 12053 35115 12087
rect 35449 12053 35483 12087
rect 38301 12053 38335 12087
rect 8953 11849 8987 11883
rect 15025 11849 15059 11883
rect 24777 11849 24811 11883
rect 25237 11849 25271 11883
rect 33701 11849 33735 11883
rect 35173 11849 35207 11883
rect 37473 11849 37507 11883
rect 37841 11849 37875 11883
rect 37933 11849 37967 11883
rect 17693 11781 17727 11815
rect 23204 11781 23238 11815
rect 25145 11781 25179 11815
rect 26157 11781 26191 11815
rect 32566 11781 32600 11815
rect 7573 11713 7607 11747
rect 7840 11713 7874 11747
rect 11161 11713 11195 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 12265 11713 12299 11747
rect 13001 11713 13035 11747
rect 14933 11713 14967 11747
rect 17325 11713 17359 11747
rect 17509 11713 17543 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 19349 11713 19383 11747
rect 19441 11713 19475 11747
rect 19699 11713 19733 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 22937 11713 22971 11747
rect 25973 11713 26007 11747
rect 26249 11713 26283 11747
rect 30297 11713 30331 11747
rect 30564 11713 30598 11747
rect 35265 11713 35299 11747
rect 36001 11713 36035 11747
rect 36553 11713 36587 11747
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 12725 11645 12759 11679
rect 15209 11645 15243 11679
rect 20637 11645 20671 11679
rect 25421 11645 25455 11679
rect 32321 11645 32355 11679
rect 35817 11645 35851 11679
rect 36277 11645 36311 11679
rect 38025 11645 38059 11679
rect 11069 11577 11103 11611
rect 12909 11577 12943 11611
rect 14565 11577 14599 11611
rect 18705 11577 18739 11611
rect 19625 11577 19659 11611
rect 24317 11577 24351 11611
rect 25973 11577 26007 11611
rect 10793 11509 10827 11543
rect 11713 11509 11747 11543
rect 12817 11509 12851 11543
rect 19165 11509 19199 11543
rect 20545 11509 20579 11543
rect 31677 11509 31711 11543
rect 10333 11305 10367 11339
rect 19441 11305 19475 11339
rect 20453 11305 20487 11339
rect 21925 11305 21959 11339
rect 25697 11305 25731 11339
rect 25881 11305 25915 11339
rect 36277 11305 36311 11339
rect 27905 11237 27939 11271
rect 32505 11237 32539 11271
rect 17141 11169 17175 11203
rect 17509 11169 17543 11203
rect 17601 11169 17635 11203
rect 18337 11169 18371 11203
rect 22569 11169 22603 11203
rect 28917 11169 28951 11203
rect 29101 11169 29135 11203
rect 29837 11169 29871 11203
rect 30481 11169 30515 11203
rect 32965 11169 32999 11203
rect 34897 11169 34931 11203
rect 10517 11101 10551 11135
rect 10701 11101 10735 11135
rect 10793 11101 10827 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 15853 11101 15887 11135
rect 16037 11101 16071 11135
rect 16681 11101 16715 11135
rect 17325 11101 17359 11135
rect 17417 11101 17451 11135
rect 18245 11101 18279 11135
rect 18429 11101 18463 11135
rect 19625 11101 19659 11135
rect 19809 11101 19843 11135
rect 19901 11101 19935 11135
rect 20361 11101 20395 11135
rect 20545 11101 20579 11135
rect 21557 11101 21591 11135
rect 21833 11101 21867 11135
rect 22753 11101 22787 11135
rect 22845 11101 22879 11135
rect 26525 11101 26559 11135
rect 29745 11101 29779 11135
rect 30665 11101 30699 11135
rect 31033 11101 31067 11135
rect 31585 11101 31619 11135
rect 32229 11101 32263 11135
rect 33149 11101 33183 11135
rect 33425 11101 33459 11135
rect 33517 11101 33551 11135
rect 36829 11101 36863 11135
rect 15945 11033 15979 11067
rect 25513 11033 25547 11067
rect 25713 11033 25747 11067
rect 26792 11033 26826 11067
rect 28825 11033 28859 11067
rect 35164 11033 35198 11067
rect 37096 11033 37130 11067
rect 11805 10965 11839 10999
rect 16589 10965 16623 10999
rect 22109 10965 22143 10999
rect 22569 10965 22603 10999
rect 28457 10965 28491 10999
rect 38209 10965 38243 10999
rect 10149 10761 10183 10795
rect 17233 10761 17267 10795
rect 17693 10761 17727 10795
rect 21189 10761 21223 10795
rect 22017 10761 22051 10795
rect 27169 10761 27203 10795
rect 27537 10761 27571 10795
rect 29745 10761 29779 10795
rect 37473 10761 37507 10795
rect 15117 10693 15151 10727
rect 17601 10693 17635 10727
rect 18889 10693 18923 10727
rect 21097 10693 21131 10727
rect 22293 10693 22327 10727
rect 22385 10693 22419 10727
rect 27629 10693 27663 10727
rect 28610 10693 28644 10727
rect 37933 10693 37967 10727
rect 8769 10625 8803 10659
rect 13645 10625 13679 10659
rect 13829 10625 13863 10659
rect 15301 10625 15335 10659
rect 22201 10625 22235 10659
rect 22569 10625 22603 10659
rect 24409 10625 24443 10659
rect 24676 10625 24710 10659
rect 28365 10625 28399 10659
rect 34161 10625 34195 10659
rect 37841 10625 37875 10659
rect 9045 10557 9079 10591
rect 15669 10557 15703 10591
rect 17877 10557 17911 10591
rect 18429 10557 18463 10591
rect 21373 10557 21407 10591
rect 27813 10557 27847 10591
rect 34253 10557 34287 10591
rect 34437 10557 34471 10591
rect 38025 10557 38059 10591
rect 18613 10489 18647 10523
rect 13461 10421 13495 10455
rect 13645 10421 13679 10455
rect 20729 10421 20763 10455
rect 25789 10421 25823 10455
rect 33793 10421 33827 10455
rect 10333 10217 10367 10251
rect 11161 10217 11195 10251
rect 17509 10217 17543 10251
rect 21833 10217 21867 10251
rect 24777 10217 24811 10251
rect 31769 10217 31803 10251
rect 14841 10149 14875 10183
rect 34345 10149 34379 10183
rect 35173 10149 35207 10183
rect 10701 10081 10735 10115
rect 12081 10081 12115 10115
rect 15485 10081 15519 10115
rect 17693 10081 17727 10115
rect 17785 10081 17819 10115
rect 18153 10081 18187 10115
rect 20361 10081 20395 10115
rect 25237 10081 25271 10115
rect 25421 10081 25455 10115
rect 35817 10081 35851 10115
rect 36277 10081 36311 10115
rect 38117 10081 38151 10115
rect 10517 10013 10551 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 12357 10013 12391 10047
rect 13737 10013 13771 10047
rect 15209 10013 15243 10047
rect 16037 10013 16071 10047
rect 16221 10013 16255 10047
rect 20177 10013 20211 10047
rect 20453 10013 20487 10047
rect 20913 10013 20947 10047
rect 21097 10013 21131 10047
rect 21741 10013 21775 10047
rect 21925 10013 21959 10047
rect 25145 10013 25179 10047
rect 32045 10013 32079 10047
rect 32137 10013 32171 10047
rect 32229 10013 32263 10047
rect 32413 10013 32447 10047
rect 32965 10013 32999 10047
rect 33232 10013 33266 10047
rect 35265 10013 35299 10047
rect 36001 10013 36035 10047
rect 36553 10013 36587 10047
rect 37841 10013 37875 10047
rect 16129 9945 16163 9979
rect 11529 9877 11563 9911
rect 15301 9877 15335 9911
rect 19993 9877 20027 9911
rect 21005 9877 21039 9911
rect 10885 9673 10919 9707
rect 13369 9673 13403 9707
rect 15301 9673 15335 9707
rect 20729 9673 20763 9707
rect 32689 9673 32723 9707
rect 34989 9673 35023 9707
rect 10425 9605 10459 9639
rect 11989 9605 12023 9639
rect 14013 9605 14047 9639
rect 14197 9605 14231 9639
rect 15393 9605 15427 9639
rect 19073 9605 19107 9639
rect 21189 9605 21223 9639
rect 24869 9605 24903 9639
rect 25605 9605 25639 9639
rect 29653 9605 29687 9639
rect 30113 9605 30147 9639
rect 38117 9605 38151 9639
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 11161 9537 11195 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 12909 9537 12943 9571
rect 13829 9537 13863 9571
rect 17049 9537 17083 9571
rect 19165 9537 19199 9571
rect 21097 9537 21131 9571
rect 22569 9537 22603 9571
rect 22836 9537 22870 9571
rect 24777 9537 24811 9571
rect 25881 9537 25915 9571
rect 27169 9537 27203 9571
rect 27436 9537 27470 9571
rect 29009 9537 29043 9571
rect 29193 9537 29227 9571
rect 29285 9537 29319 9571
rect 29377 9537 29411 9571
rect 30573 9537 30607 9571
rect 30665 9537 30699 9571
rect 34345 9537 34379 9571
rect 34529 9537 34563 9571
rect 37841 9537 37875 9571
rect 13001 9469 13035 9503
rect 15577 9469 15611 9503
rect 18981 9469 19015 9503
rect 21373 9469 21407 9503
rect 25053 9469 25087 9503
rect 25605 9469 25639 9503
rect 32781 9469 32815 9503
rect 32873 9469 32907 9503
rect 11713 9401 11747 9435
rect 24409 9401 24443 9435
rect 11069 9333 11103 9367
rect 12725 9333 12759 9367
rect 14933 9333 14967 9367
rect 16957 9333 16991 9367
rect 19533 9333 19567 9367
rect 23949 9333 23983 9367
rect 25789 9333 25823 9367
rect 28549 9333 28583 9367
rect 32321 9333 32355 9367
rect 25329 9129 25363 9163
rect 30021 9129 30055 9163
rect 20821 9061 20855 9095
rect 32321 9061 32355 9095
rect 35633 9061 35667 9095
rect 16405 8993 16439 9027
rect 19993 8993 20027 9027
rect 21189 8993 21223 9027
rect 21373 8993 21407 9027
rect 27261 8993 27295 9027
rect 33057 8993 33091 9027
rect 36277 8993 36311 9027
rect 36737 8993 36771 9027
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15393 8925 15427 8959
rect 15577 8925 15611 8959
rect 15761 8925 15795 8959
rect 16497 8925 16531 8959
rect 17601 8925 17635 8959
rect 18705 8925 18739 8959
rect 18889 8925 18923 8959
rect 19441 8925 19475 8959
rect 19809 8925 19843 8959
rect 24869 8925 24903 8959
rect 24961 8925 24995 8959
rect 25145 8925 25179 8959
rect 26709 8925 26743 8959
rect 28089 8925 28123 8959
rect 30205 8925 30239 8959
rect 30481 8925 30515 8959
rect 30941 8925 30975 8959
rect 33885 8925 33919 8959
rect 35541 8925 35575 8959
rect 36369 8925 36403 8959
rect 37013 8925 37047 8959
rect 37841 8925 37875 8959
rect 14381 8857 14415 8891
rect 16589 8857 16623 8891
rect 17509 8857 17543 8891
rect 18337 8857 18371 8891
rect 19533 8857 19567 8891
rect 21281 8857 21315 8891
rect 25881 8857 25915 8891
rect 30297 8857 30331 8891
rect 31208 8857 31242 8891
rect 38117 8857 38151 8891
rect 16957 8789 16991 8823
rect 12081 8585 12115 8619
rect 25697 8585 25731 8619
rect 27537 8585 27571 8619
rect 27905 8585 27939 8619
rect 36369 8585 36403 8619
rect 37841 8585 37875 8619
rect 12633 8517 12667 8551
rect 19809 8517 19843 8551
rect 19993 8517 20027 8551
rect 20637 8517 20671 8551
rect 31309 8517 31343 8551
rect 33793 8517 33827 8551
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 14105 8449 14139 8483
rect 14381 8449 14415 8483
rect 15945 8449 15979 8483
rect 16037 8449 16071 8483
rect 16221 8449 16255 8483
rect 16313 8449 16347 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 18337 8449 18371 8483
rect 18889 8449 18923 8483
rect 20821 8449 20855 8483
rect 24584 8449 24618 8483
rect 27997 8449 28031 8483
rect 29193 8449 29227 8483
rect 29285 8449 29319 8483
rect 30481 8449 30515 8483
rect 30757 8449 30791 8483
rect 33057 8449 33091 8483
rect 34989 8449 35023 8483
rect 35256 8449 35290 8483
rect 18521 8381 18555 8415
rect 19625 8381 19659 8415
rect 24317 8381 24351 8415
rect 28089 8381 28123 8415
rect 37933 8381 37967 8415
rect 38025 8381 38059 8415
rect 12541 8313 12575 8347
rect 14013 8313 14047 8347
rect 17325 8313 17359 8347
rect 20453 8313 20487 8347
rect 29469 8313 29503 8347
rect 37473 8313 37507 8347
rect 15761 8245 15795 8279
rect 29009 8245 29043 8279
rect 15577 8041 15611 8075
rect 16221 8041 16255 8075
rect 22937 8041 22971 8075
rect 24869 8041 24903 8075
rect 28641 8041 28675 8075
rect 33885 8041 33919 8075
rect 35265 8041 35299 8075
rect 38301 8041 38335 8075
rect 14473 7973 14507 8007
rect 32229 7973 32263 8007
rect 10609 7905 10643 7939
rect 12265 7905 12299 7939
rect 25329 7905 25363 7939
rect 25513 7905 25547 7939
rect 29745 7905 29779 7939
rect 30297 7905 30331 7939
rect 33241 7905 33275 7939
rect 35725 7905 35759 7939
rect 35817 7905 35851 7939
rect 10885 7837 10919 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 14289 7837 14323 7871
rect 14933 7837 14967 7871
rect 16313 7837 16347 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 20085 7837 20119 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 20821 7837 20855 7871
rect 21557 7837 21591 7871
rect 25237 7837 25271 7871
rect 26433 7837 26467 7871
rect 28273 7837 28307 7871
rect 30205 7837 30239 7871
rect 30849 7837 30883 7871
rect 33057 7837 33091 7871
rect 34069 7837 34103 7871
rect 34253 7837 34287 7871
rect 35633 7837 35667 7871
rect 36921 7837 36955 7871
rect 37188 7837 37222 7871
rect 21824 7769 21858 7803
rect 26700 7769 26734 7803
rect 28457 7769 28491 7803
rect 31116 7769 31150 7803
rect 33149 7769 33183 7803
rect 18153 7701 18187 7735
rect 27813 7701 27847 7735
rect 32689 7701 32723 7735
rect 11805 7497 11839 7531
rect 12173 7497 12207 7531
rect 21097 7497 21131 7531
rect 22017 7497 22051 7531
rect 24159 7497 24193 7531
rect 27169 7497 27203 7531
rect 27537 7497 27571 7531
rect 23949 7429 23983 7463
rect 27629 7429 27663 7463
rect 32956 7429 32990 7463
rect 35357 7429 35391 7463
rect 11989 7361 12023 7395
rect 12265 7361 12299 7395
rect 13737 7361 13771 7395
rect 14105 7361 14139 7395
rect 14473 7361 14507 7395
rect 15668 7361 15702 7395
rect 15761 7361 15795 7395
rect 18245 7361 18279 7395
rect 18521 7361 18555 7395
rect 18889 7361 18923 7395
rect 20177 7361 20211 7395
rect 20269 7361 20303 7395
rect 21005 7361 21039 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 32689 7361 32723 7395
rect 34713 7361 34747 7395
rect 34897 7361 34931 7395
rect 34989 7361 35023 7395
rect 35081 7361 35115 7395
rect 37841 7361 37875 7395
rect 13369 7293 13403 7327
rect 14657 7293 14691 7327
rect 18429 7293 18463 7327
rect 20453 7293 20487 7327
rect 20545 7293 20579 7327
rect 27813 7293 27847 7327
rect 38117 7293 38151 7327
rect 19257 7225 19291 7259
rect 15577 7157 15611 7191
rect 19993 7157 20027 7191
rect 24133 7157 24167 7191
rect 24317 7157 24351 7191
rect 34069 7157 34103 7191
rect 14289 6953 14323 6987
rect 18245 6953 18279 6987
rect 21465 6953 21499 6987
rect 23673 6953 23707 6987
rect 26433 6953 26467 6987
rect 33149 6953 33183 6987
rect 38117 6953 38151 6987
rect 15669 6817 15703 6851
rect 17877 6817 17911 6851
rect 25881 6817 25915 6851
rect 27537 6817 27571 6851
rect 29745 6817 29779 6851
rect 33701 6817 33735 6851
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 14841 6749 14875 6783
rect 15853 6749 15887 6783
rect 16497 6749 16531 6783
rect 18061 6749 18095 6783
rect 18337 6749 18371 6783
rect 19993 6749 20027 6783
rect 20637 6749 20671 6783
rect 20729 6749 20763 6783
rect 22293 6749 22327 6783
rect 24685 6749 24719 6783
rect 26985 6749 27019 6783
rect 27077 6749 27111 6783
rect 30205 6749 30239 6783
rect 30389 6749 30423 6783
rect 30481 6749 30515 6783
rect 36737 6749 36771 6783
rect 21281 6681 21315 6715
rect 22560 6681 22594 6715
rect 25237 6681 25271 6715
rect 26157 6681 26191 6715
rect 33517 6681 33551 6715
rect 37004 6681 37038 6715
rect 16497 6613 16531 6647
rect 21481 6613 21515 6647
rect 21649 6613 21683 6647
rect 25973 6613 26007 6647
rect 33609 6613 33643 6647
rect 23213 6409 23247 6443
rect 23581 6409 23615 6443
rect 24507 6409 24541 6443
rect 28733 6409 28767 6443
rect 29561 6409 29595 6443
rect 29929 6409 29963 6443
rect 30389 6409 30423 6443
rect 34345 6409 34379 6443
rect 35449 6409 35483 6443
rect 37473 6409 37507 6443
rect 37841 6409 37875 6443
rect 37933 6409 37967 6443
rect 24409 6341 24443 6375
rect 34161 6341 34195 6375
rect 15485 6273 15519 6307
rect 18061 6273 18095 6307
rect 18521 6273 18555 6307
rect 20361 6273 20395 6307
rect 21097 6273 21131 6307
rect 22017 6273 22051 6307
rect 22201 6273 22235 6307
rect 24593 6273 24627 6307
rect 24685 6273 24719 6307
rect 25973 6273 26007 6307
rect 26157 6273 26191 6307
rect 26249 6273 26283 6307
rect 27353 6273 27387 6307
rect 27620 6273 27654 6307
rect 29469 6273 29503 6307
rect 30757 6273 30791 6307
rect 33977 6273 34011 6307
rect 34805 6273 34839 6307
rect 34989 6273 35023 6307
rect 35081 6273 35115 6307
rect 35173 6273 35207 6307
rect 15577 6205 15611 6239
rect 16221 6205 16255 6239
rect 20085 6205 20119 6239
rect 23673 6205 23707 6239
rect 23857 6205 23891 6239
rect 29377 6205 29411 6239
rect 30849 6205 30883 6239
rect 31033 6205 31067 6239
rect 38025 6205 38059 6239
rect 20821 6137 20855 6171
rect 22017 6069 22051 6103
rect 25789 6069 25823 6103
rect 22109 5865 22143 5899
rect 25329 5865 25363 5899
rect 25421 5865 25455 5899
rect 27905 5865 27939 5899
rect 35541 5865 35575 5899
rect 19533 5797 19567 5831
rect 17325 5729 17359 5763
rect 17601 5729 17635 5763
rect 18153 5729 18187 5763
rect 19901 5729 19935 5763
rect 20729 5729 20763 5763
rect 25513 5729 25547 5763
rect 28365 5729 28399 5763
rect 28457 5729 28491 5763
rect 33057 5729 33091 5763
rect 33149 5729 33183 5763
rect 17049 5661 17083 5695
rect 17785 5661 17819 5695
rect 21005 5661 21039 5695
rect 25237 5661 25271 5695
rect 28273 5661 28307 5695
rect 30205 5661 30239 5695
rect 32965 5661 32999 5695
rect 33977 5661 34011 5695
rect 34161 5661 34195 5695
rect 34897 5661 34931 5695
rect 35081 5661 35115 5695
rect 35173 5661 35207 5695
rect 35265 5661 35299 5695
rect 37841 5661 37875 5695
rect 30472 5593 30506 5627
rect 33793 5593 33827 5627
rect 38117 5593 38151 5627
rect 19441 5525 19475 5559
rect 31585 5525 31619 5559
rect 32597 5525 32631 5559
rect 23581 5321 23615 5355
rect 30389 5321 30423 5355
rect 30757 5321 30791 5355
rect 33701 5321 33735 5355
rect 34529 5321 34563 5355
rect 36461 5321 36495 5355
rect 37841 5321 37875 5355
rect 17141 5253 17175 5287
rect 20913 5253 20947 5287
rect 34161 5253 34195 5287
rect 37933 5253 37967 5287
rect 18797 5185 18831 5219
rect 19257 5185 19291 5219
rect 22468 5185 22502 5219
rect 24869 5185 24903 5219
rect 30849 5185 30883 5219
rect 32321 5185 32355 5219
rect 32588 5185 32622 5219
rect 34345 5185 34379 5219
rect 35081 5185 35115 5219
rect 35348 5185 35382 5219
rect 18521 5117 18555 5151
rect 19533 5117 19567 5151
rect 22201 5117 22235 5151
rect 24961 5117 24995 5151
rect 25053 5117 25087 5151
rect 31033 5117 31067 5151
rect 38025 5117 38059 5151
rect 24501 4981 24535 5015
rect 37473 4981 37507 5015
rect 17785 4777 17819 4811
rect 23029 4777 23063 4811
rect 31125 4777 31159 4811
rect 34345 4777 34379 4811
rect 35541 4777 35575 4811
rect 38209 4777 38243 4811
rect 25973 4709 26007 4743
rect 26433 4709 26467 4743
rect 16221 4641 16255 4675
rect 16497 4641 16531 4675
rect 23673 4641 23707 4675
rect 28733 4641 28767 4675
rect 28917 4641 28951 4675
rect 29745 4641 29779 4675
rect 32965 4641 32999 4675
rect 36093 4641 36127 4675
rect 36829 4641 36863 4675
rect 24593 4573 24627 4607
rect 24849 4573 24883 4607
rect 27813 4573 27847 4607
rect 28641 4573 28675 4607
rect 35909 4573 35943 4607
rect 37096 4573 37130 4607
rect 23397 4505 23431 4539
rect 27546 4505 27580 4539
rect 30012 4505 30046 4539
rect 33232 4505 33266 4539
rect 36001 4505 36035 4539
rect 23489 4437 23523 4471
rect 28273 4437 28307 4471
rect 26157 4233 26191 4267
rect 26525 4233 26559 4267
rect 28917 4233 28951 4267
rect 30113 4233 30147 4267
rect 30481 4233 30515 4267
rect 33425 4233 33459 4267
rect 33793 4233 33827 4267
rect 27804 4165 27838 4199
rect 30573 4165 30607 4199
rect 26065 4097 26099 4131
rect 27537 4097 27571 4131
rect 33885 4097 33919 4131
rect 37841 4097 37875 4131
rect 38117 4097 38151 4131
rect 25881 4029 25915 4063
rect 30757 4029 30791 4063
rect 33977 4029 34011 4063
rect 37841 3009 37875 3043
rect 38117 2941 38151 2975
rect 37841 2397 37875 2431
rect 38117 2329 38151 2363
<< metal1 >>
rect 5074 39108 5080 39160
rect 5132 39148 5138 39160
rect 6638 39148 6644 39160
rect 5132 39120 6644 39148
rect 5132 39108 5138 39120
rect 6638 39108 6644 39120
rect 6696 39108 6702 39160
rect 21634 39108 21640 39160
rect 21692 39148 21698 39160
rect 22094 39148 22100 39160
rect 21692 39120 22100 39148
rect 21692 39108 21698 39120
rect 22094 39108 22100 39120
rect 22152 39108 22158 39160
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 5810 37272 5816 37324
rect 5868 37272 5874 37324
rect 9306 37272 9312 37324
rect 9364 37312 9370 37324
rect 9677 37315 9735 37321
rect 9677 37312 9689 37315
rect 9364 37284 9689 37312
rect 9364 37272 9370 37284
rect 9677 37281 9689 37284
rect 9723 37281 9735 37315
rect 9677 37275 9735 37281
rect 36630 37272 36636 37324
rect 36688 37312 36694 37324
rect 39022 37312 39028 37324
rect 36688 37284 39028 37312
rect 36688 37272 36694 37284
rect 39022 37272 39028 37284
rect 39080 37272 39086 37324
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 1949 37247 2007 37253
rect 1949 37244 1961 37247
rect 1820 37216 1961 37244
rect 1820 37204 1826 37216
rect 1949 37213 1961 37216
rect 1995 37213 2007 37247
rect 1949 37207 2007 37213
rect 6638 37204 6644 37256
rect 6696 37204 6702 37256
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 8481 37247 8539 37253
rect 8481 37244 8493 37247
rect 8444 37216 8493 37244
rect 8444 37204 8450 37216
rect 8481 37213 8493 37216
rect 8527 37213 8539 37247
rect 8481 37207 8539 37213
rect 11698 37204 11704 37256
rect 11756 37244 11762 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11756 37216 11897 37244
rect 11756 37204 11762 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 15194 37204 15200 37256
rect 15252 37204 15258 37256
rect 18233 37247 18291 37253
rect 18233 37213 18245 37247
rect 18279 37244 18291 37247
rect 18322 37244 18328 37256
rect 18279 37216 18328 37244
rect 18279 37213 18291 37216
rect 18233 37207 18291 37213
rect 18322 37204 18328 37216
rect 18380 37204 18386 37256
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 2501 37179 2559 37185
rect 2501 37145 2513 37179
rect 2547 37176 2559 37179
rect 5534 37176 5540 37188
rect 2547 37148 5540 37176
rect 2547 37145 2559 37148
rect 2501 37139 2559 37145
rect 5534 37136 5540 37148
rect 5592 37136 5598 37188
rect 7006 37136 7012 37188
rect 7064 37136 7070 37188
rect 7374 37136 7380 37188
rect 7432 37176 7438 37188
rect 7929 37179 7987 37185
rect 7929 37176 7941 37179
rect 7432 37148 7941 37176
rect 7432 37136 7438 37148
rect 7929 37145 7941 37148
rect 7975 37145 7987 37179
rect 7929 37139 7987 37145
rect 9493 37179 9551 37185
rect 9493 37145 9505 37179
rect 9539 37176 9551 37179
rect 9674 37176 9680 37188
rect 9539 37148 9680 37176
rect 9539 37145 9551 37148
rect 9493 37139 9551 37145
rect 9674 37136 9680 37148
rect 9732 37176 9738 37188
rect 9732 37148 10732 37176
rect 9732 37136 9738 37148
rect 5166 37068 5172 37120
rect 5224 37068 5230 37120
rect 5626 37068 5632 37120
rect 5684 37068 5690 37120
rect 9122 37068 9128 37120
rect 9180 37068 9186 37120
rect 9582 37068 9588 37120
rect 9640 37068 9646 37120
rect 10704 37108 10732 37148
rect 12066 37136 12072 37188
rect 12124 37176 12130 37188
rect 12253 37179 12311 37185
rect 12253 37176 12265 37179
rect 12124 37148 12265 37176
rect 12124 37136 12130 37148
rect 12253 37145 12265 37148
rect 12299 37145 12311 37179
rect 12253 37139 12311 37145
rect 15749 37179 15807 37185
rect 15749 37145 15761 37179
rect 15795 37176 15807 37179
rect 16206 37176 16212 37188
rect 15795 37148 16212 37176
rect 15795 37145 15807 37148
rect 15749 37139 15807 37145
rect 16206 37136 16212 37148
rect 16264 37136 16270 37188
rect 18782 37176 18788 37188
rect 16960 37148 18788 37176
rect 16960 37108 16988 37148
rect 18782 37136 18788 37148
rect 18840 37136 18846 37188
rect 19628 37176 19656 37207
rect 20162 37204 20168 37256
rect 20220 37204 20226 37256
rect 22094 37204 22100 37256
rect 22152 37204 22158 37256
rect 24946 37204 24952 37256
rect 25004 37244 25010 37256
rect 25041 37247 25099 37253
rect 25041 37244 25053 37247
rect 25004 37216 25053 37244
rect 25004 37204 25010 37216
rect 25041 37213 25053 37216
rect 25087 37213 25099 37247
rect 25041 37207 25099 37213
rect 27154 37204 27160 37256
rect 27212 37204 27218 37256
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 27706 37244 27712 37256
rect 27387 37216 27712 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 28316 37216 28457 37244
rect 28316 37204 28322 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 28445 37207 28503 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 31812 37216 32505 37244
rect 31812 37204 31818 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 36906 37204 36912 37256
rect 36964 37204 36970 37256
rect 38194 37204 38200 37256
rect 38252 37204 38258 37256
rect 18892 37148 19656 37176
rect 10704 37080 16988 37108
rect 17034 37068 17040 37120
rect 17092 37108 17098 37120
rect 18892 37108 18920 37148
rect 17092 37080 18920 37108
rect 17092 37068 17098 37080
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 19484 37080 19533 37108
rect 19484 37068 19490 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 19628 37108 19656 37148
rect 20441 37179 20499 37185
rect 20441 37145 20453 37179
rect 20487 37176 20499 37179
rect 20990 37176 20996 37188
rect 20487 37148 20996 37176
rect 20487 37145 20499 37148
rect 20441 37139 20499 37145
rect 20990 37136 20996 37148
rect 21048 37136 21054 37188
rect 22278 37136 22284 37188
rect 22336 37176 22342 37188
rect 22833 37179 22891 37185
rect 22833 37176 22845 37179
rect 22336 37148 22845 37176
rect 22336 37136 22342 37148
rect 22833 37145 22845 37148
rect 22879 37145 22891 37179
rect 22833 37139 22891 37145
rect 22922 37136 22928 37188
rect 22980 37176 22986 37188
rect 25869 37179 25927 37185
rect 25869 37176 25881 37179
rect 22980 37148 25881 37176
rect 22980 37136 22986 37148
rect 25869 37145 25881 37148
rect 25915 37176 25927 37179
rect 31018 37176 31024 37188
rect 25915 37148 31024 37176
rect 25915 37145 25927 37148
rect 25869 37139 25927 37145
rect 31018 37136 31024 37148
rect 31076 37136 31082 37188
rect 31846 37136 31852 37188
rect 31904 37176 31910 37188
rect 32309 37179 32367 37185
rect 32309 37176 32321 37179
rect 31904 37148 32321 37176
rect 31904 37136 31910 37148
rect 32309 37145 32321 37148
rect 32355 37145 32367 37179
rect 32309 37139 32367 37145
rect 36633 37179 36691 37185
rect 36633 37145 36645 37179
rect 36679 37145 36691 37179
rect 36633 37139 36691 37145
rect 23658 37108 23664 37120
rect 19628 37080 23664 37108
rect 19521 37071 19579 37077
rect 23658 37068 23664 37080
rect 23716 37068 23722 37120
rect 26602 37068 26608 37120
rect 26660 37108 26666 37120
rect 27157 37111 27215 37117
rect 27157 37108 27169 37111
rect 26660 37080 27169 37108
rect 26660 37068 26666 37080
rect 27157 37077 27169 37080
rect 27203 37077 27215 37111
rect 27157 37071 27215 37077
rect 28534 37068 28540 37120
rect 28592 37068 28598 37120
rect 36648 37108 36676 37139
rect 36814 37136 36820 37188
rect 36872 37176 36878 37188
rect 37645 37179 37703 37185
rect 37645 37176 37657 37179
rect 36872 37148 37657 37176
rect 36872 37136 36878 37148
rect 37645 37145 37657 37148
rect 37691 37145 37703 37179
rect 37645 37139 37703 37145
rect 39022 37108 39028 37120
rect 36648 37080 39028 37108
rect 39022 37068 39028 37080
rect 39080 37068 39086 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 5626 36864 5632 36916
rect 5684 36904 5690 36916
rect 5997 36907 6055 36913
rect 5997 36904 6009 36907
rect 5684 36876 6009 36904
rect 5684 36864 5690 36876
rect 5997 36873 6009 36876
rect 6043 36873 6055 36907
rect 5997 36867 6055 36873
rect 9582 36864 9588 36916
rect 9640 36864 9646 36916
rect 11054 36864 11060 36916
rect 11112 36904 11118 36916
rect 14182 36904 14188 36916
rect 11112 36876 14188 36904
rect 11112 36864 11118 36876
rect 14182 36864 14188 36876
rect 14240 36864 14246 36916
rect 24121 36907 24179 36913
rect 24121 36904 24133 36907
rect 14292 36876 15976 36904
rect 4884 36839 4942 36845
rect 4884 36805 4896 36839
rect 4930 36836 4942 36839
rect 5166 36836 5172 36848
rect 4930 36808 5172 36836
rect 4930 36805 4942 36808
rect 4884 36799 4942 36805
rect 5166 36796 5172 36808
rect 5224 36796 5230 36848
rect 8472 36839 8530 36845
rect 8472 36805 8484 36839
rect 8518 36836 8530 36839
rect 9122 36836 9128 36848
rect 8518 36808 9128 36836
rect 8518 36805 8530 36808
rect 8472 36799 8530 36805
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 13170 36728 13176 36780
rect 13228 36777 13234 36780
rect 13228 36731 13240 36777
rect 13228 36728 13234 36731
rect 13354 36728 13360 36780
rect 13412 36768 13418 36780
rect 14292 36777 14320 36876
rect 15948 36848 15976 36876
rect 17788 36876 22140 36904
rect 15194 36796 15200 36848
rect 15252 36796 15258 36848
rect 15930 36796 15936 36848
rect 15988 36836 15994 36848
rect 17788 36836 17816 36876
rect 19426 36836 19432 36848
rect 15988 36808 17816 36836
rect 19274 36808 19432 36836
rect 15988 36796 15994 36808
rect 13449 36771 13507 36777
rect 13449 36768 13461 36771
rect 13412 36740 13461 36768
rect 13412 36728 13418 36740
rect 13449 36737 13461 36740
rect 13495 36768 13507 36771
rect 14277 36771 14335 36777
rect 14277 36768 14289 36771
rect 13495 36740 14289 36768
rect 13495 36737 13507 36740
rect 13449 36731 13507 36737
rect 14277 36737 14289 36740
rect 14323 36737 14335 36771
rect 14277 36731 14335 36737
rect 17034 36728 17040 36780
rect 17092 36728 17098 36780
rect 17788 36777 17816 36808
rect 19426 36796 19432 36808
rect 19484 36796 19490 36848
rect 17773 36771 17831 36777
rect 17773 36737 17785 36771
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 20622 36728 20628 36780
rect 20680 36728 20686 36780
rect 20990 36728 20996 36780
rect 21048 36768 21054 36780
rect 21542 36768 21548 36780
rect 21048 36740 21548 36768
rect 21048 36728 21054 36740
rect 21542 36728 21548 36740
rect 21600 36728 21606 36780
rect 22112 36777 22140 36876
rect 22204 36876 24133 36904
rect 22097 36771 22155 36777
rect 22097 36737 22109 36771
rect 22143 36737 22155 36771
rect 22097 36731 22155 36737
rect 4614 36660 4620 36712
rect 4672 36660 4678 36712
rect 8205 36703 8263 36709
rect 8205 36669 8217 36703
rect 8251 36669 8263 36703
rect 8205 36663 8263 36669
rect 8220 36564 8248 36663
rect 14550 36660 14556 36712
rect 14608 36660 14614 36712
rect 15102 36660 15108 36712
rect 15160 36700 15166 36712
rect 17052 36700 17080 36728
rect 15160 36672 17080 36700
rect 15160 36660 15166 36672
rect 18046 36660 18052 36712
rect 18104 36660 18110 36712
rect 19978 36660 19984 36712
rect 20036 36660 20042 36712
rect 20640 36700 20668 36728
rect 22204 36700 22232 36876
rect 24121 36873 24133 36876
rect 24167 36873 24179 36907
rect 26513 36907 26571 36913
rect 26513 36904 26525 36907
rect 24121 36867 24179 36873
rect 24320 36876 26525 36904
rect 23750 36796 23756 36848
rect 23808 36836 23814 36848
rect 24320 36836 24348 36876
rect 26513 36873 26525 36876
rect 26559 36873 26571 36907
rect 26513 36867 26571 36873
rect 25590 36836 25596 36848
rect 23808 36808 24348 36836
rect 25162 36808 25596 36836
rect 23808 36796 23814 36808
rect 25590 36796 25596 36808
rect 25648 36796 25654 36848
rect 28810 36836 28816 36848
rect 27540 36808 28816 36836
rect 22370 36777 22376 36780
rect 22364 36731 22376 36777
rect 22370 36728 22376 36731
rect 22428 36728 22434 36780
rect 26326 36728 26332 36780
rect 26384 36728 26390 36780
rect 26602 36728 26608 36780
rect 26660 36728 26666 36780
rect 27540 36777 27568 36808
rect 28810 36796 28816 36808
rect 28868 36836 28874 36848
rect 32766 36836 32772 36848
rect 28868 36808 31064 36836
rect 28868 36796 28874 36808
rect 27525 36771 27583 36777
rect 27525 36737 27537 36771
rect 27571 36737 27583 36771
rect 27525 36731 27583 36737
rect 27792 36771 27850 36777
rect 27792 36737 27804 36771
rect 27838 36768 27850 36771
rect 28258 36768 28264 36780
rect 27838 36740 28264 36768
rect 27838 36737 27850 36740
rect 27792 36731 27850 36737
rect 20640 36672 22232 36700
rect 24854 36660 24860 36712
rect 24912 36700 24918 36712
rect 25593 36703 25651 36709
rect 25593 36700 25605 36703
rect 24912 36672 25605 36700
rect 24912 36660 24918 36672
rect 25593 36669 25605 36672
rect 25639 36669 25651 36703
rect 25593 36663 25651 36669
rect 25869 36703 25927 36709
rect 25869 36669 25881 36703
rect 25915 36700 25927 36703
rect 26142 36700 26148 36712
rect 25915 36672 26148 36700
rect 25915 36669 25927 36672
rect 25869 36663 25927 36669
rect 26142 36660 26148 36672
rect 26200 36700 26206 36712
rect 27540 36700 27568 36731
rect 28258 36728 28264 36740
rect 28316 36728 28322 36780
rect 31036 36777 31064 36808
rect 32324 36808 32772 36836
rect 32324 36777 32352 36808
rect 32766 36796 32772 36808
rect 32824 36796 32830 36848
rect 30765 36771 30823 36777
rect 30765 36737 30777 36771
rect 30811 36768 30823 36771
rect 31021 36771 31079 36777
rect 30811 36740 30972 36768
rect 30811 36737 30823 36740
rect 30765 36731 30823 36737
rect 26200 36672 27568 36700
rect 30944 36700 30972 36740
rect 31021 36737 31033 36771
rect 31067 36768 31079 36771
rect 32309 36771 32367 36777
rect 32309 36768 32321 36771
rect 31067 36740 32321 36768
rect 31067 36737 31079 36740
rect 31021 36731 31079 36737
rect 32309 36737 32321 36740
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 32398 36728 32404 36780
rect 32456 36768 32462 36780
rect 32565 36771 32623 36777
rect 32565 36768 32577 36771
rect 32456 36740 32577 36768
rect 32456 36728 32462 36740
rect 32565 36737 32577 36740
rect 32611 36737 32623 36771
rect 32565 36731 32623 36737
rect 33962 36728 33968 36780
rect 34020 36768 34026 36780
rect 34589 36771 34647 36777
rect 34589 36768 34601 36771
rect 34020 36740 34601 36768
rect 34020 36728 34026 36740
rect 34589 36737 34601 36740
rect 34635 36737 34647 36771
rect 34589 36731 34647 36737
rect 36449 36771 36507 36777
rect 36449 36737 36461 36771
rect 36495 36768 36507 36771
rect 36722 36768 36728 36780
rect 36495 36740 36728 36768
rect 36495 36737 36507 36740
rect 36449 36731 36507 36737
rect 36722 36728 36728 36740
rect 36780 36728 36786 36780
rect 37829 36771 37887 36777
rect 37829 36737 37841 36771
rect 37875 36768 37887 36771
rect 37918 36768 37924 36780
rect 37875 36740 37924 36768
rect 37875 36737 37887 36740
rect 37829 36731 37887 36737
rect 37918 36728 37924 36740
rect 37976 36728 37982 36780
rect 31846 36700 31852 36712
rect 30944 36672 31852 36700
rect 26200 36660 26206 36672
rect 31846 36660 31852 36672
rect 31904 36660 31910 36712
rect 34238 36660 34244 36712
rect 34296 36700 34302 36712
rect 34333 36703 34391 36709
rect 34333 36700 34345 36703
rect 34296 36672 34345 36700
rect 34296 36660 34302 36672
rect 34333 36669 34345 36672
rect 34379 36669 34391 36703
rect 34333 36663 34391 36669
rect 36630 36660 36636 36712
rect 36688 36660 36694 36712
rect 38105 36703 38163 36709
rect 38105 36669 38117 36703
rect 38151 36700 38163 36703
rect 39022 36700 39028 36712
rect 38151 36672 39028 36700
rect 38151 36669 38163 36672
rect 38105 36663 38163 36669
rect 39022 36660 39028 36672
rect 39080 36660 39086 36712
rect 9122 36564 9128 36576
rect 8220 36536 9128 36564
rect 9122 36524 9128 36536
rect 9180 36524 9186 36576
rect 12069 36567 12127 36573
rect 12069 36533 12081 36567
rect 12115 36564 12127 36567
rect 12710 36564 12716 36576
rect 12115 36536 12716 36564
rect 12115 36533 12127 36536
rect 12069 36527 12127 36533
rect 12710 36524 12716 36536
rect 12768 36524 12774 36576
rect 16022 36524 16028 36576
rect 16080 36524 16086 36576
rect 16942 36524 16948 36576
rect 17000 36524 17006 36576
rect 19521 36567 19579 36573
rect 19521 36533 19533 36567
rect 19567 36564 19579 36567
rect 20162 36564 20168 36576
rect 19567 36536 20168 36564
rect 19567 36533 19579 36536
rect 19521 36527 19579 36533
rect 20162 36524 20168 36536
rect 20220 36564 20226 36576
rect 20530 36564 20536 36576
rect 20220 36536 20536 36564
rect 20220 36524 20226 36536
rect 20530 36524 20536 36536
rect 20588 36524 20594 36576
rect 23014 36524 23020 36576
rect 23072 36564 23078 36576
rect 23477 36567 23535 36573
rect 23477 36564 23489 36567
rect 23072 36536 23489 36564
rect 23072 36524 23078 36536
rect 23477 36533 23489 36536
rect 23523 36533 23535 36567
rect 23477 36527 23535 36533
rect 26329 36567 26387 36573
rect 26329 36533 26341 36567
rect 26375 36564 26387 36567
rect 26418 36564 26424 36576
rect 26375 36536 26424 36564
rect 26375 36533 26387 36536
rect 26329 36527 26387 36533
rect 26418 36524 26424 36536
rect 26476 36524 26482 36576
rect 28718 36524 28724 36576
rect 28776 36564 28782 36576
rect 28905 36567 28963 36573
rect 28905 36564 28917 36567
rect 28776 36536 28917 36564
rect 28776 36524 28782 36536
rect 28905 36533 28917 36536
rect 28951 36533 28963 36567
rect 28905 36527 28963 36533
rect 29641 36567 29699 36573
rect 29641 36533 29653 36567
rect 29687 36564 29699 36567
rect 30098 36564 30104 36576
rect 29687 36536 30104 36564
rect 29687 36533 29699 36536
rect 29641 36527 29699 36533
rect 30098 36524 30104 36536
rect 30156 36524 30162 36576
rect 33410 36524 33416 36576
rect 33468 36564 33474 36576
rect 33689 36567 33747 36573
rect 33689 36564 33701 36567
rect 33468 36536 33701 36564
rect 33468 36524 33474 36536
rect 33689 36533 33701 36536
rect 33735 36533 33747 36567
rect 33689 36527 33747 36533
rect 35710 36524 35716 36576
rect 35768 36524 35774 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 13170 36320 13176 36372
rect 13228 36360 13234 36372
rect 13449 36363 13507 36369
rect 13449 36360 13461 36363
rect 13228 36332 13461 36360
rect 13228 36320 13234 36332
rect 13449 36329 13461 36332
rect 13495 36329 13507 36363
rect 13449 36323 13507 36329
rect 15194 36320 15200 36372
rect 15252 36320 15258 36372
rect 15764 36332 18184 36360
rect 9214 36252 9220 36304
rect 9272 36252 9278 36304
rect 14182 36252 14188 36304
rect 14240 36292 14246 36304
rect 15764 36292 15792 36332
rect 14240 36264 15792 36292
rect 14240 36252 14246 36264
rect 5626 36184 5632 36236
rect 5684 36224 5690 36236
rect 5721 36227 5779 36233
rect 5721 36224 5733 36227
rect 5684 36196 5733 36224
rect 5684 36184 5690 36196
rect 5721 36193 5733 36196
rect 5767 36193 5779 36227
rect 5721 36187 5779 36193
rect 5902 36184 5908 36236
rect 5960 36184 5966 36236
rect 9585 36227 9643 36233
rect 9585 36193 9597 36227
rect 9631 36224 9643 36227
rect 9674 36224 9680 36236
rect 9631 36196 9680 36224
rect 9631 36193 9643 36196
rect 9585 36187 9643 36193
rect 9674 36184 9680 36196
rect 9732 36184 9738 36236
rect 12894 36184 12900 36236
rect 12952 36184 12958 36236
rect 15749 36227 15807 36233
rect 15749 36193 15761 36227
rect 15795 36224 15807 36227
rect 15930 36224 15936 36236
rect 15795 36196 15936 36224
rect 15795 36193 15807 36196
rect 15749 36187 15807 36193
rect 15930 36184 15936 36196
rect 15988 36184 15994 36236
rect 16022 36184 16028 36236
rect 16080 36224 16086 36236
rect 18156 36224 18184 36332
rect 22278 36320 22284 36372
rect 22336 36360 22342 36372
rect 24946 36360 24952 36372
rect 22336 36332 24952 36360
rect 22336 36320 22342 36332
rect 24946 36320 24952 36332
rect 25004 36320 25010 36372
rect 25590 36320 25596 36372
rect 25648 36320 25654 36372
rect 27154 36360 27160 36372
rect 25700 36332 27160 36360
rect 18966 36252 18972 36304
rect 19024 36292 19030 36304
rect 21266 36292 21272 36304
rect 19024 36264 21272 36292
rect 19024 36252 19030 36264
rect 21266 36252 21272 36264
rect 21324 36252 21330 36304
rect 25700 36292 25728 36332
rect 27154 36320 27160 36332
rect 27212 36360 27218 36372
rect 27525 36363 27583 36369
rect 27525 36360 27537 36363
rect 27212 36332 27537 36360
rect 27212 36320 27218 36332
rect 27525 36329 27537 36332
rect 27571 36329 27583 36363
rect 27525 36323 27583 36329
rect 28258 36320 28264 36372
rect 28316 36320 28322 36372
rect 30098 36320 30104 36372
rect 30156 36320 30162 36372
rect 31849 36363 31907 36369
rect 31849 36329 31861 36363
rect 31895 36360 31907 36363
rect 32398 36360 32404 36372
rect 31895 36332 32404 36360
rect 31895 36329 31907 36332
rect 31849 36323 31907 36329
rect 32398 36320 32404 36332
rect 32456 36320 32462 36372
rect 33962 36320 33968 36372
rect 34020 36320 34026 36372
rect 36814 36360 36820 36372
rect 34072 36332 36820 36360
rect 34072 36292 34100 36332
rect 36814 36320 36820 36332
rect 36872 36320 36878 36372
rect 22480 36264 25728 36292
rect 28552 36264 34100 36292
rect 22480 36236 22508 36264
rect 21453 36227 21511 36233
rect 21453 36224 21465 36227
rect 16080 36196 18092 36224
rect 18156 36196 21465 36224
rect 16080 36184 16086 36196
rect 4614 36116 4620 36168
rect 4672 36156 4678 36168
rect 6457 36159 6515 36165
rect 6457 36156 6469 36159
rect 4672 36128 6469 36156
rect 4672 36116 4678 36128
rect 6457 36125 6469 36128
rect 6503 36156 6515 36159
rect 9122 36156 9128 36168
rect 6503 36128 9128 36156
rect 6503 36125 6515 36128
rect 6457 36119 6515 36125
rect 9122 36116 9128 36128
rect 9180 36156 9186 36168
rect 10505 36159 10563 36165
rect 10505 36156 10517 36159
rect 9180 36128 10517 36156
rect 9180 36116 9186 36128
rect 10505 36125 10517 36128
rect 10551 36125 10563 36159
rect 10505 36119 10563 36125
rect 12710 36116 12716 36168
rect 12768 36156 12774 36168
rect 12989 36159 13047 36165
rect 12989 36156 13001 36159
rect 12768 36128 13001 36156
rect 12768 36116 12774 36128
rect 12989 36125 13001 36128
rect 13035 36156 13047 36159
rect 13262 36156 13268 36168
rect 13035 36128 13268 36156
rect 13035 36125 13047 36128
rect 12989 36119 13047 36125
rect 13262 36116 13268 36128
rect 13320 36116 13326 36168
rect 15102 36116 15108 36168
rect 15160 36116 15166 36168
rect 16114 36116 16120 36168
rect 16172 36116 16178 36168
rect 18064 36165 18092 36196
rect 21453 36193 21465 36196
rect 21499 36193 21511 36227
rect 22278 36224 22284 36236
rect 21453 36187 21511 36193
rect 22066 36196 22284 36224
rect 18049 36159 18107 36165
rect 18049 36125 18061 36159
rect 18095 36125 18107 36159
rect 19889 36159 19947 36165
rect 18049 36119 18107 36125
rect 18156 36128 19748 36156
rect 5534 36048 5540 36100
rect 5592 36088 5598 36100
rect 5629 36091 5687 36097
rect 5629 36088 5641 36091
rect 5592 36060 5641 36088
rect 5592 36048 5598 36060
rect 5629 36057 5641 36060
rect 5675 36057 5687 36091
rect 5629 36051 5687 36057
rect 6724 36091 6782 36097
rect 6724 36057 6736 36091
rect 6770 36088 6782 36091
rect 7098 36088 7104 36100
rect 6770 36060 7104 36088
rect 6770 36057 6782 36060
rect 6724 36051 6782 36057
rect 7098 36048 7104 36060
rect 7156 36048 7162 36100
rect 9582 36048 9588 36100
rect 9640 36088 9646 36100
rect 9677 36091 9735 36097
rect 9677 36088 9689 36091
rect 9640 36060 9689 36088
rect 9640 36048 9646 36060
rect 9677 36057 9689 36060
rect 9723 36057 9735 36091
rect 9677 36051 9735 36057
rect 9769 36091 9827 36097
rect 9769 36057 9781 36091
rect 9815 36088 9827 36091
rect 10134 36088 10140 36100
rect 9815 36060 10140 36088
rect 9815 36057 9827 36060
rect 9769 36051 9827 36057
rect 10134 36048 10140 36060
rect 10192 36048 10198 36100
rect 10772 36091 10830 36097
rect 10772 36057 10784 36091
rect 10818 36088 10830 36091
rect 11698 36088 11704 36100
rect 10818 36060 11704 36088
rect 10818 36057 10830 36060
rect 10772 36051 10830 36057
rect 11698 36048 11704 36060
rect 11756 36048 11762 36100
rect 16942 36048 16948 36100
rect 17000 36048 17006 36100
rect 18156 36088 18184 36128
rect 17236 36060 18184 36088
rect 18325 36091 18383 36097
rect 5258 35980 5264 36032
rect 5316 35980 5322 36032
rect 7834 35980 7840 36032
rect 7892 35980 7898 36032
rect 11882 35980 11888 36032
rect 11940 35980 11946 36032
rect 13081 36023 13139 36029
rect 13081 35989 13093 36023
rect 13127 36020 13139 36023
rect 13446 36020 13452 36032
rect 13127 35992 13452 36020
rect 13127 35989 13139 35992
rect 13081 35983 13139 35989
rect 13446 35980 13452 35992
rect 13504 36020 13510 36032
rect 17236 36020 17264 36060
rect 18325 36057 18337 36091
rect 18371 36088 18383 36091
rect 18690 36088 18696 36100
rect 18371 36060 18696 36088
rect 18371 36057 18383 36060
rect 18325 36051 18383 36057
rect 18690 36048 18696 36060
rect 18748 36048 18754 36100
rect 18966 36048 18972 36100
rect 19024 36088 19030 36100
rect 19613 36091 19671 36097
rect 19613 36088 19625 36091
rect 19024 36060 19625 36088
rect 19024 36048 19030 36060
rect 19613 36057 19625 36060
rect 19659 36057 19671 36091
rect 19720 36088 19748 36128
rect 19889 36125 19901 36159
rect 19935 36156 19947 36159
rect 20254 36156 20260 36168
rect 19935 36128 20260 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 20254 36116 20260 36128
rect 20312 36116 20318 36168
rect 20346 36116 20352 36168
rect 20404 36156 20410 36168
rect 20441 36159 20499 36165
rect 20441 36156 20453 36159
rect 20404 36128 20453 36156
rect 20404 36116 20410 36128
rect 20441 36125 20453 36128
rect 20487 36125 20499 36159
rect 20441 36119 20499 36125
rect 20714 36116 20720 36168
rect 20772 36116 20778 36168
rect 22066 36088 22094 36196
rect 22278 36184 22284 36196
rect 22336 36184 22342 36236
rect 22462 36184 22468 36236
rect 22520 36184 22526 36236
rect 26142 36184 26148 36236
rect 26200 36184 26206 36236
rect 26326 36184 26332 36236
rect 26384 36184 26390 36236
rect 26418 36184 26424 36236
rect 26476 36184 26482 36236
rect 23014 36156 23020 36168
rect 22954 36128 23020 36156
rect 23014 36116 23020 36128
rect 23072 36116 23078 36168
rect 23382 36116 23388 36168
rect 23440 36156 23446 36168
rect 24578 36156 24584 36168
rect 23440 36128 24584 36156
rect 23440 36116 23446 36128
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25685 36159 25743 36165
rect 25685 36156 25697 36159
rect 24688 36128 25697 36156
rect 19720 36060 22094 36088
rect 19613 36051 19671 36057
rect 23658 36048 23664 36100
rect 23716 36088 23722 36100
rect 24688 36088 24716 36128
rect 25685 36125 25697 36128
rect 25731 36156 25743 36159
rect 26344 36156 26372 36184
rect 28445 36159 28503 36165
rect 28445 36156 28457 36159
rect 25731 36128 28457 36156
rect 25731 36125 25743 36128
rect 25685 36119 25743 36125
rect 28445 36125 28457 36128
rect 28491 36156 28503 36159
rect 28552 36156 28580 36264
rect 31478 36184 31484 36236
rect 31536 36184 31542 36236
rect 33042 36224 33048 36236
rect 31726 36196 33048 36224
rect 28491 36128 28580 36156
rect 28721 36159 28779 36165
rect 28491 36125 28503 36128
rect 28445 36119 28503 36125
rect 28721 36125 28733 36159
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 23716 36060 24716 36088
rect 23716 36048 23722 36060
rect 24854 36048 24860 36100
rect 24912 36048 24918 36100
rect 27706 36048 27712 36100
rect 27764 36088 27770 36100
rect 28736 36088 28764 36119
rect 30190 36116 30196 36168
rect 30248 36116 30254 36168
rect 30469 36159 30527 36165
rect 30469 36125 30481 36159
rect 30515 36125 30527 36159
rect 30469 36119 30527 36125
rect 31573 36159 31631 36165
rect 31573 36125 31585 36159
rect 31619 36156 31631 36159
rect 31726 36156 31754 36196
rect 33042 36184 33048 36196
rect 33100 36224 33106 36236
rect 33597 36227 33655 36233
rect 33597 36224 33609 36227
rect 33100 36196 33609 36224
rect 33100 36184 33106 36196
rect 33597 36193 33609 36196
rect 33643 36193 33655 36227
rect 33597 36187 33655 36193
rect 34238 36184 34244 36236
rect 34296 36224 34302 36236
rect 34885 36227 34943 36233
rect 34885 36224 34897 36227
rect 34296 36196 34897 36224
rect 34296 36184 34302 36196
rect 34885 36193 34897 36196
rect 34931 36193 34943 36227
rect 34885 36187 34943 36193
rect 31619 36128 31754 36156
rect 31619 36125 31631 36128
rect 31573 36119 31631 36125
rect 27764 36060 28764 36088
rect 30484 36088 30512 36119
rect 32674 36116 32680 36168
rect 32732 36156 32738 36168
rect 32953 36159 33011 36165
rect 32953 36156 32965 36159
rect 32732 36128 32965 36156
rect 32732 36116 32738 36128
rect 32953 36125 32965 36128
rect 32999 36125 33011 36159
rect 32953 36119 33011 36125
rect 33781 36159 33839 36165
rect 33781 36125 33793 36159
rect 33827 36125 33839 36159
rect 34900 36156 34928 36187
rect 36354 36156 36360 36168
rect 34900 36128 36360 36156
rect 33781 36119 33839 36125
rect 31846 36088 31852 36100
rect 30484 36060 31852 36088
rect 27764 36048 27770 36060
rect 31846 36048 31852 36060
rect 31904 36048 31910 36100
rect 32490 36048 32496 36100
rect 32548 36088 32554 36100
rect 32769 36091 32827 36097
rect 32769 36088 32781 36091
rect 32548 36060 32781 36088
rect 32548 36048 32554 36060
rect 32769 36057 32781 36060
rect 32815 36057 32827 36091
rect 32769 36051 32827 36057
rect 33137 36091 33195 36097
rect 33137 36057 33149 36091
rect 33183 36088 33195 36091
rect 33796 36088 33824 36119
rect 36354 36116 36360 36128
rect 36412 36156 36418 36168
rect 36817 36159 36875 36165
rect 36817 36156 36829 36159
rect 36412 36128 36829 36156
rect 36412 36116 36418 36128
rect 36817 36125 36829 36128
rect 36863 36125 36875 36159
rect 36817 36119 36875 36125
rect 33183 36060 33824 36088
rect 33183 36057 33195 36060
rect 33137 36051 33195 36057
rect 34514 36048 34520 36100
rect 34572 36088 34578 36100
rect 35130 36091 35188 36097
rect 35130 36088 35142 36091
rect 34572 36060 35142 36088
rect 34572 36048 34578 36060
rect 35130 36057 35142 36060
rect 35176 36057 35188 36091
rect 35130 36051 35188 36057
rect 37084 36091 37142 36097
rect 37084 36057 37096 36091
rect 37130 36088 37142 36091
rect 37458 36088 37464 36100
rect 37130 36060 37464 36088
rect 37130 36057 37142 36060
rect 37084 36051 37142 36057
rect 37458 36048 37464 36060
rect 37516 36048 37522 36100
rect 13504 35992 17264 36020
rect 17543 36023 17601 36029
rect 13504 35980 13510 35992
rect 17543 35989 17555 36023
rect 17589 36020 17601 36023
rect 19426 36020 19432 36032
rect 17589 35992 19432 36020
rect 17589 35989 17601 35992
rect 17543 35983 17601 35989
rect 19426 35980 19432 35992
rect 19484 35980 19490 36032
rect 20438 35980 20444 36032
rect 20496 35980 20502 36032
rect 22465 36023 22523 36029
rect 22465 35989 22477 36023
rect 22511 36020 22523 36023
rect 22922 36020 22928 36032
rect 22511 35992 22928 36020
rect 22511 35989 22523 35992
rect 22465 35983 22523 35989
rect 22922 35980 22928 35992
rect 22980 35980 22986 36032
rect 28629 36023 28687 36029
rect 28629 35989 28641 36023
rect 28675 36020 28687 36023
rect 28718 36020 28724 36032
rect 28675 35992 28724 36020
rect 28675 35989 28687 35992
rect 28629 35983 28687 35989
rect 28718 35980 28724 35992
rect 28776 35980 28782 36032
rect 29178 35980 29184 36032
rect 29236 36020 29242 36032
rect 29917 36023 29975 36029
rect 29917 36020 29929 36023
rect 29236 35992 29929 36020
rect 29236 35980 29242 35992
rect 29917 35989 29929 35992
rect 29963 35989 29975 36023
rect 29917 35983 29975 35989
rect 36078 35980 36084 36032
rect 36136 36020 36142 36032
rect 36265 36023 36323 36029
rect 36265 36020 36277 36023
rect 36136 35992 36277 36020
rect 36136 35980 36142 35992
rect 36265 35989 36277 35992
rect 36311 35989 36323 36023
rect 36265 35983 36323 35989
rect 37826 35980 37832 36032
rect 37884 36020 37890 36032
rect 38197 36023 38255 36029
rect 38197 36020 38209 36023
rect 37884 35992 38209 36020
rect 37884 35980 37890 35992
rect 38197 35989 38209 35992
rect 38243 35989 38255 36023
rect 38197 35983 38255 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 7098 35776 7104 35828
rect 7156 35776 7162 35828
rect 7558 35776 7564 35828
rect 7616 35816 7622 35828
rect 7834 35816 7840 35828
rect 7616 35788 7840 35816
rect 7616 35776 7622 35788
rect 7834 35776 7840 35788
rect 7892 35776 7898 35828
rect 11698 35776 11704 35828
rect 11756 35776 11762 35828
rect 18414 35776 18420 35828
rect 18472 35816 18478 35828
rect 20714 35816 20720 35828
rect 18472 35788 20720 35816
rect 18472 35776 18478 35788
rect 20714 35776 20720 35788
rect 20772 35816 20778 35828
rect 21358 35816 21364 35828
rect 20772 35788 21364 35816
rect 20772 35776 20778 35788
rect 21358 35776 21364 35788
rect 21416 35776 21422 35828
rect 22097 35819 22155 35825
rect 22097 35785 22109 35819
rect 22143 35816 22155 35819
rect 22370 35816 22376 35828
rect 22143 35788 22376 35816
rect 22143 35785 22155 35788
rect 22097 35779 22155 35785
rect 22370 35776 22376 35788
rect 22428 35776 22434 35828
rect 22557 35819 22615 35825
rect 22557 35785 22569 35819
rect 22603 35816 22615 35819
rect 23014 35816 23020 35828
rect 22603 35788 23020 35816
rect 22603 35785 22615 35788
rect 22557 35779 22615 35785
rect 23014 35776 23020 35788
rect 23072 35776 23078 35828
rect 32677 35819 32735 35825
rect 32677 35785 32689 35819
rect 32723 35816 32735 35819
rect 33042 35816 33048 35828
rect 32723 35788 33048 35816
rect 32723 35785 32735 35788
rect 32677 35779 32735 35785
rect 33042 35776 33048 35788
rect 33100 35776 33106 35828
rect 33413 35819 33471 35825
rect 33413 35785 33425 35819
rect 33459 35816 33471 35819
rect 34514 35816 34520 35828
rect 33459 35788 34520 35816
rect 33459 35785 33471 35788
rect 33413 35779 33471 35785
rect 34514 35776 34520 35788
rect 34572 35776 34578 35828
rect 36817 35819 36875 35825
rect 36817 35785 36829 35819
rect 36863 35816 36875 35819
rect 36906 35816 36912 35828
rect 36863 35788 36912 35816
rect 36863 35785 36875 35788
rect 36817 35779 36875 35785
rect 36906 35776 36912 35788
rect 36964 35776 36970 35828
rect 37458 35776 37464 35828
rect 37516 35776 37522 35828
rect 9306 35748 9312 35760
rect 7760 35720 9312 35748
rect 7466 35640 7472 35692
rect 7524 35640 7530 35692
rect 5810 35572 5816 35624
rect 5868 35612 5874 35624
rect 7760 35621 7788 35720
rect 9306 35708 9312 35720
rect 9364 35748 9370 35760
rect 12894 35748 12900 35760
rect 9364 35720 12900 35748
rect 9364 35708 9370 35720
rect 9858 35640 9864 35692
rect 9916 35640 9922 35692
rect 7745 35615 7803 35621
rect 7745 35612 7757 35615
rect 5868 35584 7757 35612
rect 5868 35572 5874 35584
rect 7745 35581 7757 35584
rect 7791 35581 7803 35615
rect 7745 35575 7803 35581
rect 9950 35572 9956 35624
rect 10008 35572 10014 35624
rect 10152 35621 10180 35720
rect 12066 35640 12072 35692
rect 12124 35640 12130 35692
rect 10137 35615 10195 35621
rect 10137 35581 10149 35615
rect 10183 35581 10195 35615
rect 10137 35575 10195 35581
rect 11790 35572 11796 35624
rect 11848 35612 11854 35624
rect 12360 35621 12388 35720
rect 12894 35708 12900 35720
rect 12952 35748 12958 35760
rect 12952 35720 20668 35748
rect 12952 35708 12958 35720
rect 14921 35683 14979 35689
rect 14921 35649 14933 35683
rect 14967 35680 14979 35683
rect 15102 35680 15108 35692
rect 14967 35652 15108 35680
rect 14967 35649 14979 35652
rect 14921 35643 14979 35649
rect 15102 35640 15108 35652
rect 15160 35640 15166 35692
rect 17034 35640 17040 35692
rect 17092 35640 17098 35692
rect 18233 35683 18291 35689
rect 18233 35649 18245 35683
rect 18279 35680 18291 35683
rect 18414 35680 18420 35692
rect 18279 35652 18420 35680
rect 18279 35649 18291 35652
rect 18233 35643 18291 35649
rect 18414 35640 18420 35652
rect 18472 35640 18478 35692
rect 18598 35640 18604 35692
rect 18656 35640 18662 35692
rect 18966 35640 18972 35692
rect 19024 35640 19030 35692
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35680 19671 35683
rect 20346 35680 20352 35692
rect 19659 35652 20352 35680
rect 19659 35649 19671 35652
rect 19613 35643 19671 35649
rect 12161 35615 12219 35621
rect 12161 35612 12173 35615
rect 11848 35584 12173 35612
rect 11848 35572 11854 35584
rect 12161 35581 12173 35584
rect 12207 35581 12219 35615
rect 12161 35575 12219 35581
rect 12345 35615 12403 35621
rect 12345 35581 12357 35615
rect 12391 35581 12403 35615
rect 12345 35575 12403 35581
rect 18690 35572 18696 35624
rect 18748 35612 18754 35624
rect 19628 35612 19656 35643
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20530 35640 20536 35692
rect 20588 35640 20594 35692
rect 20640 35680 20668 35720
rect 21266 35708 21272 35760
rect 21324 35748 21330 35760
rect 23382 35748 23388 35760
rect 21324 35720 23388 35748
rect 21324 35708 21330 35720
rect 23382 35708 23388 35720
rect 23440 35708 23446 35760
rect 23566 35708 23572 35760
rect 23624 35748 23630 35760
rect 23624 35720 26096 35748
rect 23624 35708 23630 35720
rect 22465 35683 22523 35689
rect 20640 35652 22094 35680
rect 18748 35584 19656 35612
rect 18748 35572 18754 35584
rect 20806 35572 20812 35624
rect 20864 35572 20870 35624
rect 9858 35504 9864 35556
rect 9916 35544 9922 35556
rect 16206 35544 16212 35556
rect 9916 35516 16212 35544
rect 9916 35504 9922 35516
rect 16206 35504 16212 35516
rect 16264 35504 16270 35556
rect 22066 35544 22094 35652
rect 22465 35649 22477 35683
rect 22511 35680 22523 35683
rect 22922 35680 22928 35692
rect 22511 35652 22928 35680
rect 22511 35649 22523 35652
rect 22465 35643 22523 35649
rect 22922 35640 22928 35652
rect 22980 35640 22986 35692
rect 23658 35640 23664 35692
rect 23716 35640 23722 35692
rect 23750 35640 23756 35692
rect 23808 35680 23814 35692
rect 23845 35683 23903 35689
rect 23845 35680 23857 35683
rect 23808 35652 23857 35680
rect 23808 35640 23814 35652
rect 23845 35649 23857 35652
rect 23891 35649 23903 35683
rect 23845 35643 23903 35649
rect 25222 35640 25228 35692
rect 25280 35680 25286 35692
rect 26068 35689 26096 35720
rect 25409 35683 25467 35689
rect 25409 35680 25421 35683
rect 25280 35652 25421 35680
rect 25280 35640 25286 35652
rect 25409 35649 25421 35652
rect 25455 35680 25467 35683
rect 26053 35683 26111 35689
rect 25455 35652 25636 35680
rect 25455 35649 25467 35652
rect 25409 35643 25467 35649
rect 22741 35615 22799 35621
rect 22741 35581 22753 35615
rect 22787 35612 22799 35615
rect 23293 35615 23351 35621
rect 23293 35612 23305 35615
rect 22787 35584 23305 35612
rect 22787 35581 22799 35584
rect 22741 35575 22799 35581
rect 23293 35581 23305 35584
rect 23339 35581 23351 35615
rect 23293 35575 23351 35581
rect 24949 35615 25007 35621
rect 24949 35581 24961 35615
rect 24995 35612 25007 35615
rect 25130 35612 25136 35624
rect 24995 35584 25136 35612
rect 24995 35581 25007 35584
rect 24949 35575 25007 35581
rect 22756 35544 22784 35575
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 25498 35572 25504 35624
rect 25556 35572 25562 35624
rect 25608 35612 25636 35652
rect 26053 35649 26065 35683
rect 26099 35649 26111 35683
rect 26053 35643 26111 35649
rect 27246 35640 27252 35692
rect 27304 35640 27310 35692
rect 28810 35640 28816 35692
rect 28868 35640 28874 35692
rect 29086 35689 29092 35692
rect 29080 35643 29092 35689
rect 29086 35640 29092 35643
rect 29144 35640 29150 35692
rect 32490 35640 32496 35692
rect 32548 35640 32554 35692
rect 32674 35640 32680 35692
rect 32732 35680 32738 35692
rect 33321 35683 33379 35689
rect 33321 35680 33333 35683
rect 32732 35652 33333 35680
rect 32732 35640 32738 35652
rect 33321 35649 33333 35652
rect 33367 35649 33379 35683
rect 33321 35643 33379 35649
rect 33502 35640 33508 35692
rect 33560 35640 33566 35692
rect 36722 35640 36728 35692
rect 36780 35640 36786 35692
rect 37642 35640 37648 35692
rect 37700 35680 37706 35692
rect 37826 35680 37832 35692
rect 37700 35652 37832 35680
rect 37700 35640 37706 35652
rect 37826 35640 37832 35652
rect 37884 35640 37890 35692
rect 26237 35615 26295 35621
rect 26237 35612 26249 35615
rect 25608 35584 26249 35612
rect 26237 35581 26249 35584
rect 26283 35581 26295 35615
rect 26237 35575 26295 35581
rect 27706 35572 27712 35624
rect 27764 35572 27770 35624
rect 37918 35572 37924 35624
rect 37976 35572 37982 35624
rect 38010 35572 38016 35624
rect 38068 35572 38074 35624
rect 22066 35516 22784 35544
rect 24857 35547 24915 35553
rect 24857 35513 24869 35547
rect 24903 35544 24915 35547
rect 26050 35544 26056 35556
rect 24903 35516 26056 35544
rect 24903 35513 24915 35516
rect 24857 35507 24915 35513
rect 26050 35504 26056 35516
rect 26108 35504 26114 35556
rect 9398 35436 9404 35488
rect 9456 35476 9462 35488
rect 9493 35479 9551 35485
rect 9493 35476 9505 35479
rect 9456 35448 9505 35476
rect 9456 35436 9462 35448
rect 9493 35445 9505 35448
rect 9539 35445 9551 35479
rect 9493 35439 9551 35445
rect 14734 35436 14740 35488
rect 14792 35476 14798 35488
rect 14829 35479 14887 35485
rect 14829 35476 14841 35479
rect 14792 35448 14841 35476
rect 14792 35436 14798 35448
rect 14829 35445 14841 35448
rect 14875 35445 14887 35479
rect 14829 35439 14887 35445
rect 16942 35436 16948 35488
rect 17000 35436 17006 35488
rect 18230 35436 18236 35488
rect 18288 35436 18294 35488
rect 23382 35436 23388 35488
rect 23440 35476 23446 35488
rect 25038 35476 25044 35488
rect 23440 35448 25044 35476
rect 23440 35436 23446 35448
rect 25038 35436 25044 35448
rect 25096 35436 25102 35488
rect 30190 35436 30196 35488
rect 30248 35436 30254 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 25222 35272 25228 35284
rect 16960 35244 23336 35272
rect 10594 35164 10600 35216
rect 10652 35204 10658 35216
rect 11333 35207 11391 35213
rect 11333 35204 11345 35207
rect 10652 35176 11345 35204
rect 10652 35164 10658 35176
rect 11333 35173 11345 35176
rect 11379 35173 11391 35207
rect 11333 35167 11391 35173
rect 5810 35096 5816 35148
rect 5868 35096 5874 35148
rect 11793 35139 11851 35145
rect 11793 35105 11805 35139
rect 11839 35136 11851 35139
rect 12066 35136 12072 35148
rect 11839 35108 12072 35136
rect 11839 35105 11851 35108
rect 11793 35099 11851 35105
rect 12066 35096 12072 35108
rect 12124 35096 12130 35148
rect 13357 35139 13415 35145
rect 13357 35105 13369 35139
rect 13403 35136 13415 35139
rect 13446 35136 13452 35148
rect 13403 35108 13452 35136
rect 13403 35105 13415 35108
rect 13357 35099 13415 35105
rect 13446 35096 13452 35108
rect 13504 35096 13510 35148
rect 15565 35139 15623 35145
rect 15565 35105 15577 35139
rect 15611 35136 15623 35139
rect 15930 35136 15936 35148
rect 15611 35108 15936 35136
rect 15611 35105 15623 35108
rect 15565 35099 15623 35105
rect 15930 35096 15936 35108
rect 15988 35096 15994 35148
rect 16206 35096 16212 35148
rect 16264 35136 16270 35148
rect 16960 35136 16988 35244
rect 22462 35204 22468 35216
rect 16264 35108 16988 35136
rect 17144 35176 22468 35204
rect 16264 35096 16270 35108
rect 9122 35028 9128 35080
rect 9180 35028 9186 35080
rect 9398 35077 9404 35080
rect 9392 35068 9404 35077
rect 9359 35040 9404 35068
rect 9392 35031 9404 35040
rect 9398 35028 9404 35031
rect 9456 35028 9462 35080
rect 10134 35028 10140 35080
rect 10192 35068 10198 35080
rect 11885 35071 11943 35077
rect 11885 35068 11897 35071
rect 10192 35040 11897 35068
rect 10192 35028 10198 35040
rect 11885 35037 11897 35040
rect 11931 35068 11943 35071
rect 13081 35071 13139 35077
rect 13081 35068 13093 35071
rect 11931 35040 13093 35068
rect 11931 35037 11943 35040
rect 11885 35031 11943 35037
rect 13081 35037 13093 35040
rect 13127 35037 13139 35071
rect 13081 35031 13139 35037
rect 5537 35003 5595 35009
rect 5537 34969 5549 35003
rect 5583 35000 5595 35003
rect 6362 35000 6368 35012
rect 5583 34972 6368 35000
rect 5583 34969 5595 34972
rect 5537 34963 5595 34969
rect 6362 34960 6368 34972
rect 6420 35000 6426 35012
rect 7006 35000 7012 35012
rect 6420 34972 7012 35000
rect 6420 34960 6426 34972
rect 7006 34960 7012 34972
rect 7064 34960 7070 35012
rect 11790 34960 11796 35012
rect 11848 34960 11854 35012
rect 12618 34960 12624 35012
rect 12676 34960 12682 35012
rect 5166 34892 5172 34944
rect 5224 34892 5230 34944
rect 5626 34892 5632 34944
rect 5684 34892 5690 34944
rect 9950 34892 9956 34944
rect 10008 34932 10014 34944
rect 10505 34935 10563 34941
rect 10505 34932 10517 34935
rect 10008 34904 10517 34932
rect 10008 34892 10014 34904
rect 10505 34901 10517 34904
rect 10551 34901 10563 34935
rect 13096 34932 13124 35031
rect 13262 35028 13268 35080
rect 13320 35028 13326 35080
rect 16942 35028 16948 35080
rect 17000 35028 17006 35080
rect 15838 34960 15844 35012
rect 15896 34960 15902 35012
rect 17144 34932 17172 35176
rect 22462 35164 22468 35176
rect 22520 35164 22526 35216
rect 17313 35139 17371 35145
rect 17313 35105 17325 35139
rect 17359 35136 17371 35139
rect 20254 35136 20260 35148
rect 17359 35108 20260 35136
rect 17359 35105 17371 35108
rect 17313 35099 17371 35105
rect 20254 35096 20260 35108
rect 20312 35096 20318 35148
rect 21082 35136 21088 35148
rect 20364 35108 21088 35136
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 18233 35071 18291 35077
rect 18233 35068 18245 35071
rect 18012 35040 18245 35068
rect 18012 35028 18018 35040
rect 18233 35037 18245 35040
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 18322 35028 18328 35080
rect 18380 35068 18386 35080
rect 18509 35071 18567 35077
rect 18509 35068 18521 35071
rect 18380 35040 18521 35068
rect 18380 35028 18386 35040
rect 18509 35037 18521 35040
rect 18555 35068 18567 35071
rect 18598 35068 18604 35080
rect 18555 35040 18604 35068
rect 18555 35037 18567 35040
rect 18509 35031 18567 35037
rect 18598 35028 18604 35040
rect 18656 35068 18662 35080
rect 18656 35040 19380 35068
rect 18656 35028 18662 35040
rect 18690 34960 18696 35012
rect 18748 35009 18754 35012
rect 18748 35003 18776 35009
rect 18764 34969 18776 35003
rect 19352 35000 19380 35040
rect 19426 35028 19432 35080
rect 19484 35028 19490 35080
rect 19705 35071 19763 35077
rect 19705 35037 19717 35071
rect 19751 35068 19763 35071
rect 20364 35068 20392 35108
rect 21082 35096 21088 35108
rect 21140 35096 21146 35148
rect 19751 35040 20392 35068
rect 19751 35037 19763 35040
rect 19705 35031 19763 35037
rect 19720 35000 19748 35031
rect 20438 35028 20444 35080
rect 20496 35028 20502 35080
rect 20622 35028 20628 35080
rect 20680 35028 20686 35080
rect 21100 35068 21128 35096
rect 22094 35068 22100 35080
rect 21100 35040 22100 35068
rect 22094 35028 22100 35040
rect 22152 35028 22158 35080
rect 23308 35068 23336 35244
rect 23400 35244 25228 35272
rect 23400 35145 23428 35244
rect 25222 35232 25228 35244
rect 25280 35232 25286 35284
rect 25958 35232 25964 35284
rect 26016 35272 26022 35284
rect 26016 35244 29040 35272
rect 26016 35232 26022 35244
rect 23474 35164 23480 35216
rect 23532 35164 23538 35216
rect 24854 35164 24860 35216
rect 24912 35204 24918 35216
rect 25317 35207 25375 35213
rect 25317 35204 25329 35207
rect 24912 35176 25329 35204
rect 24912 35164 24918 35176
rect 25317 35173 25329 35176
rect 25363 35204 25375 35207
rect 25498 35204 25504 35216
rect 25363 35176 25504 35204
rect 25363 35173 25375 35176
rect 25317 35167 25375 35173
rect 25498 35164 25504 35176
rect 25556 35164 25562 35216
rect 26881 35207 26939 35213
rect 26881 35173 26893 35207
rect 26927 35204 26939 35207
rect 27338 35204 27344 35216
rect 26927 35176 27344 35204
rect 26927 35173 26939 35176
rect 26881 35167 26939 35173
rect 27338 35164 27344 35176
rect 27396 35164 27402 35216
rect 29012 35204 29040 35244
rect 29086 35232 29092 35284
rect 29144 35232 29150 35284
rect 31481 35275 31539 35281
rect 31481 35241 31493 35275
rect 31527 35272 31539 35275
rect 32490 35272 32496 35284
rect 31527 35244 32496 35272
rect 31527 35241 31539 35244
rect 31481 35235 31539 35241
rect 32490 35232 32496 35244
rect 32548 35232 32554 35284
rect 32677 35275 32735 35281
rect 32677 35241 32689 35275
rect 32723 35272 32735 35275
rect 33502 35272 33508 35284
rect 32723 35244 33508 35272
rect 32723 35241 32735 35244
rect 32677 35235 32735 35241
rect 33502 35232 33508 35244
rect 33560 35232 33566 35284
rect 31202 35204 31208 35216
rect 29012 35176 31208 35204
rect 31202 35164 31208 35176
rect 31260 35164 31266 35216
rect 23385 35139 23443 35145
rect 23385 35105 23397 35139
rect 23431 35105 23443 35139
rect 23385 35099 23443 35105
rect 23860 35108 24992 35136
rect 23860 35080 23888 35108
rect 23658 35068 23664 35080
rect 23308 35040 23664 35068
rect 23658 35028 23664 35040
rect 23716 35028 23722 35080
rect 23842 35028 23848 35080
rect 23900 35028 23906 35080
rect 24964 35077 24992 35108
rect 25222 35096 25228 35148
rect 25280 35136 25286 35148
rect 25409 35139 25467 35145
rect 25409 35136 25421 35139
rect 25280 35108 25421 35136
rect 25280 35096 25286 35108
rect 25409 35105 25421 35108
rect 25455 35105 25467 35139
rect 25409 35099 25467 35105
rect 26142 35096 26148 35148
rect 26200 35136 26206 35148
rect 26200 35108 27476 35136
rect 26200 35096 26206 35108
rect 23937 35071 23995 35077
rect 23937 35037 23949 35071
rect 23983 35037 23995 35071
rect 23937 35031 23995 35037
rect 24857 35071 24915 35077
rect 24857 35037 24869 35071
rect 24903 35037 24915 35071
rect 24857 35031 24915 35037
rect 24949 35071 25007 35077
rect 24949 35037 24961 35071
rect 24995 35068 25007 35071
rect 25130 35068 25136 35080
rect 24995 35040 25136 35068
rect 24995 35037 25007 35040
rect 24949 35031 25007 35037
rect 19352 34972 19748 35000
rect 18748 34963 18776 34969
rect 18748 34960 18754 34963
rect 20530 34960 20536 35012
rect 20588 34960 20594 35012
rect 21085 35003 21143 35009
rect 21085 34969 21097 35003
rect 21131 35000 21143 35003
rect 21174 35000 21180 35012
rect 21131 34972 21180 35000
rect 21131 34969 21143 34972
rect 21085 34963 21143 34969
rect 21174 34960 21180 34972
rect 21232 34960 21238 35012
rect 22373 35003 22431 35009
rect 22373 34969 22385 35003
rect 22419 34969 22431 35003
rect 22373 34963 22431 34969
rect 13096 34904 17172 34932
rect 10505 34895 10563 34901
rect 18414 34892 18420 34944
rect 18472 34932 18478 34944
rect 18601 34935 18659 34941
rect 18601 34932 18613 34935
rect 18472 34904 18613 34932
rect 18472 34892 18478 34904
rect 18601 34901 18613 34904
rect 18647 34901 18659 34935
rect 18601 34895 18659 34901
rect 18877 34935 18935 34941
rect 18877 34901 18889 34935
rect 18923 34932 18935 34935
rect 20346 34932 20352 34944
rect 18923 34904 20352 34932
rect 18923 34901 18935 34904
rect 18877 34895 18935 34901
rect 20346 34892 20352 34904
rect 20404 34892 20410 34944
rect 22388 34932 22416 34963
rect 23014 34960 23020 35012
rect 23072 34960 23078 35012
rect 23382 34932 23388 34944
rect 22388 34904 23388 34932
rect 23382 34892 23388 34904
rect 23440 34892 23446 34944
rect 23952 34932 23980 35031
rect 24872 35000 24900 35031
rect 25130 35028 25136 35040
rect 25188 35028 25194 35080
rect 26602 35028 26608 35080
rect 26660 35028 26666 35080
rect 27448 35077 27476 35108
rect 29178 35096 29184 35148
rect 29236 35096 29242 35148
rect 35710 35136 35716 35148
rect 31220 35108 35716 35136
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 26896 35040 27353 35068
rect 26896 35012 26924 35040
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 27341 35031 27399 35037
rect 27434 35071 27492 35077
rect 27434 35037 27446 35071
rect 27480 35037 27492 35071
rect 27434 35031 27492 35037
rect 28902 35028 28908 35080
rect 28960 35028 28966 35080
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35068 29055 35071
rect 29270 35068 29276 35080
rect 29043 35040 29276 35068
rect 29043 35037 29055 35040
rect 28997 35031 29055 35037
rect 29270 35028 29276 35040
rect 29328 35028 29334 35080
rect 30834 35028 30840 35080
rect 30892 35028 30898 35080
rect 30926 35028 30932 35080
rect 30984 35068 30990 35080
rect 31220 35068 31248 35108
rect 35710 35096 35716 35108
rect 35768 35136 35774 35148
rect 35894 35136 35900 35148
rect 35768 35108 35900 35136
rect 35768 35096 35774 35108
rect 35894 35096 35900 35108
rect 35952 35096 35958 35148
rect 36354 35096 36360 35148
rect 36412 35096 36418 35148
rect 30984 35040 31248 35068
rect 31343 35071 31401 35077
rect 30984 35028 30990 35040
rect 31343 35037 31355 35071
rect 31389 35068 31401 35071
rect 31570 35068 31576 35080
rect 31389 35040 31576 35068
rect 31389 35037 31401 35040
rect 31343 35031 31401 35037
rect 31570 35028 31576 35040
rect 31628 35028 31634 35080
rect 32950 35028 32956 35080
rect 33008 35028 33014 35080
rect 24872 34972 24992 35000
rect 24854 34932 24860 34944
rect 23952 34904 24860 34932
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 24964 34932 24992 34972
rect 25498 34960 25504 35012
rect 25556 35000 25562 35012
rect 26050 35000 26056 35012
rect 25556 34972 26056 35000
rect 25556 34960 25562 34972
rect 26050 34960 26056 34972
rect 26108 35000 26114 35012
rect 26697 35003 26755 35009
rect 26697 35000 26709 35003
rect 26108 34972 26709 35000
rect 26108 34960 26114 34972
rect 26697 34969 26709 34972
rect 26743 34969 26755 35003
rect 26697 34963 26755 34969
rect 26878 34960 26884 35012
rect 26936 34960 26942 35012
rect 31113 35003 31171 35009
rect 31113 34969 31125 35003
rect 31159 34969 31171 35003
rect 31113 34963 31171 34969
rect 25038 34932 25044 34944
rect 24964 34904 25044 34932
rect 25038 34892 25044 34904
rect 25096 34932 25102 34944
rect 25590 34932 25596 34944
rect 25096 34904 25596 34932
rect 25096 34892 25102 34904
rect 25590 34892 25596 34904
rect 25648 34892 25654 34944
rect 25682 34892 25688 34944
rect 25740 34892 25746 34944
rect 27709 34935 27767 34941
rect 27709 34901 27721 34935
rect 27755 34932 27767 34935
rect 28626 34932 28632 34944
rect 27755 34904 28632 34932
rect 27755 34901 27767 34904
rect 27709 34895 27767 34901
rect 28626 34892 28632 34904
rect 28684 34892 28690 34944
rect 30926 34892 30932 34944
rect 30984 34932 30990 34944
rect 31128 34932 31156 34963
rect 31202 34960 31208 35012
rect 31260 34960 31266 35012
rect 32490 34960 32496 35012
rect 32548 35000 32554 35012
rect 32677 35003 32735 35009
rect 32677 35000 32689 35003
rect 32548 34972 32689 35000
rect 32548 34960 32554 34972
rect 32677 34969 32689 34972
rect 32723 34969 32735 35003
rect 34790 35000 34796 35012
rect 32677 34963 32735 34969
rect 32784 34972 34796 35000
rect 30984 34904 31156 34932
rect 31220 34932 31248 34960
rect 32784 34932 32812 34972
rect 34790 34960 34796 34972
rect 34848 34960 34854 35012
rect 36624 35003 36682 35009
rect 36624 34969 36636 35003
rect 36670 35000 36682 35003
rect 37458 35000 37464 35012
rect 36670 34972 37464 35000
rect 36670 34969 36682 34972
rect 36624 34963 36682 34969
rect 37458 34960 37464 34972
rect 37516 34960 37522 35012
rect 31220 34904 32812 34932
rect 32861 34935 32919 34941
rect 30984 34892 30990 34904
rect 32861 34901 32873 34935
rect 32907 34932 32919 34935
rect 33042 34932 33048 34944
rect 32907 34904 33048 34932
rect 32907 34901 32919 34904
rect 32861 34895 32919 34901
rect 33042 34892 33048 34904
rect 33100 34892 33106 34944
rect 37734 34892 37740 34944
rect 37792 34892 37798 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 4614 34728 4620 34740
rect 4356 34700 4620 34728
rect 4356 34601 4384 34700
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 5626 34688 5632 34740
rect 5684 34728 5690 34740
rect 5721 34731 5779 34737
rect 5721 34728 5733 34731
rect 5684 34700 5733 34728
rect 5684 34688 5690 34700
rect 5721 34697 5733 34700
rect 5767 34697 5779 34731
rect 5721 34691 5779 34697
rect 7098 34688 7104 34740
rect 7156 34728 7162 34740
rect 9493 34731 9551 34737
rect 9493 34728 9505 34731
rect 7156 34700 9505 34728
rect 7156 34688 7162 34700
rect 9493 34697 9505 34700
rect 9539 34697 9551 34731
rect 9493 34691 9551 34697
rect 9858 34688 9864 34740
rect 9916 34688 9922 34740
rect 9950 34688 9956 34740
rect 10008 34688 10014 34740
rect 19797 34731 19855 34737
rect 19797 34697 19809 34731
rect 19843 34728 19855 34731
rect 20070 34728 20076 34740
rect 19843 34700 20076 34728
rect 19843 34697 19855 34700
rect 19797 34691 19855 34697
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 20622 34728 20628 34740
rect 20180 34700 20628 34728
rect 5534 34620 5540 34672
rect 5592 34660 5598 34672
rect 5902 34660 5908 34672
rect 5592 34632 5908 34660
rect 5592 34620 5598 34632
rect 5902 34620 5908 34632
rect 5960 34660 5966 34672
rect 20180 34660 20208 34700
rect 20622 34688 20628 34700
rect 20680 34728 20686 34740
rect 20901 34731 20959 34737
rect 20901 34728 20913 34731
rect 20680 34700 20913 34728
rect 20680 34688 20686 34700
rect 20901 34697 20913 34700
rect 20947 34697 20959 34731
rect 20901 34691 20959 34697
rect 22094 34688 22100 34740
rect 22152 34728 22158 34740
rect 24486 34728 24492 34740
rect 22152 34700 24492 34728
rect 22152 34688 22158 34700
rect 24486 34688 24492 34700
rect 24544 34688 24550 34740
rect 25317 34731 25375 34737
rect 25317 34697 25329 34731
rect 25363 34728 25375 34731
rect 27246 34728 27252 34740
rect 25363 34700 27252 34728
rect 25363 34697 25375 34700
rect 25317 34691 25375 34697
rect 27246 34688 27252 34700
rect 27304 34688 27310 34740
rect 28902 34688 28908 34740
rect 28960 34728 28966 34740
rect 30101 34731 30159 34737
rect 30101 34728 30113 34731
rect 28960 34700 30113 34728
rect 28960 34688 28966 34700
rect 30101 34697 30113 34700
rect 30147 34697 30159 34731
rect 30101 34691 30159 34697
rect 31297 34731 31355 34737
rect 31297 34697 31309 34731
rect 31343 34728 31355 34731
rect 31478 34728 31484 34740
rect 31343 34700 31484 34728
rect 31343 34697 31355 34700
rect 31297 34691 31355 34697
rect 31478 34688 31484 34700
rect 31536 34688 31542 34740
rect 32232 34700 32628 34728
rect 5960 34632 7788 34660
rect 5960 34620 5966 34632
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34561 4399 34595
rect 4341 34555 4399 34561
rect 4608 34595 4666 34601
rect 4608 34561 4620 34595
rect 4654 34592 4666 34595
rect 5166 34592 5172 34604
rect 4654 34564 5172 34592
rect 4654 34561 4666 34564
rect 4608 34555 4666 34561
rect 5166 34552 5172 34564
rect 5224 34552 5230 34604
rect 7558 34552 7564 34604
rect 7616 34552 7622 34604
rect 7760 34601 7788 34632
rect 20088 34632 20208 34660
rect 20303 34663 20361 34669
rect 7745 34595 7803 34601
rect 7745 34561 7757 34595
rect 7791 34592 7803 34595
rect 7791 34564 10180 34592
rect 7791 34561 7803 34564
rect 7745 34555 7803 34561
rect 10152 34536 10180 34564
rect 13354 34552 13360 34604
rect 13412 34552 13418 34604
rect 14734 34552 14740 34604
rect 14792 34552 14798 34604
rect 19978 34552 19984 34604
rect 20036 34552 20042 34604
rect 20088 34601 20116 34632
rect 20303 34629 20315 34663
rect 20349 34660 20361 34663
rect 20438 34660 20444 34672
rect 20349 34632 20444 34660
rect 20349 34629 20361 34632
rect 20303 34623 20361 34629
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 26142 34660 26148 34672
rect 21192 34632 26148 34660
rect 20073 34595 20131 34601
rect 20073 34561 20085 34595
rect 20119 34561 20131 34595
rect 20073 34555 20131 34561
rect 20165 34595 20223 34601
rect 20165 34561 20177 34595
rect 20211 34592 20223 34595
rect 20622 34592 20628 34604
rect 20211 34564 20628 34592
rect 20211 34561 20223 34564
rect 20165 34555 20223 34561
rect 20622 34552 20628 34564
rect 20680 34552 20686 34604
rect 21082 34552 21088 34604
rect 21140 34552 21146 34604
rect 7466 34484 7472 34536
rect 7524 34524 7530 34536
rect 7926 34524 7932 34536
rect 7524 34496 7932 34524
rect 7524 34484 7530 34496
rect 7926 34484 7932 34496
rect 7984 34484 7990 34536
rect 8202 34484 8208 34536
rect 8260 34484 8266 34536
rect 10134 34484 10140 34536
rect 10192 34484 10198 34536
rect 12066 34484 12072 34536
rect 12124 34524 12130 34536
rect 13170 34524 13176 34536
rect 12124 34496 13176 34524
rect 12124 34484 12130 34496
rect 13170 34484 13176 34496
rect 13228 34484 13234 34536
rect 13630 34484 13636 34536
rect 13688 34484 13694 34536
rect 15010 34484 15016 34536
rect 15068 34524 15074 34536
rect 15105 34527 15163 34533
rect 15105 34524 15117 34527
rect 15068 34496 15117 34524
rect 15068 34484 15074 34496
rect 15105 34493 15117 34496
rect 15151 34493 15163 34527
rect 15105 34487 15163 34493
rect 19996 34456 20024 34552
rect 20346 34484 20352 34536
rect 20404 34524 20410 34536
rect 20441 34527 20499 34533
rect 20441 34524 20453 34527
rect 20404 34496 20453 34524
rect 20404 34484 20410 34496
rect 20441 34493 20453 34496
rect 20487 34493 20499 34527
rect 20441 34487 20499 34493
rect 20530 34484 20536 34536
rect 20588 34524 20594 34536
rect 20806 34524 20812 34536
rect 20588 34496 20812 34524
rect 20588 34484 20594 34496
rect 20806 34484 20812 34496
rect 20864 34524 20870 34536
rect 21192 34524 21220 34632
rect 26142 34620 26148 34632
rect 26200 34660 26206 34672
rect 26421 34663 26479 34669
rect 26421 34660 26433 34663
rect 26200 34632 26433 34660
rect 26200 34620 26206 34632
rect 26421 34629 26433 34632
rect 26467 34629 26479 34663
rect 26878 34660 26884 34672
rect 26421 34623 26479 34629
rect 26528 34632 26884 34660
rect 21266 34552 21272 34604
rect 21324 34552 21330 34604
rect 21358 34552 21364 34604
rect 21416 34592 21422 34604
rect 23661 34595 23719 34601
rect 23661 34592 23673 34595
rect 21416 34564 23673 34592
rect 21416 34552 21422 34564
rect 23661 34561 23673 34564
rect 23707 34561 23719 34595
rect 23661 34555 23719 34561
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25038 34592 25044 34604
rect 24903 34564 25044 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25130 34552 25136 34604
rect 25188 34552 25194 34604
rect 26050 34552 26056 34604
rect 26108 34592 26114 34604
rect 26237 34595 26295 34601
rect 26237 34592 26249 34595
rect 26108 34564 26249 34592
rect 26108 34552 26114 34564
rect 26237 34561 26249 34564
rect 26283 34592 26295 34595
rect 26528 34592 26556 34632
rect 26878 34620 26884 34632
rect 26936 34620 26942 34672
rect 32232 34660 32260 34700
rect 30852 34632 32260 34660
rect 32309 34663 32367 34669
rect 26283 34564 26556 34592
rect 26605 34595 26663 34601
rect 26283 34561 26295 34564
rect 26237 34555 26295 34561
rect 26605 34561 26617 34595
rect 26651 34592 26663 34595
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 26651 34564 27169 34592
rect 26651 34561 26663 34564
rect 26605 34555 26663 34561
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 27157 34555 27215 34561
rect 29454 34552 29460 34604
rect 29512 34552 29518 34604
rect 30190 34552 30196 34604
rect 30248 34552 30254 34604
rect 30650 34552 30656 34604
rect 30708 34552 30714 34604
rect 30742 34552 30748 34604
rect 30800 34592 30806 34604
rect 30852 34592 30880 34632
rect 32309 34629 32321 34663
rect 32355 34629 32367 34663
rect 32309 34623 32367 34629
rect 30800 34564 30880 34592
rect 30800 34552 30806 34564
rect 30926 34552 30932 34604
rect 30984 34552 30990 34604
rect 31018 34552 31024 34604
rect 31076 34552 31082 34604
rect 31159 34595 31217 34601
rect 31159 34561 31171 34595
rect 31205 34592 31217 34595
rect 31570 34592 31576 34604
rect 31205 34564 31576 34592
rect 31205 34561 31217 34564
rect 31159 34555 31217 34561
rect 31570 34552 31576 34564
rect 31628 34552 31634 34604
rect 32324 34592 32352 34623
rect 32490 34620 32496 34672
rect 32548 34669 32554 34672
rect 32548 34663 32567 34669
rect 32555 34629 32567 34663
rect 32600 34660 32628 34700
rect 32674 34688 32680 34740
rect 32732 34688 32738 34740
rect 37458 34688 37464 34740
rect 37516 34688 37522 34740
rect 33410 34660 33416 34672
rect 32600 34632 33416 34660
rect 32548 34623 32567 34629
rect 32548 34620 32554 34623
rect 33410 34620 33416 34632
rect 33468 34620 33474 34672
rect 33042 34592 33048 34604
rect 32324 34564 33048 34592
rect 33042 34552 33048 34564
rect 33100 34592 33106 34604
rect 33321 34595 33379 34601
rect 33321 34592 33333 34595
rect 33100 34564 33333 34592
rect 33100 34552 33106 34564
rect 33321 34561 33333 34564
rect 33367 34561 33379 34595
rect 33321 34555 33379 34561
rect 34238 34552 34244 34604
rect 34296 34552 34302 34604
rect 34497 34595 34555 34601
rect 34497 34592 34509 34595
rect 34348 34564 34509 34592
rect 20864 34496 21220 34524
rect 21284 34524 21312 34552
rect 22370 34524 22376 34536
rect 21284 34496 22376 34524
rect 20864 34484 20870 34496
rect 22370 34484 22376 34496
rect 22428 34484 22434 34536
rect 22649 34527 22707 34533
rect 22649 34493 22661 34527
rect 22695 34524 22707 34527
rect 23474 34524 23480 34536
rect 22695 34496 23480 34524
rect 22695 34493 22707 34496
rect 22649 34487 22707 34493
rect 23474 34484 23480 34496
rect 23532 34524 23538 34536
rect 23842 34524 23848 34536
rect 23532 34496 23848 34524
rect 23532 34484 23538 34496
rect 23842 34484 23848 34496
rect 23900 34484 23906 34536
rect 24946 34484 24952 34536
rect 25004 34484 25010 34536
rect 27614 34484 27620 34536
rect 27672 34484 27678 34536
rect 31036 34524 31064 34552
rect 32214 34524 32220 34536
rect 31036 34496 32220 34524
rect 32214 34484 32220 34496
rect 32272 34484 32278 34536
rect 32950 34524 32956 34536
rect 32508 34496 32956 34524
rect 20162 34456 20168 34468
rect 19996 34428 20168 34456
rect 20162 34416 20168 34428
rect 20220 34416 20226 34468
rect 20254 34416 20260 34468
rect 20312 34456 20318 34468
rect 20312 34428 22876 34456
rect 20312 34416 20318 34428
rect 17034 34348 17040 34400
rect 17092 34388 17098 34400
rect 22186 34388 22192 34400
rect 17092 34360 22192 34388
rect 17092 34348 17098 34360
rect 22186 34348 22192 34360
rect 22244 34348 22250 34400
rect 22554 34348 22560 34400
rect 22612 34348 22618 34400
rect 22738 34348 22744 34400
rect 22796 34348 22802 34400
rect 22848 34397 22876 34428
rect 23198 34416 23204 34468
rect 23256 34456 23262 34468
rect 23382 34456 23388 34468
rect 23256 34428 23388 34456
rect 23256 34416 23262 34428
rect 23382 34416 23388 34428
rect 23440 34416 23446 34468
rect 23658 34416 23664 34468
rect 23716 34456 23722 34468
rect 31386 34456 31392 34468
rect 23716 34428 31392 34456
rect 23716 34416 23722 34428
rect 31386 34416 31392 34428
rect 31444 34416 31450 34468
rect 22833 34391 22891 34397
rect 22833 34357 22845 34391
rect 22879 34388 22891 34391
rect 24670 34388 24676 34400
rect 22879 34360 24676 34388
rect 22879 34357 22891 34360
rect 22833 34351 22891 34357
rect 24670 34348 24676 34360
rect 24728 34348 24734 34400
rect 25133 34391 25191 34397
rect 25133 34357 25145 34391
rect 25179 34388 25191 34391
rect 25222 34388 25228 34400
rect 25179 34360 25228 34388
rect 25179 34357 25191 34360
rect 25133 34351 25191 34357
rect 25222 34348 25228 34360
rect 25280 34348 25286 34400
rect 29178 34348 29184 34400
rect 29236 34348 29242 34400
rect 32398 34348 32404 34400
rect 32456 34388 32462 34400
rect 32508 34397 32536 34496
rect 32950 34484 32956 34496
rect 33008 34524 33014 34536
rect 33229 34527 33287 34533
rect 33229 34524 33241 34527
rect 33008 34496 33241 34524
rect 33008 34484 33014 34496
rect 33229 34493 33241 34496
rect 33275 34493 33287 34527
rect 33229 34487 33287 34493
rect 33689 34527 33747 34533
rect 33689 34493 33701 34527
rect 33735 34524 33747 34527
rect 34348 34524 34376 34564
rect 34497 34561 34509 34564
rect 34543 34561 34555 34595
rect 34497 34555 34555 34561
rect 37734 34552 37740 34604
rect 37792 34592 37798 34604
rect 37829 34595 37887 34601
rect 37829 34592 37841 34595
rect 37792 34564 37841 34592
rect 37792 34552 37798 34564
rect 37829 34561 37841 34564
rect 37875 34561 37887 34595
rect 37829 34555 37887 34561
rect 33735 34496 34376 34524
rect 37921 34527 37979 34533
rect 33735 34493 33747 34496
rect 33689 34487 33747 34493
rect 37921 34493 37933 34527
rect 37967 34493 37979 34527
rect 37921 34487 37979 34493
rect 37826 34416 37832 34468
rect 37884 34456 37890 34468
rect 37936 34456 37964 34487
rect 38010 34484 38016 34536
rect 38068 34484 38074 34536
rect 37884 34428 37964 34456
rect 37884 34416 37890 34428
rect 32493 34391 32551 34397
rect 32493 34388 32505 34391
rect 32456 34360 32505 34388
rect 32456 34348 32462 34360
rect 32493 34357 32505 34360
rect 32539 34357 32551 34391
rect 32493 34351 32551 34357
rect 35342 34348 35348 34400
rect 35400 34388 35406 34400
rect 35621 34391 35679 34397
rect 35621 34388 35633 34391
rect 35400 34360 35633 34388
rect 35400 34348 35406 34360
rect 35621 34357 35633 34360
rect 35667 34357 35679 34391
rect 35621 34351 35679 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 8294 34144 8300 34196
rect 8352 34184 8358 34196
rect 10413 34187 10471 34193
rect 10413 34184 10425 34187
rect 8352 34156 10425 34184
rect 8352 34144 8358 34156
rect 10413 34153 10425 34156
rect 10459 34153 10471 34187
rect 10413 34147 10471 34153
rect 10873 34187 10931 34193
rect 10873 34153 10885 34187
rect 10919 34184 10931 34187
rect 10919 34156 18644 34184
rect 10919 34153 10931 34156
rect 10873 34147 10931 34153
rect 15010 34076 15016 34128
rect 15068 34116 15074 34128
rect 15068 34088 17540 34116
rect 15068 34076 15074 34088
rect 5534 34008 5540 34060
rect 5592 34008 5598 34060
rect 5626 34008 5632 34060
rect 5684 34008 5690 34060
rect 7668 34020 9444 34048
rect 7374 33940 7380 33992
rect 7432 33980 7438 33992
rect 7668 33989 7696 34020
rect 9416 33992 9444 34020
rect 10594 34008 10600 34060
rect 10652 34008 10658 34060
rect 15286 34008 15292 34060
rect 15344 34048 15350 34060
rect 15344 34020 15608 34048
rect 15344 34008 15350 34020
rect 7653 33983 7711 33989
rect 7653 33980 7665 33983
rect 7432 33952 7665 33980
rect 7432 33940 7438 33952
rect 7653 33949 7665 33952
rect 7699 33949 7711 33983
rect 7653 33943 7711 33949
rect 7834 33940 7840 33992
rect 7892 33940 7898 33992
rect 8202 33940 8208 33992
rect 8260 33980 8266 33992
rect 8481 33983 8539 33989
rect 8481 33980 8493 33983
rect 8260 33952 8493 33980
rect 8260 33940 8266 33952
rect 8481 33949 8493 33952
rect 8527 33980 8539 33983
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 8527 33952 9321 33980
rect 8527 33949 8539 33952
rect 8481 33943 8539 33949
rect 9309 33949 9321 33952
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 9398 33940 9404 33992
rect 9456 33940 9462 33992
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33980 10747 33983
rect 11514 33980 11520 33992
rect 10735 33952 11520 33980
rect 10735 33949 10747 33952
rect 10689 33943 10747 33949
rect 11514 33940 11520 33952
rect 11572 33940 11578 33992
rect 11882 33940 11888 33992
rect 11940 33980 11946 33992
rect 11977 33983 12035 33989
rect 11977 33980 11989 33983
rect 11940 33952 11989 33980
rect 11940 33940 11946 33952
rect 11977 33949 11989 33952
rect 12023 33949 12035 33983
rect 11977 33943 12035 33949
rect 12161 33983 12219 33989
rect 12161 33949 12173 33983
rect 12207 33980 12219 33983
rect 12526 33980 12532 33992
rect 12207 33952 12532 33980
rect 12207 33949 12219 33952
rect 12161 33943 12219 33949
rect 12526 33940 12532 33952
rect 12584 33940 12590 33992
rect 14734 33940 14740 33992
rect 14792 33980 14798 33992
rect 15580 33989 15608 34020
rect 15381 33983 15439 33989
rect 15381 33980 15393 33983
rect 14792 33952 15393 33980
rect 14792 33940 14798 33952
rect 15381 33949 15393 33952
rect 15427 33949 15439 33983
rect 15381 33943 15439 33949
rect 15565 33983 15623 33989
rect 15565 33949 15577 33983
rect 15611 33980 15623 33983
rect 16206 33980 16212 33992
rect 15611 33952 16212 33980
rect 15611 33949 15623 33952
rect 15565 33943 15623 33949
rect 16206 33940 16212 33952
rect 16264 33940 16270 33992
rect 16853 33983 16911 33989
rect 16853 33949 16865 33983
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 5721 33915 5779 33921
rect 5721 33881 5733 33915
rect 5767 33912 5779 33915
rect 6362 33912 6368 33924
rect 5767 33884 6368 33912
rect 5767 33881 5779 33884
rect 5721 33875 5779 33881
rect 6362 33872 6368 33884
rect 6420 33872 6426 33924
rect 9858 33872 9864 33924
rect 9916 33912 9922 33924
rect 10413 33915 10471 33921
rect 10413 33912 10425 33915
rect 9916 33884 10425 33912
rect 9916 33872 9922 33884
rect 10413 33881 10425 33884
rect 10459 33881 10471 33915
rect 10413 33875 10471 33881
rect 13722 33872 13728 33924
rect 13780 33912 13786 33924
rect 16868 33912 16896 33943
rect 17034 33940 17040 33992
rect 17092 33940 17098 33992
rect 17512 33989 17540 34088
rect 18616 33992 18644 34156
rect 20438 34144 20444 34196
rect 20496 34144 20502 34196
rect 21266 34144 21272 34196
rect 21324 34184 21330 34196
rect 22738 34184 22744 34196
rect 21324 34156 22744 34184
rect 21324 34144 21330 34156
rect 22738 34144 22744 34156
rect 22796 34184 22802 34196
rect 23566 34184 23572 34196
rect 22796 34156 23572 34184
rect 22796 34144 22802 34156
rect 23566 34144 23572 34156
rect 23624 34184 23630 34196
rect 23842 34184 23848 34196
rect 23624 34156 23848 34184
rect 23624 34144 23630 34156
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 30377 34187 30435 34193
rect 30377 34153 30389 34187
rect 30423 34184 30435 34187
rect 30834 34184 30840 34196
rect 30423 34156 30840 34184
rect 30423 34153 30435 34156
rect 30377 34147 30435 34153
rect 30834 34144 30840 34156
rect 30892 34144 30898 34196
rect 31849 34187 31907 34193
rect 31849 34153 31861 34187
rect 31895 34184 31907 34187
rect 32490 34184 32496 34196
rect 31895 34156 32496 34184
rect 31895 34153 31907 34156
rect 31849 34147 31907 34153
rect 32490 34144 32496 34156
rect 32548 34144 32554 34196
rect 33134 34144 33140 34196
rect 33192 34184 33198 34196
rect 37642 34184 37648 34196
rect 33192 34156 37648 34184
rect 33192 34144 33198 34156
rect 37642 34144 37648 34156
rect 37700 34144 37706 34196
rect 19613 34119 19671 34125
rect 19613 34085 19625 34119
rect 19659 34116 19671 34119
rect 19978 34116 19984 34128
rect 19659 34088 19984 34116
rect 19659 34085 19671 34088
rect 19613 34079 19671 34085
rect 19978 34076 19984 34088
rect 20036 34076 20042 34128
rect 20254 34076 20260 34128
rect 20312 34116 20318 34128
rect 20530 34116 20536 34128
rect 20312 34088 20536 34116
rect 20312 34076 20318 34088
rect 20530 34076 20536 34088
rect 20588 34076 20594 34128
rect 22646 34076 22652 34128
rect 22704 34116 22710 34128
rect 24946 34116 24952 34128
rect 22704 34088 24952 34116
rect 22704 34076 22710 34088
rect 24946 34076 24952 34088
rect 25004 34076 25010 34128
rect 28074 34076 28080 34128
rect 28132 34116 28138 34128
rect 28718 34116 28724 34128
rect 28132 34088 28724 34116
rect 28132 34076 28138 34088
rect 28718 34076 28724 34088
rect 28776 34076 28782 34128
rect 28902 34076 28908 34128
rect 28960 34076 28966 34128
rect 35710 34116 35716 34128
rect 30024 34088 35716 34116
rect 21177 34051 21235 34057
rect 21177 34048 21189 34051
rect 19444 34020 20024 34048
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33949 17555 33983
rect 18417 33983 18475 33989
rect 18417 33980 18429 33983
rect 17497 33943 17555 33949
rect 17604 33952 18429 33980
rect 17604 33912 17632 33952
rect 18417 33949 18429 33952
rect 18463 33949 18475 33983
rect 18417 33943 18475 33949
rect 18598 33940 18604 33992
rect 18656 33940 18662 33992
rect 19444 33989 19472 34020
rect 19429 33983 19487 33989
rect 19429 33949 19441 33983
rect 19475 33949 19487 33983
rect 19613 33983 19671 33989
rect 19613 33980 19625 33983
rect 19429 33943 19487 33949
rect 19536 33952 19625 33980
rect 13780 33884 17632 33912
rect 13780 33872 13786 33884
rect 17770 33872 17776 33924
rect 17828 33872 17834 33924
rect 17862 33872 17868 33924
rect 17920 33912 17926 33924
rect 19242 33912 19248 33924
rect 17920 33884 19248 33912
rect 17920 33872 17926 33884
rect 19242 33872 19248 33884
rect 19300 33912 19306 33924
rect 19536 33912 19564 33952
rect 19613 33949 19625 33952
rect 19659 33949 19671 33983
rect 19996 33980 20024 34020
rect 20180 34020 21189 34048
rect 20180 33980 20208 34020
rect 21177 34017 21189 34020
rect 21223 34048 21235 34051
rect 21358 34048 21364 34060
rect 21223 34020 21364 34048
rect 21223 34017 21235 34020
rect 21177 34011 21235 34017
rect 21358 34008 21364 34020
rect 21416 34008 21422 34060
rect 22097 34051 22155 34057
rect 22097 34017 22109 34051
rect 22143 34017 22155 34051
rect 24302 34048 24308 34060
rect 22097 34011 22155 34017
rect 23032 34020 24308 34048
rect 19996 33952 20208 33980
rect 19613 33943 19671 33949
rect 20254 33940 20260 33992
rect 20312 33940 20318 33992
rect 20438 33940 20444 33992
rect 20496 33980 20502 33992
rect 20714 33980 20720 33992
rect 20496 33952 20720 33980
rect 20496 33940 20502 33952
rect 20714 33940 20720 33952
rect 20772 33940 20778 33992
rect 21269 33983 21327 33989
rect 21269 33949 21281 33983
rect 21315 33980 21327 33983
rect 22112 33980 22140 34011
rect 23032 33992 23060 34020
rect 24302 34008 24308 34020
rect 24360 34008 24366 34060
rect 24964 34048 24992 34076
rect 26694 34048 26700 34060
rect 24964 34020 26700 34048
rect 21315 33952 22140 33980
rect 21315 33949 21327 33952
rect 21269 33943 21327 33949
rect 22370 33940 22376 33992
rect 22428 33940 22434 33992
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33949 22523 33983
rect 22465 33943 22523 33949
rect 19300 33884 19564 33912
rect 19300 33872 19306 33884
rect 21542 33872 21548 33924
rect 21600 33872 21606 33924
rect 21634 33872 21640 33924
rect 21692 33872 21698 33924
rect 22480 33912 22508 33943
rect 22554 33940 22560 33992
rect 22612 33940 22618 33992
rect 22741 33983 22799 33989
rect 22741 33949 22753 33983
rect 22787 33980 22799 33983
rect 23014 33980 23020 33992
rect 22787 33952 23020 33980
rect 22787 33949 22799 33952
rect 22741 33943 22799 33949
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 23293 33983 23351 33989
rect 23293 33949 23305 33983
rect 23339 33980 23351 33983
rect 23474 33980 23480 33992
rect 23339 33952 23480 33980
rect 23339 33949 23351 33952
rect 23293 33943 23351 33949
rect 23474 33940 23480 33952
rect 23532 33940 23538 33992
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23201 33915 23259 33921
rect 23201 33912 23213 33915
rect 22480 33884 23213 33912
rect 23201 33881 23213 33884
rect 23247 33912 23259 33915
rect 23382 33912 23388 33924
rect 23247 33884 23388 33912
rect 23247 33881 23259 33884
rect 23201 33875 23259 33881
rect 23382 33872 23388 33884
rect 23440 33872 23446 33924
rect 23584 33912 23612 33943
rect 24670 33940 24676 33992
rect 24728 33940 24734 33992
rect 25038 33940 25044 33992
rect 25096 33940 25102 33992
rect 25409 33983 25467 33989
rect 25409 33949 25421 33983
rect 25455 33980 25467 33983
rect 25590 33980 25596 33992
rect 25455 33952 25596 33980
rect 25455 33949 25467 33952
rect 25409 33943 25467 33949
rect 25590 33940 25596 33952
rect 25648 33940 25654 33992
rect 26160 33989 26188 34020
rect 26694 34008 26700 34020
rect 26752 34048 26758 34060
rect 27065 34051 27123 34057
rect 27065 34048 27077 34051
rect 26752 34020 27077 34048
rect 26752 34008 26758 34020
rect 27065 34017 27077 34020
rect 27111 34017 27123 34051
rect 28920 34048 28948 34076
rect 27065 34011 27123 34017
rect 28644 34020 28948 34048
rect 26145 33983 26203 33989
rect 26145 33949 26157 33983
rect 26191 33949 26203 33983
rect 26145 33943 26203 33949
rect 26421 33983 26479 33989
rect 26421 33949 26433 33983
rect 26467 33980 26479 33983
rect 26878 33980 26884 33992
rect 26467 33952 26884 33980
rect 26467 33949 26479 33952
rect 26421 33943 26479 33949
rect 25222 33912 25228 33924
rect 23584 33884 25228 33912
rect 25222 33872 25228 33884
rect 25280 33872 25286 33924
rect 25682 33872 25688 33924
rect 25740 33912 25746 33924
rect 26436 33912 26464 33943
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 28644 33989 28672 34020
rect 28629 33983 28687 33989
rect 28629 33949 28641 33983
rect 28675 33949 28687 33983
rect 28629 33943 28687 33949
rect 28905 33983 28963 33989
rect 28905 33949 28917 33983
rect 28951 33980 28963 33983
rect 29178 33980 29184 33992
rect 28951 33952 29184 33980
rect 28951 33949 28963 33952
rect 28905 33943 28963 33949
rect 29178 33940 29184 33952
rect 29236 33980 29242 33992
rect 29730 33980 29736 33992
rect 29236 33952 29736 33980
rect 29236 33940 29242 33952
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 29822 33940 29828 33992
rect 29880 33980 29886 33992
rect 30024 33980 30052 34088
rect 35710 34076 35716 34088
rect 35768 34076 35774 34128
rect 33226 34048 33232 34060
rect 31496 34020 33232 34048
rect 30282 33989 30288 33992
rect 29880 33952 30052 33980
rect 30239 33983 30288 33989
rect 29880 33940 29886 33952
rect 30239 33949 30251 33983
rect 30285 33949 30288 33983
rect 30239 33943 30288 33949
rect 30282 33940 30288 33943
rect 30340 33940 30346 33992
rect 31202 33940 31208 33992
rect 31260 33940 31266 33992
rect 31353 33983 31411 33989
rect 31353 33949 31365 33983
rect 31399 33980 31411 33983
rect 31496 33980 31524 34020
rect 33226 34008 33232 34020
rect 33284 34048 33290 34060
rect 36078 34048 36084 34060
rect 33284 34020 36084 34048
rect 33284 34008 33290 34020
rect 36078 34008 36084 34020
rect 36136 34008 36142 34060
rect 38102 34008 38108 34060
rect 38160 34008 38166 34060
rect 31662 33980 31668 33992
rect 31720 33989 31726 33992
rect 31399 33952 31524 33980
rect 31628 33952 31668 33980
rect 31399 33949 31411 33952
rect 31353 33943 31411 33949
rect 31662 33940 31668 33952
rect 31720 33943 31728 33989
rect 31720 33940 31726 33943
rect 37826 33940 37832 33992
rect 37884 33940 37890 33992
rect 25740 33884 26464 33912
rect 25740 33872 25746 33884
rect 26510 33872 26516 33924
rect 26568 33872 26574 33924
rect 27614 33872 27620 33924
rect 27672 33912 27678 33924
rect 27893 33915 27951 33921
rect 27893 33912 27905 33915
rect 27672 33884 27905 33912
rect 27672 33872 27678 33884
rect 27893 33881 27905 33884
rect 27939 33881 27951 33915
rect 27893 33875 27951 33881
rect 30006 33872 30012 33924
rect 30064 33872 30070 33924
rect 30098 33872 30104 33924
rect 30156 33872 30162 33924
rect 30300 33884 30512 33912
rect 6086 33804 6092 33856
rect 6144 33804 6150 33856
rect 8754 33804 8760 33856
rect 8812 33844 8818 33856
rect 9125 33847 9183 33853
rect 9125 33844 9137 33847
rect 8812 33816 9137 33844
rect 8812 33804 8818 33816
rect 9125 33813 9137 33816
rect 9171 33813 9183 33847
rect 9125 33807 9183 33813
rect 12069 33847 12127 33853
rect 12069 33813 12081 33847
rect 12115 33844 12127 33847
rect 14182 33844 14188 33856
rect 12115 33816 14188 33844
rect 12115 33813 12127 33816
rect 12069 33807 12127 33813
rect 14182 33804 14188 33816
rect 14240 33804 14246 33856
rect 15470 33804 15476 33856
rect 15528 33804 15534 33856
rect 17037 33847 17095 33853
rect 17037 33813 17049 33847
rect 17083 33844 17095 33847
rect 17586 33844 17592 33856
rect 17083 33816 17592 33844
rect 17083 33813 17095 33816
rect 17037 33807 17095 33813
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 18506 33804 18512 33856
rect 18564 33804 18570 33856
rect 19334 33804 19340 33856
rect 19392 33844 19398 33856
rect 20993 33847 21051 33853
rect 20993 33844 21005 33847
rect 19392 33816 21005 33844
rect 19392 33804 19398 33816
rect 20993 33813 21005 33816
rect 21039 33813 21051 33847
rect 20993 33807 21051 33813
rect 29089 33847 29147 33853
rect 29089 33813 29101 33847
rect 29135 33844 29147 33847
rect 30300 33844 30328 33884
rect 29135 33816 30328 33844
rect 30484 33844 30512 33884
rect 30926 33872 30932 33924
rect 30984 33912 30990 33924
rect 31481 33915 31539 33921
rect 31481 33912 31493 33915
rect 30984 33884 31493 33912
rect 30984 33872 30990 33884
rect 31481 33881 31493 33884
rect 31527 33881 31539 33915
rect 31481 33875 31539 33881
rect 31573 33915 31631 33921
rect 31573 33881 31585 33915
rect 31619 33912 31631 33915
rect 31754 33912 31760 33924
rect 31619 33884 31760 33912
rect 31619 33881 31631 33884
rect 31573 33875 31631 33881
rect 31754 33872 31760 33884
rect 31812 33872 31818 33924
rect 32122 33844 32128 33856
rect 30484 33816 32128 33844
rect 29135 33813 29147 33816
rect 29089 33807 29147 33813
rect 32122 33804 32128 33816
rect 32180 33804 32186 33856
rect 32674 33804 32680 33856
rect 32732 33844 32738 33856
rect 35342 33844 35348 33856
rect 32732 33816 35348 33844
rect 32732 33804 32738 33816
rect 35342 33804 35348 33816
rect 35400 33804 35406 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 13630 33600 13636 33652
rect 13688 33600 13694 33652
rect 14734 33600 14740 33652
rect 14792 33600 14798 33652
rect 16025 33643 16083 33649
rect 15212 33612 15976 33640
rect 7098 33532 7104 33584
rect 7156 33532 7162 33584
rect 9398 33532 9404 33584
rect 9456 33572 9462 33584
rect 15212 33572 15240 33612
rect 9456 33544 10180 33572
rect 9456 33532 9462 33544
rect 5905 33507 5963 33513
rect 5905 33473 5917 33507
rect 5951 33504 5963 33507
rect 6546 33504 6552 33516
rect 5951 33476 6552 33504
rect 5951 33473 5963 33476
rect 5905 33467 5963 33473
rect 6546 33464 6552 33476
rect 6604 33464 6610 33516
rect 8573 33507 8631 33513
rect 8573 33473 8585 33507
rect 8619 33473 8631 33507
rect 8573 33467 8631 33473
rect 5994 33396 6000 33448
rect 6052 33396 6058 33448
rect 6822 33396 6828 33448
rect 6880 33436 6886 33448
rect 8205 33439 8263 33445
rect 8205 33436 8217 33439
rect 6880 33408 8217 33436
rect 6880 33396 6886 33408
rect 8205 33405 8217 33408
rect 8251 33405 8263 33439
rect 8205 33399 8263 33405
rect 6012 33368 6040 33396
rect 7374 33368 7380 33380
rect 6012 33340 7380 33368
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 8386 33328 8392 33380
rect 8444 33368 8450 33380
rect 8588 33368 8616 33467
rect 8754 33464 8760 33516
rect 8812 33464 8818 33516
rect 9674 33464 9680 33516
rect 9732 33464 9738 33516
rect 10152 33513 10180 33544
rect 13280 33544 15240 33572
rect 10137 33507 10195 33513
rect 10137 33473 10149 33507
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 10594 33464 10600 33516
rect 10652 33464 10658 33516
rect 11514 33464 11520 33516
rect 11572 33504 11578 33516
rect 12161 33507 12219 33513
rect 12161 33504 12173 33507
rect 11572 33476 12173 33504
rect 11572 33464 11578 33476
rect 12161 33473 12173 33476
rect 12207 33473 12219 33507
rect 12161 33467 12219 33473
rect 12250 33464 12256 33516
rect 12308 33504 12314 33516
rect 13280 33513 13308 33544
rect 12345 33507 12403 33513
rect 12345 33504 12357 33507
rect 12308 33476 12357 33504
rect 12308 33464 12314 33476
rect 12345 33473 12357 33476
rect 12391 33473 12403 33507
rect 12345 33467 12403 33473
rect 13265 33507 13323 33513
rect 13265 33473 13277 33507
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 13357 33507 13415 33513
rect 13357 33473 13369 33507
rect 13403 33473 13415 33507
rect 13357 33467 13415 33473
rect 13449 33507 13507 33513
rect 13449 33473 13461 33507
rect 13495 33504 13507 33507
rect 14090 33504 14096 33516
rect 13495 33476 14096 33504
rect 13495 33473 13507 33476
rect 13449 33467 13507 33473
rect 9306 33396 9312 33448
rect 9364 33436 9370 33448
rect 9401 33439 9459 33445
rect 9401 33436 9413 33439
rect 9364 33408 9413 33436
rect 9364 33396 9370 33408
rect 9401 33405 9413 33408
rect 9447 33405 9459 33439
rect 9401 33399 9459 33405
rect 10042 33396 10048 33448
rect 10100 33436 10106 33448
rect 10505 33439 10563 33445
rect 10505 33436 10517 33439
rect 10100 33408 10517 33436
rect 10100 33396 10106 33408
rect 10505 33405 10517 33408
rect 10551 33405 10563 33439
rect 13372 33436 13400 33467
rect 14090 33464 14096 33476
rect 14148 33464 14154 33516
rect 14550 33464 14556 33516
rect 14608 33504 14614 33516
rect 15194 33504 15200 33516
rect 14608 33476 15200 33504
rect 14608 33464 14614 33476
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 15378 33464 15384 33516
rect 15436 33464 15442 33516
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33473 15899 33507
rect 15948 33504 15976 33612
rect 16025 33609 16037 33643
rect 16071 33640 16083 33643
rect 16114 33640 16120 33652
rect 16071 33612 16120 33640
rect 16071 33609 16083 33612
rect 16025 33603 16083 33609
rect 16114 33600 16120 33612
rect 16172 33600 16178 33652
rect 16758 33600 16764 33652
rect 16816 33640 16822 33652
rect 17405 33643 17463 33649
rect 17405 33640 17417 33643
rect 16816 33612 17417 33640
rect 16816 33600 16822 33612
rect 17405 33609 17417 33612
rect 17451 33640 17463 33643
rect 17862 33640 17868 33652
rect 17451 33612 17868 33640
rect 17451 33609 17463 33612
rect 17405 33603 17463 33609
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 17954 33600 17960 33652
rect 18012 33640 18018 33652
rect 18966 33640 18972 33652
rect 18012 33612 18972 33640
rect 18012 33600 18018 33612
rect 18966 33600 18972 33612
rect 19024 33600 19030 33652
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 20257 33643 20315 33649
rect 20257 33640 20269 33643
rect 19484 33612 20269 33640
rect 19484 33600 19490 33612
rect 20257 33609 20269 33612
rect 20303 33640 20315 33643
rect 20346 33640 20352 33652
rect 20303 33612 20352 33640
rect 20303 33609 20315 33612
rect 20257 33603 20315 33609
rect 20346 33600 20352 33612
rect 20404 33600 20410 33652
rect 21361 33643 21419 33649
rect 21361 33609 21373 33643
rect 21407 33640 21419 33643
rect 21634 33640 21640 33652
rect 21407 33612 21640 33640
rect 21407 33609 21419 33612
rect 21361 33603 21419 33609
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 25682 33640 25688 33652
rect 22066 33612 25688 33640
rect 16206 33532 16212 33584
rect 16264 33572 16270 33584
rect 19153 33575 19211 33581
rect 19153 33572 19165 33575
rect 16264 33544 19165 33572
rect 16264 33532 16270 33544
rect 19153 33541 19165 33544
rect 19199 33541 19211 33575
rect 19153 33535 19211 33541
rect 19352 33544 20208 33572
rect 16942 33504 16948 33516
rect 15948 33476 16948 33504
rect 15841 33467 15899 33473
rect 13538 33436 13544 33448
rect 13372 33408 13544 33436
rect 10505 33399 10563 33405
rect 13538 33396 13544 33408
rect 13596 33396 13602 33448
rect 14458 33396 14464 33448
rect 14516 33396 14522 33448
rect 15654 33396 15660 33448
rect 15712 33396 15718 33448
rect 10060 33368 10088 33396
rect 8444 33340 10088 33368
rect 12345 33371 12403 33377
rect 8444 33328 8450 33340
rect 12345 33337 12357 33371
rect 12391 33368 12403 33371
rect 15562 33368 15568 33380
rect 12391 33340 15568 33368
rect 12391 33337 12403 33340
rect 12345 33331 12403 33337
rect 15562 33328 15568 33340
rect 15620 33328 15626 33380
rect 15856 33368 15884 33467
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 17770 33464 17776 33516
rect 17828 33504 17834 33516
rect 18141 33507 18199 33513
rect 17828 33476 18092 33504
rect 17828 33464 17834 33476
rect 17681 33439 17739 33445
rect 17681 33405 17693 33439
rect 17727 33436 17739 33439
rect 17954 33436 17960 33448
rect 17727 33408 17960 33436
rect 17727 33405 17739 33408
rect 17681 33399 17739 33405
rect 17954 33396 17960 33408
rect 18012 33396 18018 33448
rect 18064 33436 18092 33476
rect 18141 33473 18153 33507
rect 18187 33504 18199 33507
rect 18690 33504 18696 33516
rect 18187 33476 18696 33504
rect 18187 33473 18199 33476
rect 18141 33467 18199 33473
rect 18690 33464 18696 33476
rect 18748 33504 18754 33516
rect 18874 33504 18880 33516
rect 18748 33476 18880 33504
rect 18748 33464 18754 33476
rect 18874 33464 18880 33476
rect 18932 33464 18938 33516
rect 19352 33513 19380 33544
rect 20180 33516 20208 33544
rect 20530 33532 20536 33584
rect 20588 33572 20594 33584
rect 22066 33572 22094 33612
rect 25682 33600 25688 33612
rect 25740 33600 25746 33652
rect 26602 33640 26608 33652
rect 25792 33612 26608 33640
rect 20588 33544 22094 33572
rect 20588 33532 20594 33544
rect 22370 33532 22376 33584
rect 22428 33572 22434 33584
rect 24857 33575 24915 33581
rect 22428 33544 23520 33572
rect 22428 33532 22434 33544
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33473 19395 33507
rect 19337 33467 19395 33473
rect 19426 33464 19432 33516
rect 19484 33464 19490 33516
rect 19610 33464 19616 33516
rect 19668 33464 19674 33516
rect 19702 33464 19708 33516
rect 19760 33504 19766 33516
rect 19978 33504 19984 33516
rect 19760 33476 19984 33504
rect 19760 33464 19766 33476
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 20162 33464 20168 33516
rect 20220 33464 20226 33516
rect 20441 33507 20499 33513
rect 20441 33473 20453 33507
rect 20487 33473 20499 33507
rect 20441 33467 20499 33473
rect 21453 33507 21511 33513
rect 21453 33473 21465 33507
rect 21499 33504 21511 33507
rect 22388 33504 22416 33532
rect 21499 33476 22416 33504
rect 22465 33507 22523 33513
rect 21499 33473 21511 33476
rect 21453 33467 21511 33473
rect 22465 33473 22477 33507
rect 22511 33504 22523 33507
rect 22830 33504 22836 33516
rect 22511 33476 22836 33504
rect 22511 33473 22523 33476
rect 22465 33467 22523 33473
rect 18233 33439 18291 33445
rect 18233 33436 18245 33439
rect 18064 33408 18245 33436
rect 18233 33405 18245 33408
rect 18279 33436 18291 33439
rect 18414 33436 18420 33448
rect 18279 33408 18420 33436
rect 18279 33405 18291 33408
rect 18233 33399 18291 33405
rect 18414 33396 18420 33408
rect 18472 33396 18478 33448
rect 19886 33396 19892 33448
rect 19944 33436 19950 33448
rect 20456 33436 20484 33467
rect 22830 33464 22836 33476
rect 22888 33464 22894 33516
rect 23109 33507 23167 33513
rect 23109 33473 23121 33507
rect 23155 33504 23167 33507
rect 23382 33504 23388 33516
rect 23155 33476 23388 33504
rect 23155 33473 23167 33476
rect 23109 33467 23167 33473
rect 19944 33408 20484 33436
rect 22373 33439 22431 33445
rect 19944 33396 19950 33408
rect 22373 33405 22385 33439
rect 22419 33436 22431 33439
rect 23124 33436 23152 33467
rect 23382 33464 23388 33476
rect 23440 33464 23446 33516
rect 23492 33504 23520 33544
rect 24857 33541 24869 33575
rect 24903 33572 24915 33575
rect 25590 33572 25596 33584
rect 24903 33544 25596 33572
rect 24903 33541 24915 33544
rect 24857 33535 24915 33541
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 25792 33504 25820 33612
rect 26602 33600 26608 33612
rect 26660 33640 26666 33652
rect 27430 33640 27436 33652
rect 26660 33612 27436 33640
rect 26660 33600 26666 33612
rect 27430 33600 27436 33612
rect 27488 33600 27494 33652
rect 30098 33600 30104 33652
rect 30156 33640 30162 33652
rect 31665 33643 31723 33649
rect 30156 33612 31432 33640
rect 30156 33600 30162 33612
rect 26510 33532 26516 33584
rect 26568 33572 26574 33584
rect 29454 33572 29460 33584
rect 26568 33544 29460 33572
rect 26568 33532 26574 33544
rect 29454 33532 29460 33544
rect 29512 33572 29518 33584
rect 29512 33544 29868 33572
rect 29512 33532 29518 33544
rect 23492 33476 25820 33504
rect 22419 33408 23152 33436
rect 22419 33405 22431 33408
rect 22373 33399 22431 33405
rect 23198 33396 23204 33448
rect 23256 33396 23262 33448
rect 23293 33439 23351 33445
rect 23293 33405 23305 33439
rect 23339 33436 23351 33439
rect 23566 33436 23572 33448
rect 23339 33408 23572 33436
rect 23339 33405 23351 33408
rect 23293 33399 23351 33405
rect 23566 33396 23572 33408
rect 23624 33396 23630 33448
rect 23661 33439 23719 33445
rect 23661 33405 23673 33439
rect 23707 33436 23719 33439
rect 23707 33408 24900 33436
rect 23707 33405 23719 33408
rect 23661 33399 23719 33405
rect 19610 33368 19616 33380
rect 15856 33340 19616 33368
rect 19610 33328 19616 33340
rect 19668 33328 19674 33380
rect 24872 33312 24900 33408
rect 25130 33396 25136 33448
rect 25188 33436 25194 33448
rect 25225 33439 25283 33445
rect 25225 33436 25237 33439
rect 25188 33408 25237 33436
rect 25188 33396 25194 33408
rect 25225 33405 25237 33408
rect 25271 33405 25283 33439
rect 25225 33399 25283 33405
rect 25593 33439 25651 33445
rect 25593 33405 25605 33439
rect 25639 33436 25651 33439
rect 25792 33436 25820 33476
rect 26142 33464 26148 33516
rect 26200 33464 26206 33516
rect 27433 33507 27491 33513
rect 27433 33504 27445 33507
rect 26252 33476 27445 33504
rect 25639 33408 25820 33436
rect 25639 33405 25651 33408
rect 25593 33399 25651 33405
rect 25774 33368 25780 33380
rect 25148 33340 25780 33368
rect 5626 33260 5632 33312
rect 5684 33300 5690 33312
rect 5721 33303 5779 33309
rect 5721 33300 5733 33303
rect 5684 33272 5733 33300
rect 5684 33260 5690 33272
rect 5721 33269 5733 33272
rect 5767 33269 5779 33303
rect 5721 33263 5779 33269
rect 6546 33260 6552 33312
rect 6604 33300 6610 33312
rect 7193 33303 7251 33309
rect 7193 33300 7205 33303
rect 6604 33272 7205 33300
rect 6604 33260 6610 33272
rect 7193 33269 7205 33272
rect 7239 33269 7251 33303
rect 7193 33263 7251 33269
rect 14182 33260 14188 33312
rect 14240 33260 14246 33312
rect 15470 33260 15476 33312
rect 15528 33260 15534 33312
rect 17773 33303 17831 33309
rect 17773 33269 17785 33303
rect 17819 33300 17831 33303
rect 18322 33300 18328 33312
rect 17819 33272 18328 33300
rect 17819 33269 17831 33272
rect 17773 33263 17831 33269
rect 18322 33260 18328 33272
rect 18380 33260 18386 33312
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20625 33303 20683 33309
rect 20625 33300 20637 33303
rect 20036 33272 20637 33300
rect 20036 33260 20042 33272
rect 20625 33269 20637 33272
rect 20671 33269 20683 33303
rect 20625 33263 20683 33269
rect 22097 33303 22155 33309
rect 22097 33269 22109 33303
rect 22143 33300 22155 33303
rect 22186 33300 22192 33312
rect 22143 33272 22192 33300
rect 22143 33269 22155 33272
rect 22097 33263 22155 33269
rect 22186 33260 22192 33272
rect 22244 33260 22250 33312
rect 22465 33303 22523 33309
rect 22465 33269 22477 33303
rect 22511 33300 22523 33303
rect 22646 33300 22652 33312
rect 22511 33272 22652 33300
rect 22511 33269 22523 33272
rect 22465 33263 22523 33269
rect 22646 33260 22652 33272
rect 22704 33260 22710 33312
rect 24854 33260 24860 33312
rect 24912 33300 24918 33312
rect 25148 33309 25176 33340
rect 25774 33328 25780 33340
rect 25832 33328 25838 33380
rect 24995 33303 25053 33309
rect 24995 33300 25007 33303
rect 24912 33272 25007 33300
rect 24912 33260 24918 33272
rect 24995 33269 25007 33272
rect 25041 33269 25053 33303
rect 24995 33263 25053 33269
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25222 33300 25228 33312
rect 25179 33272 25228 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25222 33260 25228 33272
rect 25280 33260 25286 33312
rect 25866 33260 25872 33312
rect 25924 33300 25930 33312
rect 26252 33309 26280 33476
rect 27433 33473 27445 33476
rect 27479 33473 27491 33507
rect 27433 33467 27491 33473
rect 28626 33464 28632 33516
rect 28684 33464 28690 33516
rect 29840 33513 29868 33544
rect 30926 33532 30932 33584
rect 30984 33572 30990 33584
rect 31297 33575 31355 33581
rect 31297 33572 31309 33575
rect 30984 33544 31309 33572
rect 30984 33532 30990 33544
rect 31297 33541 31309 33544
rect 31343 33541 31355 33575
rect 31404 33572 31432 33612
rect 31665 33609 31677 33643
rect 31711 33640 31723 33643
rect 32398 33640 32404 33652
rect 31711 33612 32404 33640
rect 31711 33609 31723 33612
rect 31665 33603 31723 33609
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 33336 33612 34376 33640
rect 33336 33572 33364 33612
rect 31404 33544 33364 33572
rect 31297 33535 31355 33541
rect 33410 33532 33416 33584
rect 33468 33532 33474 33584
rect 34348 33572 34376 33612
rect 34422 33600 34428 33652
rect 34480 33640 34486 33652
rect 35986 33640 35992 33652
rect 34480 33612 35992 33640
rect 34480 33600 34486 33612
rect 35986 33600 35992 33612
rect 36044 33600 36050 33652
rect 36173 33643 36231 33649
rect 36173 33609 36185 33643
rect 36219 33640 36231 33643
rect 37826 33640 37832 33652
rect 36219 33612 37832 33640
rect 36219 33609 36231 33612
rect 36173 33603 36231 33609
rect 37826 33600 37832 33612
rect 37884 33600 37890 33652
rect 37918 33572 37924 33584
rect 34348 33544 34560 33572
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 29825 33467 29883 33473
rect 31018 33464 31024 33516
rect 31076 33464 31082 33516
rect 31114 33507 31172 33513
rect 31114 33473 31126 33507
rect 31160 33473 31172 33507
rect 31114 33467 31172 33473
rect 26326 33396 26332 33448
rect 26384 33436 26390 33448
rect 26421 33439 26479 33445
rect 26421 33436 26433 33439
rect 26384 33408 26433 33436
rect 26384 33396 26390 33408
rect 26421 33405 26433 33408
rect 26467 33405 26479 33439
rect 26421 33399 26479 33405
rect 27154 33396 27160 33448
rect 27212 33436 27218 33448
rect 27709 33439 27767 33445
rect 27709 33436 27721 33439
rect 27212 33408 27721 33436
rect 27212 33396 27218 33408
rect 27709 33405 27721 33408
rect 27755 33405 27767 33439
rect 27709 33399 27767 33405
rect 28994 33396 29000 33448
rect 29052 33396 29058 33448
rect 30282 33396 30288 33448
rect 30340 33396 30346 33448
rect 31128 33436 31156 33467
rect 31386 33464 31392 33516
rect 31444 33464 31450 33516
rect 31570 33513 31576 33516
rect 31527 33507 31576 33513
rect 31527 33473 31539 33507
rect 31573 33473 31576 33507
rect 31527 33467 31576 33473
rect 31570 33464 31576 33467
rect 31628 33464 31634 33516
rect 33042 33464 33048 33516
rect 33100 33464 33106 33516
rect 33134 33464 33140 33516
rect 33192 33504 33198 33516
rect 33321 33507 33379 33513
rect 33192 33476 33237 33504
rect 33192 33464 33198 33476
rect 33321 33473 33333 33507
rect 33367 33473 33379 33507
rect 33321 33467 33379 33473
rect 33551 33507 33609 33513
rect 33551 33473 33563 33507
rect 33597 33504 33609 33507
rect 34422 33504 34428 33516
rect 33597 33476 34428 33504
rect 33597 33473 33609 33476
rect 33551 33467 33609 33473
rect 32674 33436 32680 33448
rect 31128 33408 32680 33436
rect 28626 33328 28632 33380
rect 28684 33368 28690 33380
rect 31128 33368 31156 33408
rect 32674 33396 32680 33408
rect 32732 33396 32738 33448
rect 28684 33340 31156 33368
rect 28684 33328 28690 33340
rect 26237 33303 26295 33309
rect 26237 33300 26249 33303
rect 25924 33272 26249 33300
rect 25924 33260 25930 33272
rect 26237 33269 26249 33272
rect 26283 33269 26295 33303
rect 33336 33300 33364 33467
rect 34422 33464 34428 33476
rect 34480 33464 34486 33516
rect 34532 33513 34560 33544
rect 34624 33544 37924 33572
rect 34517 33507 34575 33513
rect 34517 33473 34529 33507
rect 34563 33473 34575 33507
rect 34517 33467 34575 33473
rect 34624 33436 34652 33544
rect 37918 33532 37924 33544
rect 37976 33532 37982 33584
rect 34698 33464 34704 33516
rect 34756 33464 34762 33516
rect 34790 33464 34796 33516
rect 34848 33464 34854 33516
rect 34885 33507 34943 33513
rect 34885 33473 34897 33507
rect 34931 33473 34943 33507
rect 35529 33507 35587 33513
rect 35529 33504 35541 33507
rect 34885 33467 34943 33473
rect 35084 33476 35541 33504
rect 34900 33436 34928 33467
rect 33704 33408 34652 33436
rect 34716 33408 34928 33436
rect 33704 33377 33732 33408
rect 34716 33380 34744 33408
rect 33689 33371 33747 33377
rect 33689 33337 33701 33371
rect 33735 33337 33747 33371
rect 33689 33331 33747 33337
rect 34698 33328 34704 33380
rect 34756 33328 34762 33380
rect 35084 33377 35112 33476
rect 35529 33473 35541 33476
rect 35575 33473 35587 33507
rect 35529 33467 35587 33473
rect 35622 33507 35680 33513
rect 35622 33473 35634 33507
rect 35668 33473 35680 33507
rect 35622 33467 35680 33473
rect 35636 33436 35664 33467
rect 35802 33464 35808 33516
rect 35860 33464 35866 33516
rect 35894 33464 35900 33516
rect 35952 33464 35958 33516
rect 35986 33464 35992 33516
rect 36044 33513 36050 33516
rect 36044 33507 36093 33513
rect 36044 33473 36047 33507
rect 36081 33504 36093 33507
rect 36262 33504 36268 33516
rect 36081 33476 36268 33504
rect 36081 33473 36093 33476
rect 36044 33467 36093 33473
rect 36044 33464 36050 33467
rect 36262 33464 36268 33476
rect 36320 33464 36326 33516
rect 37826 33464 37832 33516
rect 37884 33464 37890 33516
rect 35710 33436 35716 33448
rect 35636 33408 35716 33436
rect 35710 33396 35716 33408
rect 35768 33436 35774 33448
rect 37734 33436 37740 33448
rect 35768 33408 37740 33436
rect 35768 33396 35774 33408
rect 37734 33396 37740 33408
rect 37792 33396 37798 33448
rect 37918 33396 37924 33448
rect 37976 33396 37982 33448
rect 38010 33396 38016 33448
rect 38068 33396 38074 33448
rect 35069 33371 35127 33377
rect 35069 33337 35081 33371
rect 35115 33337 35127 33371
rect 35069 33331 35127 33337
rect 35802 33300 35808 33312
rect 33336 33272 35808 33300
rect 26237 33263 26295 33269
rect 35802 33260 35808 33272
rect 35860 33260 35866 33312
rect 37090 33260 37096 33312
rect 37148 33300 37154 33312
rect 37461 33303 37519 33309
rect 37461 33300 37473 33303
rect 37148 33272 37473 33300
rect 37148 33260 37154 33272
rect 37461 33269 37473 33272
rect 37507 33269 37519 33303
rect 37461 33263 37519 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 4982 33056 4988 33108
rect 5040 33096 5046 33108
rect 5445 33099 5503 33105
rect 5445 33096 5457 33099
rect 5040 33068 5457 33096
rect 5040 33056 5046 33068
rect 5445 33065 5457 33068
rect 5491 33065 5503 33099
rect 5445 33059 5503 33065
rect 7561 33099 7619 33105
rect 7561 33065 7573 33099
rect 7607 33096 7619 33099
rect 8754 33096 8760 33108
rect 7607 33068 8760 33096
rect 7607 33065 7619 33068
rect 7561 33059 7619 33065
rect 8754 33056 8760 33068
rect 8812 33056 8818 33108
rect 10781 33099 10839 33105
rect 10781 33096 10793 33099
rect 9692 33068 10793 33096
rect 9692 33040 9720 33068
rect 10781 33065 10793 33068
rect 10827 33065 10839 33099
rect 10781 33059 10839 33065
rect 11241 33099 11299 33105
rect 11241 33065 11253 33099
rect 11287 33096 11299 33099
rect 13722 33096 13728 33108
rect 11287 33068 13728 33096
rect 11287 33065 11299 33068
rect 11241 33059 11299 33065
rect 13722 33056 13728 33068
rect 13780 33056 13786 33108
rect 14090 33056 14096 33108
rect 14148 33096 14154 33108
rect 14369 33099 14427 33105
rect 14369 33096 14381 33099
rect 14148 33068 14381 33096
rect 14148 33056 14154 33068
rect 14369 33065 14381 33068
rect 14415 33065 14427 33099
rect 14369 33059 14427 33065
rect 15286 33056 15292 33108
rect 15344 33056 15350 33108
rect 15657 33099 15715 33105
rect 15657 33065 15669 33099
rect 15703 33096 15715 33099
rect 15838 33096 15844 33108
rect 15703 33068 15844 33096
rect 15703 33065 15715 33068
rect 15657 33059 15715 33065
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 17589 33099 17647 33105
rect 17589 33065 17601 33099
rect 17635 33065 17647 33099
rect 17589 33059 17647 33065
rect 17773 33099 17831 33105
rect 17773 33065 17785 33099
rect 17819 33096 17831 33099
rect 18046 33096 18052 33108
rect 17819 33068 18052 33096
rect 17819 33065 17831 33068
rect 17773 33059 17831 33065
rect 6917 33031 6975 33037
rect 6917 32997 6929 33031
rect 6963 33028 6975 33031
rect 9674 33028 9680 33040
rect 6963 33000 9680 33028
rect 6963 32997 6975 33000
rect 6917 32991 6975 32997
rect 9674 32988 9680 33000
rect 9732 32988 9738 33040
rect 10134 32988 10140 33040
rect 10192 33028 10198 33040
rect 10321 33031 10379 33037
rect 10321 33028 10333 33031
rect 10192 33000 10333 33028
rect 10192 32988 10198 33000
rect 10321 32997 10333 33000
rect 10367 33028 10379 33031
rect 12345 33031 12403 33037
rect 12345 33028 12357 33031
rect 10367 33000 12357 33028
rect 10367 32997 10379 33000
rect 10321 32991 10379 32997
rect 12345 32997 12357 33000
rect 12391 32997 12403 33031
rect 17604 33028 17632 33059
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 18230 33056 18236 33108
rect 18288 33096 18294 33108
rect 18325 33099 18383 33105
rect 18325 33096 18337 33099
rect 18288 33068 18337 33096
rect 18288 33056 18294 33068
rect 18325 33065 18337 33068
rect 18371 33065 18383 33099
rect 22738 33096 22744 33108
rect 18325 33059 18383 33065
rect 19444 33068 22744 33096
rect 19334 33028 19340 33040
rect 12345 32991 12403 32997
rect 13740 33000 17540 33028
rect 17604 33000 19340 33028
rect 5994 32960 6000 32972
rect 5184 32932 6000 32960
rect 4522 32852 4528 32904
rect 4580 32892 4586 32904
rect 5184 32901 5212 32932
rect 5994 32920 6000 32932
rect 6052 32920 6058 32972
rect 7745 32963 7803 32969
rect 7745 32929 7757 32963
rect 7791 32960 7803 32963
rect 7791 32932 8432 32960
rect 7791 32929 7803 32932
rect 7745 32923 7803 32929
rect 8404 32904 8432 32932
rect 10594 32920 10600 32972
rect 10652 32960 10658 32972
rect 10873 32963 10931 32969
rect 10873 32960 10885 32963
rect 10652 32932 10885 32960
rect 10652 32920 10658 32932
rect 10873 32929 10885 32932
rect 10919 32929 10931 32963
rect 10873 32923 10931 32929
rect 5169 32895 5227 32901
rect 5169 32892 5181 32895
rect 4580 32864 5181 32892
rect 4580 32852 4586 32864
rect 5169 32861 5181 32864
rect 5215 32861 5227 32895
rect 5169 32855 5227 32861
rect 5258 32852 5264 32904
rect 5316 32852 5322 32904
rect 6546 32852 6552 32904
rect 6604 32892 6610 32904
rect 6825 32895 6883 32901
rect 6825 32892 6837 32895
rect 6604 32864 6837 32892
rect 6604 32852 6610 32864
rect 6825 32861 6837 32864
rect 6871 32861 6883 32895
rect 6825 32855 6883 32861
rect 7009 32895 7067 32901
rect 7009 32861 7021 32895
rect 7055 32892 7067 32895
rect 7374 32892 7380 32904
rect 7055 32864 7380 32892
rect 7055 32861 7067 32864
rect 7009 32855 7067 32861
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 7469 32895 7527 32901
rect 7469 32861 7481 32895
rect 7515 32861 7527 32895
rect 7469 32855 7527 32861
rect 6178 32784 6184 32836
rect 6236 32824 6242 32836
rect 7484 32824 7512 32855
rect 7558 32852 7564 32904
rect 7616 32892 7622 32904
rect 7834 32892 7840 32904
rect 7616 32864 7840 32892
rect 7616 32852 7622 32864
rect 7834 32852 7840 32864
rect 7892 32892 7898 32904
rect 7892 32864 8340 32892
rect 7892 32852 7898 32864
rect 6236 32796 7512 32824
rect 6236 32784 6242 32796
rect 8110 32784 8116 32836
rect 8168 32824 8174 32836
rect 8205 32827 8263 32833
rect 8205 32824 8217 32827
rect 8168 32796 8217 32824
rect 8168 32784 8174 32796
rect 8205 32793 8217 32796
rect 8251 32793 8263 32827
rect 8312 32824 8340 32864
rect 8386 32852 8392 32904
rect 8444 32852 8450 32904
rect 9858 32892 9864 32904
rect 8588 32864 9864 32892
rect 8588 32833 8616 32864
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 10042 32852 10048 32904
rect 10100 32892 10106 32904
rect 10137 32895 10195 32901
rect 10137 32892 10149 32895
rect 10100 32864 10149 32892
rect 10100 32852 10106 32864
rect 10137 32861 10149 32864
rect 10183 32861 10195 32895
rect 10137 32855 10195 32861
rect 11057 32895 11115 32901
rect 11057 32861 11069 32895
rect 11103 32892 11115 32895
rect 11514 32892 11520 32904
rect 11103 32864 11520 32892
rect 11103 32861 11115 32864
rect 11057 32855 11115 32861
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 12253 32895 12311 32901
rect 12253 32861 12265 32895
rect 12299 32861 12311 32895
rect 12253 32855 12311 32861
rect 8573 32827 8631 32833
rect 8573 32824 8585 32827
rect 8312 32796 8585 32824
rect 8205 32787 8263 32793
rect 8573 32793 8585 32796
rect 8619 32793 8631 32827
rect 9876 32824 9904 32852
rect 10781 32827 10839 32833
rect 10781 32824 10793 32827
rect 9876 32796 10793 32824
rect 8573 32787 8631 32793
rect 10781 32793 10793 32796
rect 10827 32793 10839 32827
rect 12268 32824 12296 32855
rect 12434 32852 12440 32904
rect 12492 32852 12498 32904
rect 12526 32852 12532 32904
rect 12584 32852 12590 32904
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32892 12771 32895
rect 13538 32892 13544 32904
rect 12759 32864 13544 32892
rect 12759 32861 12771 32864
rect 12713 32855 12771 32861
rect 13538 32852 13544 32864
rect 13596 32852 13602 32904
rect 13740 32901 13768 33000
rect 14553 32963 14611 32969
rect 14553 32929 14565 32963
rect 14599 32960 14611 32963
rect 14826 32960 14832 32972
rect 14599 32932 14832 32960
rect 14599 32929 14611 32932
rect 14553 32923 14611 32929
rect 14826 32920 14832 32932
rect 14884 32920 14890 32972
rect 15470 32960 15476 32972
rect 15120 32932 15476 32960
rect 13725 32895 13783 32901
rect 13725 32861 13737 32895
rect 13771 32861 13783 32895
rect 14645 32895 14703 32901
rect 14645 32892 14657 32895
rect 13725 32855 13783 32861
rect 14568 32864 14657 32892
rect 12544 32824 12572 32852
rect 14568 32836 14596 32864
rect 14645 32861 14657 32864
rect 14691 32861 14703 32895
rect 14645 32855 14703 32861
rect 14734 32852 14740 32904
rect 14792 32892 14798 32904
rect 15120 32892 15148 32932
rect 15470 32920 15476 32932
rect 15528 32920 15534 32972
rect 17218 32920 17224 32972
rect 17276 32960 17282 32972
rect 17405 32963 17463 32969
rect 17405 32960 17417 32963
rect 17276 32932 17417 32960
rect 17276 32920 17282 32932
rect 17405 32929 17417 32932
rect 17451 32929 17463 32963
rect 17512 32960 17540 33000
rect 19334 32988 19340 33000
rect 19392 32988 19398 33040
rect 18509 32963 18567 32969
rect 17512 32932 18460 32960
rect 17405 32923 17463 32929
rect 14792 32864 15148 32892
rect 14792 32852 14798 32864
rect 15194 32852 15200 32904
rect 15252 32892 15258 32904
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 15252 32864 15301 32892
rect 15252 32852 15258 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 15289 32855 15347 32861
rect 15381 32895 15439 32901
rect 15381 32861 15393 32895
rect 15427 32861 15439 32895
rect 15381 32855 15439 32861
rect 12802 32824 12808 32836
rect 12268 32796 12434 32824
rect 12544 32796 12808 32824
rect 10781 32787 10839 32793
rect 7745 32759 7803 32765
rect 7745 32725 7757 32759
rect 7791 32756 7803 32759
rect 9490 32756 9496 32768
rect 7791 32728 9496 32756
rect 7791 32725 7803 32728
rect 7745 32719 7803 32725
rect 9490 32716 9496 32728
rect 9548 32716 9554 32768
rect 9953 32759 10011 32765
rect 9953 32725 9965 32759
rect 9999 32756 10011 32759
rect 10594 32756 10600 32768
rect 9999 32728 10600 32756
rect 9999 32725 10011 32728
rect 9953 32719 10011 32725
rect 10594 32716 10600 32728
rect 10652 32716 10658 32768
rect 12406 32756 12434 32796
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 14550 32784 14556 32836
rect 14608 32824 14614 32836
rect 15396 32824 15424 32855
rect 15562 32852 15568 32904
rect 15620 32892 15626 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 15620 32864 17325 32892
rect 15620 32852 15626 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17313 32855 17371 32861
rect 17586 32852 17592 32904
rect 17644 32852 17650 32904
rect 18233 32895 18291 32901
rect 18233 32861 18245 32895
rect 18279 32892 18291 32895
rect 18322 32892 18328 32904
rect 18279 32864 18328 32892
rect 18279 32861 18291 32864
rect 18233 32855 18291 32861
rect 18322 32852 18328 32864
rect 18380 32852 18386 32904
rect 18432 32892 18460 32932
rect 18509 32929 18521 32963
rect 18555 32960 18567 32963
rect 18598 32960 18604 32972
rect 18555 32932 18604 32960
rect 18555 32929 18567 32932
rect 18509 32923 18567 32929
rect 18598 32920 18604 32932
rect 18656 32920 18662 32972
rect 19444 32892 19472 33068
rect 22738 33056 22744 33068
rect 22796 33056 22802 33108
rect 25225 33099 25283 33105
rect 25225 33065 25237 33099
rect 25271 33096 25283 33099
rect 25682 33096 25688 33108
rect 25271 33068 25688 33096
rect 25271 33065 25283 33068
rect 25225 33059 25283 33065
rect 25682 33056 25688 33068
rect 25740 33056 25746 33108
rect 30377 33099 30435 33105
rect 30377 33065 30389 33099
rect 30423 33096 30435 33099
rect 30650 33096 30656 33108
rect 30423 33068 30656 33096
rect 30423 33065 30435 33068
rect 30377 33059 30435 33065
rect 30650 33056 30656 33068
rect 30708 33056 30714 33108
rect 30837 33099 30895 33105
rect 30837 33065 30849 33099
rect 30883 33096 30895 33099
rect 31202 33096 31208 33108
rect 30883 33068 31208 33096
rect 30883 33065 30895 33068
rect 30837 33059 30895 33065
rect 31202 33056 31208 33068
rect 31260 33056 31266 33108
rect 31294 33056 31300 33108
rect 31352 33096 31358 33108
rect 32493 33099 32551 33105
rect 31352 33068 32444 33096
rect 31352 33056 31358 33068
rect 20346 32988 20352 33040
rect 20404 33028 20410 33040
rect 20714 33028 20720 33040
rect 20404 33000 20720 33028
rect 20404 32988 20410 33000
rect 20714 32988 20720 33000
rect 20772 32988 20778 33040
rect 25406 32988 25412 33040
rect 25464 32988 25470 33040
rect 27614 33028 27620 33040
rect 26252 33000 27620 33028
rect 20254 32960 20260 32972
rect 19628 32932 20260 32960
rect 19628 32901 19656 32932
rect 20254 32920 20260 32932
rect 20312 32920 20318 32972
rect 20548 32960 20668 32968
rect 20456 32940 20668 32960
rect 20456 32932 20576 32940
rect 18432 32864 19472 32892
rect 19613 32895 19671 32901
rect 19613 32861 19625 32895
rect 19659 32861 19671 32895
rect 19613 32855 19671 32861
rect 19797 32895 19855 32901
rect 19797 32861 19809 32895
rect 19843 32861 19855 32895
rect 19797 32855 19855 32861
rect 14608 32796 15424 32824
rect 19812 32824 19840 32855
rect 20346 32852 20352 32904
rect 20404 32892 20410 32904
rect 20456 32901 20484 32932
rect 20441 32895 20499 32901
rect 20441 32892 20453 32895
rect 20404 32864 20453 32892
rect 20404 32852 20410 32864
rect 20441 32861 20453 32864
rect 20487 32861 20499 32895
rect 20441 32855 20499 32861
rect 20530 32852 20536 32904
rect 20588 32852 20594 32904
rect 20640 32892 20668 32940
rect 20901 32963 20959 32969
rect 20901 32929 20913 32963
rect 20947 32960 20959 32963
rect 21634 32960 21640 32972
rect 20947 32932 21640 32960
rect 20947 32929 20959 32932
rect 20901 32923 20959 32929
rect 21634 32920 21640 32932
rect 21692 32920 21698 32972
rect 22830 32920 22836 32972
rect 22888 32960 22894 32972
rect 23109 32963 23167 32969
rect 22888 32932 23060 32960
rect 22888 32920 22894 32932
rect 22554 32892 22560 32904
rect 20640 32864 22560 32892
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22922 32852 22928 32904
rect 22980 32852 22986 32904
rect 23032 32892 23060 32932
rect 23109 32929 23121 32963
rect 23155 32960 23167 32963
rect 23382 32960 23388 32972
rect 23155 32932 23388 32960
rect 23155 32929 23167 32932
rect 23109 32923 23167 32929
rect 23382 32920 23388 32932
rect 23440 32920 23446 32972
rect 24765 32963 24823 32969
rect 24765 32929 24777 32963
rect 24811 32960 24823 32963
rect 24946 32960 24952 32972
rect 24811 32932 24952 32960
rect 24811 32929 24823 32932
rect 24765 32923 24823 32929
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 26252 32960 26280 33000
rect 27614 32988 27620 33000
rect 27672 32988 27678 33040
rect 30282 33028 30288 33040
rect 29748 33000 30288 33028
rect 25332 32932 26280 32960
rect 23201 32895 23259 32901
rect 23032 32886 23152 32892
rect 23201 32886 23213 32895
rect 23032 32864 23213 32886
rect 23124 32861 23213 32864
rect 23247 32861 23259 32895
rect 23124 32858 23259 32861
rect 23201 32855 23259 32858
rect 24578 32852 24584 32904
rect 24636 32892 24642 32904
rect 24857 32895 24915 32901
rect 24857 32892 24869 32895
rect 24636 32864 24869 32892
rect 24636 32852 24642 32864
rect 24857 32861 24869 32864
rect 24903 32861 24915 32895
rect 24857 32855 24915 32861
rect 25222 32852 25228 32904
rect 25280 32852 25286 32904
rect 20548 32824 20576 32852
rect 19812 32796 20576 32824
rect 14608 32784 14614 32796
rect 20806 32784 20812 32836
rect 20864 32784 20870 32836
rect 25332 32824 25360 32932
rect 26234 32892 26240 32904
rect 22066 32796 25360 32824
rect 25424 32864 26240 32892
rect 13630 32756 13636 32768
rect 12406 32728 13636 32756
rect 13630 32716 13636 32728
rect 13688 32716 13694 32768
rect 13725 32759 13783 32765
rect 13725 32725 13737 32759
rect 13771 32756 13783 32759
rect 14274 32756 14280 32768
rect 13771 32728 14280 32756
rect 13771 32725 13783 32728
rect 13725 32719 13783 32725
rect 14274 32716 14280 32728
rect 14332 32716 14338 32768
rect 14366 32716 14372 32768
rect 14424 32756 14430 32768
rect 18414 32756 18420 32768
rect 14424 32728 18420 32756
rect 14424 32716 14430 32728
rect 18414 32716 18420 32728
rect 18472 32716 18478 32768
rect 18509 32759 18567 32765
rect 18509 32725 18521 32759
rect 18555 32756 18567 32759
rect 19334 32756 19340 32768
rect 18555 32728 19340 32756
rect 18555 32725 18567 32728
rect 18509 32719 18567 32725
rect 19334 32716 19340 32728
rect 19392 32716 19398 32768
rect 19426 32716 19432 32768
rect 19484 32756 19490 32768
rect 19705 32759 19763 32765
rect 19705 32756 19717 32759
rect 19484 32728 19717 32756
rect 19484 32716 19490 32728
rect 19705 32725 19717 32728
rect 19751 32756 19763 32759
rect 19886 32756 19892 32768
rect 19751 32728 19892 32756
rect 19751 32725 19763 32728
rect 19705 32719 19763 32725
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 20254 32716 20260 32768
rect 20312 32716 20318 32768
rect 20898 32716 20904 32768
rect 20956 32756 20962 32768
rect 22066 32756 22094 32796
rect 20956 32728 22094 32756
rect 20956 32716 20962 32728
rect 22738 32716 22744 32768
rect 22796 32716 22802 32768
rect 23566 32716 23572 32768
rect 23624 32756 23630 32768
rect 25424 32756 25452 32864
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 26694 32852 26700 32904
rect 26752 32852 26758 32904
rect 27801 32895 27859 32901
rect 27801 32861 27813 32895
rect 27847 32861 27859 32895
rect 27801 32855 27859 32861
rect 26050 32784 26056 32836
rect 26108 32824 26114 32836
rect 27816 32824 27844 32855
rect 28166 32852 28172 32904
rect 28224 32852 28230 32904
rect 28718 32852 28724 32904
rect 28776 32852 28782 32904
rect 29748 32901 29776 33000
rect 30282 32988 30288 33000
rect 30340 33028 30346 33040
rect 31938 33028 31944 33040
rect 30340 33000 31944 33028
rect 30340 32988 30346 33000
rect 31938 32988 31944 33000
rect 31996 32988 32002 33040
rect 32416 33028 32444 33068
rect 32493 33065 32505 33099
rect 32539 33096 32551 33099
rect 33042 33096 33048 33108
rect 32539 33068 33048 33096
rect 32539 33065 32551 33068
rect 32493 33059 32551 33065
rect 33042 33056 33048 33068
rect 33100 33056 33106 33108
rect 37826 33096 37832 33108
rect 35866 33068 37832 33096
rect 35866 33028 35894 33068
rect 37826 33056 37832 33068
rect 37884 33096 37890 33108
rect 38197 33099 38255 33105
rect 38197 33096 38209 33099
rect 37884 33068 38209 33096
rect 37884 33056 37890 33068
rect 38197 33065 38209 33068
rect 38243 33065 38255 33099
rect 38197 33059 38255 33065
rect 32416 33000 35894 33028
rect 32582 32960 32588 32972
rect 30116 32932 32588 32960
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29826 32895 29884 32901
rect 29826 32861 29838 32895
rect 29872 32892 29884 32895
rect 29914 32892 29920 32904
rect 29872 32864 29920 32892
rect 29872 32861 29884 32864
rect 29826 32855 29884 32861
rect 26108 32796 27844 32824
rect 26108 32784 26114 32796
rect 28810 32784 28816 32836
rect 28868 32824 28874 32836
rect 28905 32827 28963 32833
rect 28905 32824 28917 32827
rect 28868 32796 28917 32824
rect 28868 32784 28874 32796
rect 28905 32793 28917 32796
rect 28951 32793 28963 32827
rect 28905 32787 28963 32793
rect 23624 32728 25452 32756
rect 23624 32716 23630 32728
rect 26142 32716 26148 32768
rect 26200 32756 26206 32768
rect 26237 32759 26295 32765
rect 26237 32756 26249 32759
rect 26200 32728 26249 32756
rect 26200 32716 26206 32728
rect 26237 32725 26249 32728
rect 26283 32725 26295 32759
rect 26237 32719 26295 32725
rect 26602 32716 26608 32768
rect 26660 32756 26666 32768
rect 29840 32756 29868 32855
rect 29914 32852 29920 32864
rect 29972 32852 29978 32904
rect 30116 32901 30144 32932
rect 30282 32901 30288 32904
rect 30101 32895 30159 32901
rect 30101 32861 30113 32895
rect 30147 32861 30159 32895
rect 30101 32855 30159 32861
rect 30239 32895 30288 32901
rect 30239 32861 30251 32895
rect 30285 32861 30288 32895
rect 30239 32855 30288 32861
rect 30282 32852 30288 32855
rect 30340 32892 30346 32904
rect 30975 32895 31033 32901
rect 30975 32892 30987 32895
rect 30340 32864 30987 32892
rect 30340 32852 30346 32864
rect 30975 32861 30987 32864
rect 31021 32861 31033 32895
rect 30975 32855 31033 32861
rect 31294 32852 31300 32904
rect 31352 32901 31358 32904
rect 31352 32895 31391 32901
rect 31379 32861 31391 32895
rect 31352 32855 31391 32861
rect 31352 32852 31358 32855
rect 31478 32852 31484 32904
rect 31536 32852 31542 32904
rect 31956 32901 31984 32932
rect 32582 32920 32588 32932
rect 32640 32920 32646 32972
rect 31941 32895 31999 32901
rect 31941 32861 31953 32895
rect 31987 32861 31999 32895
rect 31941 32855 31999 32861
rect 32214 32852 32220 32904
rect 32272 32852 32278 32904
rect 32306 32852 32312 32904
rect 32364 32852 32370 32904
rect 35434 32852 35440 32904
rect 35492 32892 35498 32904
rect 35866 32901 35894 33000
rect 36354 32920 36360 32972
rect 36412 32960 36418 32972
rect 36817 32963 36875 32969
rect 36817 32960 36829 32963
rect 36412 32932 36829 32960
rect 36412 32920 36418 32932
rect 36817 32929 36829 32932
rect 36863 32929 36875 32963
rect 36817 32923 36875 32929
rect 35713 32895 35771 32901
rect 35713 32892 35725 32895
rect 35492 32864 35725 32892
rect 35492 32852 35498 32864
rect 35713 32861 35725 32864
rect 35759 32861 35771 32895
rect 35713 32855 35771 32861
rect 35851 32895 35909 32901
rect 35851 32861 35863 32895
rect 35897 32861 35909 32895
rect 35851 32855 35909 32861
rect 36078 32852 36084 32904
rect 36136 32852 36142 32904
rect 36262 32901 36268 32904
rect 36219 32895 36268 32901
rect 36219 32861 36231 32895
rect 36265 32861 36268 32895
rect 36219 32855 36268 32861
rect 36262 32852 36268 32855
rect 36320 32852 36326 32904
rect 37090 32901 37096 32904
rect 37084 32892 37096 32901
rect 37051 32864 37096 32892
rect 37084 32855 37096 32864
rect 37090 32852 37096 32855
rect 37148 32852 37154 32904
rect 30006 32784 30012 32836
rect 30064 32784 30070 32836
rect 31110 32784 31116 32836
rect 31168 32784 31174 32836
rect 31205 32827 31263 32833
rect 31205 32793 31217 32827
rect 31251 32793 31263 32827
rect 31205 32787 31263 32793
rect 26660 32728 29868 32756
rect 30024 32756 30052 32784
rect 31220 32756 31248 32787
rect 31662 32784 31668 32836
rect 31720 32824 31726 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 31720 32796 32137 32824
rect 31720 32784 31726 32796
rect 32125 32793 32137 32796
rect 32171 32793 32183 32827
rect 32125 32787 32183 32793
rect 30024 32728 31248 32756
rect 26660 32716 26666 32728
rect 31754 32716 31760 32768
rect 31812 32756 31818 32768
rect 32232 32756 32260 32852
rect 35989 32827 36047 32833
rect 35989 32824 36001 32827
rect 35912 32796 36001 32824
rect 35912 32768 35940 32796
rect 35989 32793 36001 32796
rect 36035 32793 36047 32827
rect 35989 32787 36047 32793
rect 31812 32728 32260 32756
rect 31812 32716 31818 32728
rect 35802 32716 35808 32768
rect 35860 32756 35866 32768
rect 35894 32756 35900 32768
rect 35860 32728 35900 32756
rect 35860 32716 35866 32728
rect 35894 32716 35900 32728
rect 35952 32716 35958 32768
rect 36357 32759 36415 32765
rect 36357 32725 36369 32759
rect 36403 32756 36415 32759
rect 37918 32756 37924 32768
rect 36403 32728 37924 32756
rect 36403 32725 36415 32728
rect 36357 32719 36415 32725
rect 37918 32716 37924 32728
rect 37976 32716 37982 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 12437 32555 12495 32561
rect 12437 32521 12449 32555
rect 12483 32552 12495 32555
rect 13722 32552 13728 32564
rect 12483 32524 13728 32552
rect 12483 32521 12495 32524
rect 12437 32515 12495 32521
rect 13722 32512 13728 32524
rect 13780 32512 13786 32564
rect 14366 32552 14372 32564
rect 13832 32524 14372 32552
rect 6917 32487 6975 32493
rect 6917 32484 6929 32487
rect 6012 32456 6929 32484
rect 4522 32376 4528 32428
rect 4580 32376 4586 32428
rect 4617 32419 4675 32425
rect 4617 32385 4629 32419
rect 4663 32385 4675 32419
rect 4617 32379 4675 32385
rect 4632 32348 4660 32379
rect 4982 32376 4988 32428
rect 5040 32416 5046 32428
rect 5261 32419 5319 32425
rect 5261 32416 5273 32419
rect 5040 32388 5273 32416
rect 5040 32376 5046 32388
rect 5261 32385 5273 32388
rect 5307 32385 5319 32419
rect 5261 32379 5319 32385
rect 5810 32376 5816 32428
rect 5868 32416 5874 32428
rect 6012 32425 6040 32456
rect 6917 32453 6929 32456
rect 6963 32453 6975 32487
rect 6917 32447 6975 32453
rect 8021 32487 8079 32493
rect 8021 32453 8033 32487
rect 8067 32484 8079 32487
rect 9122 32484 9128 32496
rect 8067 32456 9128 32484
rect 8067 32453 8079 32456
rect 8021 32447 8079 32453
rect 9122 32444 9128 32456
rect 9180 32444 9186 32496
rect 9674 32444 9680 32496
rect 9732 32484 9738 32496
rect 10505 32487 10563 32493
rect 9732 32456 10364 32484
rect 9732 32444 9738 32456
rect 5997 32419 6055 32425
rect 5997 32416 6009 32419
rect 5868 32388 6009 32416
rect 5868 32376 5874 32388
rect 5997 32385 6009 32388
rect 6043 32385 6055 32419
rect 5997 32379 6055 32385
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32416 6883 32419
rect 7374 32416 7380 32428
rect 6871 32388 7380 32416
rect 6871 32385 6883 32388
rect 6825 32379 6883 32385
rect 6086 32348 6092 32360
rect 4632 32320 6092 32348
rect 6086 32308 6092 32320
rect 6144 32348 6150 32360
rect 6564 32348 6592 32379
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 8754 32376 8760 32428
rect 8812 32376 8818 32428
rect 9766 32376 9772 32428
rect 9824 32376 9830 32428
rect 9858 32376 9864 32428
rect 9916 32416 9922 32428
rect 9953 32419 10011 32425
rect 9953 32416 9965 32419
rect 9916 32388 9965 32416
rect 9916 32376 9922 32388
rect 9953 32385 9965 32388
rect 9999 32385 10011 32419
rect 9953 32379 10011 32385
rect 10134 32376 10140 32428
rect 10192 32376 10198 32428
rect 10336 32425 10364 32456
rect 10505 32453 10517 32487
rect 10551 32484 10563 32487
rect 12253 32487 12311 32493
rect 12253 32484 12265 32487
rect 10551 32456 12265 32484
rect 10551 32453 10563 32456
rect 10505 32447 10563 32453
rect 12253 32453 12265 32456
rect 12299 32453 12311 32487
rect 12253 32447 12311 32453
rect 13630 32444 13636 32496
rect 13688 32484 13694 32496
rect 13832 32484 13860 32524
rect 14366 32512 14372 32524
rect 14424 32512 14430 32564
rect 14458 32512 14464 32564
rect 14516 32552 14522 32564
rect 14737 32555 14795 32561
rect 14737 32552 14749 32555
rect 14516 32524 14749 32552
rect 14516 32512 14522 32524
rect 14737 32521 14749 32524
rect 14783 32521 14795 32555
rect 17586 32552 17592 32564
rect 14737 32515 14795 32521
rect 17144 32524 17592 32552
rect 13688 32456 13860 32484
rect 13688 32444 13694 32456
rect 14274 32444 14280 32496
rect 14332 32444 14338 32496
rect 17144 32484 17172 32524
rect 17586 32512 17592 32524
rect 17644 32512 17650 32564
rect 18322 32512 18328 32564
rect 18380 32552 18386 32564
rect 20898 32552 20904 32564
rect 18380 32524 20904 32552
rect 18380 32512 18386 32524
rect 20898 32512 20904 32524
rect 20956 32512 20962 32564
rect 23474 32512 23480 32564
rect 23532 32552 23538 32564
rect 24118 32552 24124 32564
rect 23532 32524 24124 32552
rect 23532 32512 23538 32524
rect 24118 32512 24124 32524
rect 24176 32512 24182 32564
rect 24504 32524 24808 32552
rect 20254 32484 20260 32496
rect 14476 32456 17172 32484
rect 17236 32456 20260 32484
rect 10321 32419 10379 32425
rect 10321 32385 10333 32419
rect 10367 32385 10379 32419
rect 10321 32379 10379 32385
rect 12066 32376 12072 32428
rect 12124 32376 12130 32428
rect 12158 32376 12164 32428
rect 12216 32376 12222 32428
rect 14476 32425 14504 32456
rect 14461 32419 14519 32425
rect 14461 32385 14473 32419
rect 14507 32385 14519 32419
rect 14461 32379 14519 32385
rect 14550 32376 14556 32428
rect 14608 32376 14614 32428
rect 14918 32376 14924 32428
rect 14976 32416 14982 32428
rect 15197 32419 15255 32425
rect 15197 32416 15209 32419
rect 14976 32388 15209 32416
rect 14976 32376 14982 32388
rect 15197 32385 15209 32388
rect 15243 32385 15255 32419
rect 15197 32379 15255 32385
rect 15378 32376 15384 32428
rect 15436 32376 15442 32428
rect 16298 32376 16304 32428
rect 16356 32376 16362 32428
rect 17236 32425 17264 32456
rect 20254 32444 20260 32456
rect 20312 32444 20318 32496
rect 21542 32444 21548 32496
rect 21600 32484 21606 32496
rect 24504 32484 24532 32524
rect 21600 32456 24532 32484
rect 24780 32484 24808 32524
rect 25222 32512 25228 32564
rect 25280 32552 25286 32564
rect 25869 32555 25927 32561
rect 25869 32552 25881 32555
rect 25280 32524 25881 32552
rect 25280 32512 25286 32524
rect 25869 32521 25881 32524
rect 25915 32552 25927 32555
rect 25915 32524 27384 32552
rect 25915 32521 25927 32524
rect 25869 32515 25927 32521
rect 24780 32456 26556 32484
rect 21600 32444 21606 32456
rect 16853 32419 16911 32425
rect 16853 32385 16865 32419
rect 16899 32385 16911 32419
rect 16853 32379 16911 32385
rect 17221 32419 17279 32425
rect 17221 32385 17233 32419
rect 17267 32385 17279 32419
rect 17221 32379 17279 32385
rect 6144 32320 6592 32348
rect 6144 32308 6150 32320
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 10045 32351 10103 32357
rect 10045 32348 10057 32351
rect 9732 32320 10057 32348
rect 9732 32308 9738 32320
rect 10045 32317 10057 32320
rect 10091 32317 10103 32351
rect 10045 32311 10103 32317
rect 11514 32308 11520 32360
rect 11572 32348 11578 32360
rect 15102 32348 15108 32360
rect 11572 32320 15108 32348
rect 11572 32308 11578 32320
rect 15102 32308 15108 32320
rect 15160 32308 15166 32360
rect 16868 32348 16896 32379
rect 17310 32376 17316 32428
rect 17368 32376 17374 32428
rect 20438 32376 20444 32428
rect 20496 32416 20502 32428
rect 22204 32425 22232 32456
rect 22189 32419 22247 32425
rect 20496 32388 22140 32416
rect 20496 32376 20502 32388
rect 17126 32348 17132 32360
rect 15304 32320 17132 32348
rect 5626 32240 5632 32292
rect 5684 32280 5690 32292
rect 7006 32280 7012 32292
rect 5684 32252 7012 32280
rect 5684 32240 5690 32252
rect 7006 32240 7012 32252
rect 7064 32240 7070 32292
rect 9306 32240 9312 32292
rect 9364 32280 9370 32292
rect 9364 32252 10732 32280
rect 9364 32240 9370 32252
rect 4801 32215 4859 32221
rect 4801 32181 4813 32215
rect 4847 32212 4859 32215
rect 4890 32212 4896 32224
rect 4847 32184 4896 32212
rect 4847 32181 4859 32184
rect 4801 32175 4859 32181
rect 4890 32172 4896 32184
rect 4948 32172 4954 32224
rect 5718 32172 5724 32224
rect 5776 32212 5782 32224
rect 5905 32215 5963 32221
rect 5905 32212 5917 32215
rect 5776 32184 5917 32212
rect 5776 32172 5782 32184
rect 5905 32181 5917 32184
rect 5951 32181 5963 32215
rect 5905 32175 5963 32181
rect 8018 32172 8024 32224
rect 8076 32212 8082 32224
rect 10594 32212 10600 32224
rect 8076 32184 10600 32212
rect 8076 32172 8082 32184
rect 10594 32172 10600 32184
rect 10652 32172 10658 32224
rect 10704 32212 10732 32252
rect 11882 32240 11888 32292
rect 11940 32240 11946 32292
rect 12986 32240 12992 32292
rect 13044 32280 13050 32292
rect 15304 32280 15332 32320
rect 17126 32308 17132 32320
rect 17184 32308 17190 32360
rect 20625 32351 20683 32357
rect 20625 32317 20637 32351
rect 20671 32348 20683 32351
rect 20714 32348 20720 32360
rect 20671 32320 20720 32348
rect 20671 32317 20683 32320
rect 20625 32311 20683 32317
rect 20714 32308 20720 32320
rect 20772 32348 20778 32360
rect 21910 32348 21916 32360
rect 20772 32320 21916 32348
rect 20772 32308 20778 32320
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 22112 32348 22140 32388
rect 22189 32385 22201 32419
rect 22235 32385 22247 32419
rect 22189 32379 22247 32385
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 22296 32348 22324 32379
rect 23474 32376 23480 32428
rect 23532 32376 23538 32428
rect 23842 32376 23848 32428
rect 23900 32376 23906 32428
rect 24394 32376 24400 32428
rect 24452 32376 24458 32428
rect 24486 32376 24492 32428
rect 24544 32376 24550 32428
rect 24670 32376 24676 32428
rect 24728 32376 24734 32428
rect 25777 32419 25835 32425
rect 25777 32416 25789 32419
rect 24780 32388 25789 32416
rect 24780 32348 24808 32388
rect 25777 32385 25789 32388
rect 25823 32416 25835 32419
rect 26050 32416 26056 32428
rect 25823 32388 26056 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26234 32376 26240 32428
rect 26292 32376 26298 32428
rect 22112 32320 24808 32348
rect 25133 32351 25191 32357
rect 25133 32317 25145 32351
rect 25179 32348 25191 32351
rect 25222 32348 25228 32360
rect 25179 32320 25228 32348
rect 25179 32317 25191 32320
rect 25133 32311 25191 32317
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 13044 32252 15332 32280
rect 13044 32240 13050 32252
rect 16022 32240 16028 32292
rect 16080 32280 16086 32292
rect 17497 32283 17555 32289
rect 17497 32280 17509 32283
rect 16080 32252 17509 32280
rect 16080 32240 16086 32252
rect 17497 32249 17509 32252
rect 17543 32249 17555 32283
rect 26528 32280 26556 32456
rect 27356 32416 27384 32524
rect 28718 32512 28724 32564
rect 28776 32561 28782 32564
rect 28776 32555 28789 32561
rect 28777 32552 28789 32555
rect 30745 32555 30803 32561
rect 28777 32524 28821 32552
rect 29932 32524 30696 32552
rect 28777 32521 28789 32524
rect 28776 32515 28789 32521
rect 28776 32512 28782 32515
rect 27617 32419 27675 32425
rect 27617 32416 27629 32419
rect 27356 32388 27629 32416
rect 27617 32385 27629 32388
rect 27663 32416 27675 32419
rect 27890 32416 27896 32428
rect 27663 32388 27896 32416
rect 27663 32385 27675 32388
rect 27617 32379 27675 32385
rect 27890 32376 27896 32388
rect 27948 32376 27954 32428
rect 27982 32376 27988 32428
rect 28040 32376 28046 32428
rect 28629 32419 28687 32425
rect 28629 32416 28641 32419
rect 28184 32388 28641 32416
rect 27706 32308 27712 32360
rect 27764 32348 27770 32360
rect 28184 32348 28212 32388
rect 28629 32385 28641 32388
rect 28675 32385 28687 32419
rect 28629 32379 28687 32385
rect 29730 32376 29736 32428
rect 29788 32416 29794 32428
rect 29932 32416 29960 32524
rect 30006 32444 30012 32496
rect 30064 32484 30070 32496
rect 30377 32487 30435 32493
rect 30377 32484 30389 32487
rect 30064 32456 30389 32484
rect 30064 32444 30070 32456
rect 30377 32453 30389 32456
rect 30423 32453 30435 32487
rect 30668 32484 30696 32524
rect 30745 32521 30757 32555
rect 30791 32552 30803 32555
rect 31018 32552 31024 32564
rect 30791 32524 31024 32552
rect 30791 32521 30803 32524
rect 30745 32515 30803 32521
rect 31018 32512 31024 32524
rect 31076 32512 31082 32564
rect 31662 32512 31668 32564
rect 31720 32552 31726 32564
rect 34514 32552 34520 32564
rect 31720 32524 34520 32552
rect 31720 32512 31726 32524
rect 34514 32512 34520 32524
rect 34572 32552 34578 32564
rect 34572 32524 35112 32552
rect 34572 32512 34578 32524
rect 30668 32456 31064 32484
rect 30377 32447 30435 32453
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 29788 32388 30113 32416
rect 29788 32376 29794 32388
rect 30101 32385 30113 32388
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 30194 32419 30252 32425
rect 30194 32385 30206 32419
rect 30240 32385 30252 32419
rect 30194 32379 30252 32385
rect 27764 32320 28212 32348
rect 27764 32308 27770 32320
rect 28258 32308 28264 32360
rect 28316 32348 28322 32360
rect 28316 32320 28382 32348
rect 28316 32308 28322 32320
rect 29454 32308 29460 32360
rect 29512 32348 29518 32360
rect 30208 32348 30236 32379
rect 30466 32376 30472 32428
rect 30524 32376 30530 32428
rect 30566 32419 30624 32425
rect 30566 32385 30578 32419
rect 30612 32385 30624 32419
rect 31036 32416 31064 32456
rect 31110 32444 31116 32496
rect 31168 32484 31174 32496
rect 35084 32493 35112 32524
rect 35434 32512 35440 32564
rect 35492 32512 35498 32564
rect 35069 32487 35127 32493
rect 31168 32456 34928 32484
rect 31168 32444 31174 32456
rect 31478 32416 31484 32428
rect 31036 32388 31484 32416
rect 30566 32379 30624 32385
rect 30282 32348 30288 32360
rect 29512 32320 30288 32348
rect 29512 32308 29518 32320
rect 30282 32308 30288 32320
rect 30340 32308 30346 32360
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 30576 32348 30604 32379
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 32858 32376 32864 32428
rect 32916 32416 32922 32428
rect 34900 32425 34928 32456
rect 35069 32453 35081 32487
rect 35115 32453 35127 32487
rect 35069 32447 35127 32453
rect 35161 32487 35219 32493
rect 35161 32453 35173 32487
rect 35207 32484 35219 32487
rect 35526 32484 35532 32496
rect 35207 32456 35532 32484
rect 35207 32453 35219 32456
rect 35161 32447 35219 32453
rect 35526 32444 35532 32456
rect 35584 32484 35590 32496
rect 35710 32484 35716 32496
rect 35584 32456 35716 32484
rect 35584 32444 35590 32456
rect 35710 32444 35716 32456
rect 35768 32444 35774 32496
rect 38102 32444 38108 32496
rect 38160 32444 38166 32496
rect 33025 32419 33083 32425
rect 33025 32416 33037 32419
rect 32916 32388 33037 32416
rect 32916 32376 32922 32388
rect 33025 32385 33037 32388
rect 33071 32385 33083 32419
rect 33025 32379 33083 32385
rect 34885 32419 34943 32425
rect 34885 32385 34897 32419
rect 34931 32385 34943 32419
rect 34885 32379 34943 32385
rect 30432 32320 30604 32348
rect 30432 32308 30438 32320
rect 31846 32308 31852 32360
rect 31904 32348 31910 32360
rect 32766 32348 32772 32360
rect 31904 32320 32772 32348
rect 31904 32308 31910 32320
rect 32766 32308 32772 32320
rect 32824 32308 32830 32360
rect 34900 32348 34928 32379
rect 35250 32376 35256 32428
rect 35308 32376 35314 32428
rect 37829 32419 37887 32425
rect 37829 32385 37841 32419
rect 37875 32416 37887 32419
rect 37918 32416 37924 32428
rect 37875 32388 37924 32416
rect 37875 32385 37887 32388
rect 37829 32379 37887 32385
rect 37918 32376 37924 32388
rect 37976 32376 37982 32428
rect 35618 32348 35624 32360
rect 34900 32320 35624 32348
rect 35618 32308 35624 32320
rect 35676 32308 35682 32360
rect 27982 32280 27988 32292
rect 26528 32252 27988 32280
rect 17497 32243 17555 32249
rect 27982 32240 27988 32252
rect 28040 32240 28046 32292
rect 31294 32280 31300 32292
rect 28368 32252 31300 32280
rect 28368 32224 28396 32252
rect 31294 32240 31300 32252
rect 31352 32240 31358 32292
rect 34698 32280 34704 32292
rect 34072 32252 34704 32280
rect 12434 32212 12440 32224
rect 10704 32184 12440 32212
rect 12434 32172 12440 32184
rect 12492 32212 12498 32224
rect 12710 32212 12716 32224
rect 12492 32184 12716 32212
rect 12492 32172 12498 32184
rect 12710 32172 12716 32184
rect 12768 32172 12774 32224
rect 13814 32172 13820 32224
rect 13872 32212 13878 32224
rect 14277 32215 14335 32221
rect 14277 32212 14289 32215
rect 13872 32184 14289 32212
rect 13872 32172 13878 32184
rect 14277 32181 14289 32184
rect 14323 32181 14335 32215
rect 14277 32175 14335 32181
rect 14366 32172 14372 32224
rect 14424 32212 14430 32224
rect 14918 32212 14924 32224
rect 14424 32184 14924 32212
rect 14424 32172 14430 32184
rect 14918 32172 14924 32184
rect 14976 32172 14982 32224
rect 15286 32172 15292 32224
rect 15344 32172 15350 32224
rect 15565 32215 15623 32221
rect 15565 32181 15577 32215
rect 15611 32212 15623 32215
rect 15930 32212 15936 32224
rect 15611 32184 15936 32212
rect 15611 32181 15623 32184
rect 15565 32175 15623 32181
rect 15930 32172 15936 32184
rect 15988 32172 15994 32224
rect 16114 32172 16120 32224
rect 16172 32172 16178 32224
rect 16942 32172 16948 32224
rect 17000 32212 17006 32224
rect 17402 32212 17408 32224
rect 17000 32184 17408 32212
rect 17000 32172 17006 32184
rect 17402 32172 17408 32184
rect 17460 32172 17466 32224
rect 20257 32215 20315 32221
rect 20257 32181 20269 32215
rect 20303 32212 20315 32215
rect 20438 32212 20444 32224
rect 20303 32184 20444 32212
rect 20303 32181 20315 32184
rect 20257 32175 20315 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 20806 32172 20812 32224
rect 20864 32212 20870 32224
rect 21450 32212 21456 32224
rect 20864 32184 21456 32212
rect 20864 32172 20870 32184
rect 21450 32172 21456 32184
rect 21508 32172 21514 32224
rect 22278 32172 22284 32224
rect 22336 32172 22342 32224
rect 23842 32172 23848 32224
rect 23900 32172 23906 32224
rect 25130 32172 25136 32224
rect 25188 32212 25194 32224
rect 28166 32212 28172 32224
rect 25188 32184 28172 32212
rect 25188 32172 25194 32184
rect 28166 32172 28172 32184
rect 28224 32172 28230 32224
rect 28350 32172 28356 32224
rect 28408 32172 28414 32224
rect 28810 32172 28816 32224
rect 28868 32212 28874 32224
rect 32306 32212 32312 32224
rect 28868 32184 32312 32212
rect 28868 32172 28874 32184
rect 32306 32172 32312 32184
rect 32364 32212 32370 32224
rect 34072 32212 34100 32252
rect 34698 32240 34704 32252
rect 34756 32280 34762 32292
rect 35250 32280 35256 32292
rect 34756 32252 35256 32280
rect 34756 32240 34762 32252
rect 35250 32240 35256 32252
rect 35308 32240 35314 32292
rect 32364 32184 34100 32212
rect 32364 32172 32370 32184
rect 34146 32172 34152 32224
rect 34204 32172 34210 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 5718 31968 5724 32020
rect 5776 32008 5782 32020
rect 8018 32008 8024 32020
rect 5776 31980 8024 32008
rect 5776 31968 5782 31980
rect 3418 31900 3424 31952
rect 3476 31940 3482 31952
rect 3476 31912 5396 31940
rect 3476 31900 3482 31912
rect 5368 31881 5396 31912
rect 6822 31900 6828 31952
rect 6880 31900 6886 31952
rect 6932 31949 6960 31980
rect 8018 31968 8024 31980
rect 8076 31968 8082 32020
rect 9309 32011 9367 32017
rect 9309 31977 9321 32011
rect 9355 32008 9367 32011
rect 9674 32008 9680 32020
rect 9355 31980 9680 32008
rect 9355 31977 9367 31980
rect 9309 31971 9367 31977
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 9766 31968 9772 32020
rect 9824 32008 9830 32020
rect 9953 32011 10011 32017
rect 9953 32008 9965 32011
rect 9824 31980 9965 32008
rect 9824 31968 9830 31980
rect 9953 31977 9965 31980
rect 9999 31977 10011 32011
rect 9953 31971 10011 31977
rect 10318 31968 10324 32020
rect 10376 32008 10382 32020
rect 10413 32011 10471 32017
rect 10413 32008 10425 32011
rect 10376 31980 10425 32008
rect 10376 31968 10382 31980
rect 10413 31977 10425 31980
rect 10459 31977 10471 32011
rect 10413 31971 10471 31977
rect 12161 32011 12219 32017
rect 12161 31977 12173 32011
rect 12207 32008 12219 32011
rect 12207 31980 12434 32008
rect 12207 31977 12219 31980
rect 12161 31971 12219 31977
rect 6917 31943 6975 31949
rect 6917 31909 6929 31943
rect 6963 31940 6975 31943
rect 7193 31943 7251 31949
rect 6963 31912 6997 31940
rect 6963 31909 6975 31912
rect 6917 31903 6975 31909
rect 7193 31909 7205 31943
rect 7239 31940 7251 31943
rect 9582 31940 9588 31952
rect 7239 31912 9588 31940
rect 7239 31909 7251 31912
rect 7193 31903 7251 31909
rect 9582 31900 9588 31912
rect 9640 31900 9646 31952
rect 10781 31943 10839 31949
rect 10781 31909 10793 31943
rect 10827 31940 10839 31943
rect 11974 31940 11980 31952
rect 10827 31912 11980 31940
rect 10827 31909 10839 31912
rect 10781 31903 10839 31909
rect 11974 31900 11980 31912
rect 12032 31900 12038 31952
rect 12406 31940 12434 31980
rect 12710 31968 12716 32020
rect 12768 31968 12774 32020
rect 14734 32008 14740 32020
rect 12912 31980 14740 32008
rect 12912 31940 12940 31980
rect 14734 31968 14740 31980
rect 14792 31968 14798 32020
rect 14826 31968 14832 32020
rect 14884 31968 14890 32020
rect 15194 31968 15200 32020
rect 15252 31968 15258 32020
rect 15396 31980 15792 32008
rect 12406 31912 12940 31940
rect 12986 31900 12992 31952
rect 13044 31900 13050 31952
rect 13725 31943 13783 31949
rect 13725 31909 13737 31943
rect 13771 31940 13783 31943
rect 15396 31940 15424 31980
rect 13771 31912 15424 31940
rect 13771 31909 13783 31912
rect 13725 31903 13783 31909
rect 15562 31900 15568 31952
rect 15620 31940 15626 31952
rect 15657 31943 15715 31949
rect 15657 31940 15669 31943
rect 15620 31912 15669 31940
rect 15620 31900 15626 31912
rect 15657 31909 15669 31912
rect 15703 31909 15715 31943
rect 15764 31940 15792 31980
rect 15838 31968 15844 32020
rect 15896 31968 15902 32020
rect 17221 32011 17279 32017
rect 16592 31980 16804 32008
rect 16592 31940 16620 31980
rect 15764 31912 16620 31940
rect 16669 31943 16727 31949
rect 15657 31903 15715 31909
rect 16669 31909 16681 31943
rect 16715 31909 16727 31943
rect 16776 31940 16804 31980
rect 17221 31977 17233 32011
rect 17267 32008 17279 32011
rect 18046 32008 18052 32020
rect 17267 31980 18052 32008
rect 17267 31977 17279 31980
rect 17221 31971 17279 31977
rect 18046 31968 18052 31980
rect 18104 31968 18110 32020
rect 19613 32011 19671 32017
rect 19613 31977 19625 32011
rect 19659 32008 19671 32011
rect 22094 32008 22100 32020
rect 19659 31980 22100 32008
rect 19659 31977 19671 31980
rect 19613 31971 19671 31977
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 22554 31968 22560 32020
rect 22612 32008 22618 32020
rect 22830 32008 22836 32020
rect 22612 31980 22836 32008
rect 22612 31968 22618 31980
rect 22830 31968 22836 31980
rect 22888 31968 22894 32020
rect 23753 32011 23811 32017
rect 23753 31977 23765 32011
rect 23799 32008 23811 32011
rect 26694 32008 26700 32020
rect 23799 31980 26700 32008
rect 23799 31977 23811 31980
rect 23753 31971 23811 31977
rect 26694 31968 26700 31980
rect 26752 31968 26758 32020
rect 27816 31980 30236 32008
rect 16776 31912 18644 31940
rect 16669 31903 16727 31909
rect 5353 31875 5411 31881
rect 4172 31844 4936 31872
rect 4172 31813 4200 31844
rect 4908 31813 4936 31844
rect 5353 31841 5365 31875
rect 5399 31872 5411 31875
rect 6086 31872 6092 31884
rect 5399 31844 6092 31872
rect 5399 31841 5411 31844
rect 5353 31835 5411 31841
rect 6086 31832 6092 31844
rect 6144 31832 6150 31884
rect 6181 31875 6239 31881
rect 6181 31841 6193 31875
rect 6227 31872 6239 31875
rect 10318 31872 10324 31884
rect 6227 31844 7972 31872
rect 6227 31841 6239 31844
rect 6181 31835 6239 31841
rect 6932 31816 6960 31844
rect 4157 31807 4215 31813
rect 4157 31773 4169 31807
rect 4203 31773 4215 31807
rect 4157 31767 4215 31773
rect 4341 31807 4399 31813
rect 4341 31773 4353 31807
rect 4387 31804 4399 31807
rect 4801 31807 4859 31813
rect 4801 31804 4813 31807
rect 4387 31776 4813 31804
rect 4387 31773 4399 31776
rect 4341 31767 4399 31773
rect 4801 31773 4813 31776
rect 4847 31773 4859 31807
rect 4801 31767 4859 31773
rect 4893 31807 4951 31813
rect 4893 31773 4905 31807
rect 4939 31804 4951 31807
rect 5810 31804 5816 31816
rect 4939 31776 5816 31804
rect 4939 31773 4951 31776
rect 4893 31767 4951 31773
rect 4816 31736 4844 31767
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 6733 31807 6791 31813
rect 6733 31773 6745 31807
rect 6779 31773 6791 31807
rect 6733 31767 6791 31773
rect 4982 31736 4988 31748
rect 4816 31708 4988 31736
rect 4982 31696 4988 31708
rect 5040 31736 5046 31748
rect 5997 31739 6055 31745
rect 5997 31736 6009 31739
rect 5040 31708 6009 31736
rect 5040 31696 5046 31708
rect 5997 31705 6009 31708
rect 6043 31705 6055 31739
rect 6748 31736 6776 31767
rect 6914 31764 6920 31816
rect 6972 31764 6978 31816
rect 7006 31764 7012 31816
rect 7064 31804 7070 31816
rect 7944 31813 7972 31844
rect 8220 31844 10324 31872
rect 7929 31807 7987 31813
rect 7064 31776 7880 31804
rect 7064 31764 7070 31776
rect 7852 31736 7880 31776
rect 7929 31773 7941 31807
rect 7975 31773 7987 31807
rect 7929 31767 7987 31773
rect 8018 31764 8024 31816
rect 8076 31764 8082 31816
rect 8110 31764 8116 31816
rect 8168 31804 8174 31816
rect 8220 31813 8248 31844
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 11790 31872 11796 31884
rect 10428 31844 11796 31872
rect 8205 31807 8263 31813
rect 8205 31804 8217 31807
rect 8168 31776 8217 31804
rect 8168 31764 8174 31776
rect 8205 31773 8217 31776
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 8294 31764 8300 31816
rect 8352 31764 8358 31816
rect 9217 31807 9275 31813
rect 9217 31773 9229 31807
rect 9263 31804 9275 31807
rect 9306 31804 9312 31816
rect 9263 31776 9312 31804
rect 9263 31773 9275 31776
rect 9217 31767 9275 31773
rect 9306 31764 9312 31776
rect 9364 31764 9370 31816
rect 9490 31764 9496 31816
rect 9548 31764 9554 31816
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31773 9735 31807
rect 9677 31767 9735 31773
rect 8312 31736 8340 31764
rect 6748 31708 7052 31736
rect 7852 31708 8340 31736
rect 9692 31736 9720 31767
rect 9766 31764 9772 31816
rect 9824 31804 9830 31816
rect 10428 31813 10456 31844
rect 11790 31832 11796 31844
rect 11848 31872 11854 31884
rect 11848 31844 12020 31872
rect 11848 31832 11854 31844
rect 10413 31807 10471 31813
rect 10413 31804 10425 31807
rect 9824 31776 10425 31804
rect 9824 31764 9830 31776
rect 10413 31773 10425 31776
rect 10459 31773 10471 31807
rect 10413 31767 10471 31773
rect 10502 31764 10508 31816
rect 10560 31764 10566 31816
rect 11606 31764 11612 31816
rect 11664 31764 11670 31816
rect 11698 31764 11704 31816
rect 11756 31764 11762 31816
rect 11992 31813 12020 31844
rect 12066 31832 12072 31884
rect 12124 31872 12130 31884
rect 12124 31844 13492 31872
rect 12124 31832 12130 31844
rect 11885 31807 11943 31813
rect 11885 31773 11897 31807
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 11977 31807 12035 31813
rect 11977 31773 11989 31807
rect 12023 31773 12035 31807
rect 11977 31767 12035 31773
rect 10134 31736 10140 31748
rect 9692 31708 10140 31736
rect 5997 31699 6055 31705
rect 7024 31680 7052 31708
rect 10134 31696 10140 31708
rect 10192 31696 10198 31748
rect 4062 31628 4068 31680
rect 4120 31628 4126 31680
rect 7006 31628 7012 31680
rect 7064 31628 7070 31680
rect 7742 31628 7748 31680
rect 7800 31628 7806 31680
rect 9582 31628 9588 31680
rect 9640 31628 9646 31680
rect 11698 31628 11704 31680
rect 11756 31668 11762 31680
rect 11900 31668 11928 31767
rect 12342 31764 12348 31816
rect 12400 31804 12406 31816
rect 12621 31807 12679 31813
rect 12621 31804 12633 31807
rect 12400 31776 12633 31804
rect 12400 31764 12406 31776
rect 12621 31773 12633 31776
rect 12667 31773 12679 31807
rect 12621 31767 12679 31773
rect 12802 31764 12808 31816
rect 12860 31804 12866 31816
rect 13464 31813 13492 31844
rect 14550 31832 14556 31884
rect 14608 31872 14614 31884
rect 14826 31872 14832 31884
rect 14608 31844 14832 31872
rect 14608 31832 14614 31844
rect 14826 31832 14832 31844
rect 14884 31832 14890 31884
rect 15930 31872 15936 31884
rect 15028 31844 15936 31872
rect 15028 31813 15056 31844
rect 15930 31832 15936 31844
rect 15988 31832 15994 31884
rect 16684 31872 16712 31903
rect 16132 31844 16712 31872
rect 17037 31875 17095 31881
rect 13449 31807 13507 31813
rect 12860 31776 12940 31804
rect 12860 31764 12866 31776
rect 12912 31736 12940 31776
rect 13449 31773 13461 31807
rect 13495 31773 13507 31807
rect 13449 31767 13507 31773
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 15013 31807 15071 31813
rect 14783 31776 14964 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 13725 31739 13783 31745
rect 13725 31736 13737 31739
rect 12912 31708 13737 31736
rect 13725 31705 13737 31708
rect 13771 31705 13783 31739
rect 14936 31736 14964 31776
rect 15013 31773 15025 31807
rect 15059 31773 15071 31807
rect 15013 31767 15071 31773
rect 15120 31776 15976 31804
rect 15120 31736 15148 31776
rect 14936 31708 15148 31736
rect 15948 31736 15976 31776
rect 16022 31764 16028 31816
rect 16080 31764 16086 31816
rect 16132 31736 16160 31844
rect 17037 31841 17049 31875
rect 17083 31872 17095 31875
rect 17586 31872 17592 31884
rect 17083 31844 17592 31872
rect 17083 31841 17095 31844
rect 17037 31835 17095 31841
rect 17586 31832 17592 31844
rect 17644 31872 17650 31884
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17644 31844 18521 31872
rect 17644 31832 17650 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18616 31872 18644 31912
rect 18874 31900 18880 31952
rect 18932 31940 18938 31952
rect 18932 31912 19656 31940
rect 18932 31900 18938 31912
rect 19521 31875 19579 31881
rect 19521 31872 19533 31875
rect 18616 31844 19533 31872
rect 18509 31835 18567 31841
rect 19521 31841 19533 31844
rect 19567 31841 19579 31875
rect 19628 31872 19656 31912
rect 19794 31900 19800 31952
rect 19852 31900 19858 31952
rect 20346 31900 20352 31952
rect 20404 31940 20410 31952
rect 20530 31940 20536 31952
rect 20404 31912 20536 31940
rect 20404 31900 20410 31912
rect 20530 31900 20536 31912
rect 20588 31900 20594 31952
rect 21450 31900 21456 31952
rect 21508 31940 21514 31952
rect 22925 31943 22983 31949
rect 21508 31912 22876 31940
rect 21508 31900 21514 31912
rect 21266 31872 21272 31884
rect 19628 31844 21272 31872
rect 19521 31835 19579 31841
rect 16850 31764 16856 31816
rect 16908 31764 16914 31816
rect 17126 31764 17132 31816
rect 17184 31804 17190 31816
rect 17313 31807 17371 31813
rect 17313 31804 17325 31807
rect 17184 31776 17325 31804
rect 17184 31764 17190 31776
rect 17313 31773 17325 31776
rect 17359 31773 17371 31807
rect 17313 31767 17371 31773
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31804 18751 31807
rect 19334 31804 19340 31816
rect 18739 31776 19340 31804
rect 18739 31773 18751 31776
rect 18693 31767 18751 31773
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 21192 31813 21220 31844
rect 21266 31832 21272 31844
rect 21324 31832 21330 31884
rect 21545 31875 21603 31881
rect 21545 31841 21557 31875
rect 21591 31872 21603 31875
rect 22554 31872 22560 31884
rect 21591 31844 22560 31872
rect 21591 31841 21603 31844
rect 21545 31835 21603 31841
rect 22554 31832 22560 31844
rect 22612 31832 22618 31884
rect 22848 31881 22876 31912
rect 22925 31909 22937 31943
rect 22971 31940 22983 31943
rect 23106 31940 23112 31952
rect 22971 31912 23112 31940
rect 22971 31909 22983 31912
rect 22925 31903 22983 31909
rect 23106 31900 23112 31912
rect 23164 31900 23170 31952
rect 25682 31940 25688 31952
rect 23952 31912 25688 31940
rect 22833 31875 22891 31881
rect 22833 31841 22845 31875
rect 22879 31872 22891 31875
rect 23952 31872 23980 31912
rect 25682 31900 25688 31912
rect 25740 31900 25746 31952
rect 26142 31900 26148 31952
rect 26200 31940 26206 31952
rect 27816 31940 27844 31980
rect 29178 31940 29184 31952
rect 26200 31912 27844 31940
rect 27908 31912 29184 31940
rect 26200 31900 26206 31912
rect 27908 31884 27936 31912
rect 29178 31900 29184 31912
rect 29236 31900 29242 31952
rect 22879 31844 23980 31872
rect 22879 31841 22891 31844
rect 22833 31835 22891 31841
rect 24302 31832 24308 31884
rect 24360 31872 24366 31884
rect 24360 31844 24624 31872
rect 24360 31832 24366 31844
rect 21177 31807 21235 31813
rect 19536 31776 21036 31804
rect 15948 31708 16160 31736
rect 18877 31739 18935 31745
rect 13725 31699 13783 31705
rect 18877 31705 18889 31739
rect 18923 31736 18935 31739
rect 19536 31736 19564 31776
rect 18923 31708 19564 31736
rect 21008 31736 21036 31776
rect 21177 31773 21189 31807
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 21358 31764 21364 31816
rect 21416 31764 21422 31816
rect 22922 31764 22928 31816
rect 22980 31804 22986 31816
rect 22980 31776 23796 31804
rect 22980 31764 22986 31776
rect 22649 31739 22707 31745
rect 21008 31708 21312 31736
rect 18923 31705 18935 31708
rect 18877 31699 18935 31705
rect 11756 31640 11928 31668
rect 11756 31628 11762 31640
rect 13538 31628 13544 31680
rect 13596 31628 13602 31680
rect 15194 31628 15200 31680
rect 15252 31668 15258 31680
rect 15746 31668 15752 31680
rect 15252 31640 15752 31668
rect 15252 31628 15258 31640
rect 15746 31628 15752 31640
rect 15804 31668 15810 31680
rect 16114 31668 16120 31680
rect 15804 31640 16120 31668
rect 15804 31628 15810 31640
rect 16114 31628 16120 31640
rect 16172 31628 16178 31680
rect 18690 31628 18696 31680
rect 18748 31668 18754 31680
rect 20254 31668 20260 31680
rect 18748 31640 20260 31668
rect 18748 31628 18754 31640
rect 20254 31628 20260 31640
rect 20312 31628 20318 31680
rect 21174 31628 21180 31680
rect 21232 31628 21238 31680
rect 21284 31668 21312 31708
rect 22649 31705 22661 31739
rect 22695 31736 22707 31739
rect 23382 31736 23388 31748
rect 22695 31708 23388 31736
rect 22695 31705 22707 31708
rect 22649 31699 22707 31705
rect 23382 31696 23388 31708
rect 23440 31696 23446 31748
rect 23768 31736 23796 31776
rect 23842 31764 23848 31816
rect 23900 31804 23906 31816
rect 24486 31804 24492 31816
rect 23900 31776 24492 31804
rect 23900 31764 23906 31776
rect 24486 31764 24492 31776
rect 24544 31764 24550 31816
rect 24596 31813 24624 31844
rect 24780 31844 26234 31872
rect 24780 31813 24808 31844
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 25501 31807 25559 31813
rect 25501 31773 25513 31807
rect 25547 31804 25559 31807
rect 25682 31804 25688 31816
rect 25547 31776 25688 31804
rect 25547 31773 25559 31776
rect 25501 31767 25559 31773
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 25866 31764 25872 31816
rect 25924 31764 25930 31816
rect 24029 31739 24087 31745
rect 24029 31736 24041 31739
rect 23768 31708 24041 31736
rect 24029 31705 24041 31708
rect 24075 31736 24087 31739
rect 25038 31736 25044 31748
rect 24075 31708 25044 31736
rect 24075 31705 24087 31708
rect 24029 31699 24087 31705
rect 25038 31696 25044 31708
rect 25096 31696 25102 31748
rect 26206 31736 26234 31844
rect 27890 31832 27896 31884
rect 27948 31832 27954 31884
rect 28258 31832 28264 31884
rect 28316 31832 28322 31884
rect 29825 31875 29883 31881
rect 29825 31872 29837 31875
rect 28368 31844 29837 31872
rect 27154 31764 27160 31816
rect 27212 31764 27218 31816
rect 27246 31764 27252 31816
rect 27304 31764 27310 31816
rect 27982 31764 27988 31816
rect 28040 31764 28046 31816
rect 28368 31813 28396 31844
rect 29825 31841 29837 31844
rect 29871 31841 29883 31875
rect 30208 31872 30236 31980
rect 30282 31968 30288 32020
rect 30340 32008 30346 32020
rect 32769 32011 32827 32017
rect 30340 31980 32720 32008
rect 30340 31968 30346 31980
rect 32309 31943 32367 31949
rect 32309 31909 32321 31943
rect 32355 31909 32367 31943
rect 32309 31903 32367 31909
rect 30282 31872 30288 31884
rect 30208 31844 30288 31872
rect 29825 31835 29883 31841
rect 30282 31832 30288 31844
rect 30340 31832 30346 31884
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31773 28411 31807
rect 28353 31767 28411 31773
rect 28626 31764 28632 31816
rect 28684 31804 28690 31816
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 28684 31776 29745 31804
rect 28684 31764 28690 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29911 31807 29969 31813
rect 29911 31804 29923 31807
rect 29733 31767 29791 31773
rect 29840 31776 29923 31804
rect 26973 31739 27031 31745
rect 26973 31736 26985 31739
rect 26206 31708 26985 31736
rect 26973 31705 26985 31708
rect 27019 31736 27031 31739
rect 27062 31736 27068 31748
rect 27019 31708 27068 31736
rect 27019 31705 27031 31708
rect 26973 31699 27031 31705
rect 27062 31696 27068 31708
rect 27120 31736 27126 31748
rect 28644 31736 28672 31764
rect 27120 31708 28672 31736
rect 28997 31739 29055 31745
rect 27120 31696 27126 31708
rect 28997 31705 29009 31739
rect 29043 31705 29055 31739
rect 28997 31699 29055 31705
rect 22462 31668 22468 31680
rect 21284 31640 22468 31668
rect 22462 31628 22468 31640
rect 22520 31668 22526 31680
rect 24673 31671 24731 31677
rect 24673 31668 24685 31671
rect 22520 31640 24685 31668
rect 22520 31628 22526 31640
rect 24673 31637 24685 31640
rect 24719 31637 24731 31671
rect 29012 31668 29040 31699
rect 29362 31696 29368 31748
rect 29420 31736 29426 31748
rect 29840 31736 29868 31776
rect 29911 31773 29923 31776
rect 29957 31773 29969 31807
rect 29911 31767 29969 31773
rect 32030 31764 32036 31816
rect 32088 31764 32094 31816
rect 32324 31804 32352 31903
rect 32692 31872 32720 31980
rect 32769 31977 32781 32011
rect 32815 32008 32827 32011
rect 32858 32008 32864 32020
rect 32815 31980 32864 32008
rect 32815 31977 32827 31980
rect 32769 31971 32827 31977
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 36538 32008 36544 32020
rect 35360 31980 36544 32008
rect 35360 31872 35388 31980
rect 36538 31968 36544 31980
rect 36596 32008 36602 32020
rect 37737 32011 37795 32017
rect 37737 32008 37749 32011
rect 36596 31980 37749 32008
rect 36596 31968 36602 31980
rect 37737 31977 37749 31980
rect 37783 31977 37795 32011
rect 37737 31971 37795 31977
rect 35986 31872 35992 31884
rect 32692 31844 35388 31872
rect 32769 31807 32827 31813
rect 32769 31804 32781 31807
rect 32324 31776 32781 31804
rect 32769 31773 32781 31776
rect 32815 31773 32827 31807
rect 32769 31767 32827 31773
rect 32950 31764 32956 31816
rect 33008 31764 33014 31816
rect 35250 31764 35256 31816
rect 35308 31764 35314 31816
rect 35360 31813 35388 31844
rect 35544 31844 35992 31872
rect 35346 31807 35404 31813
rect 35346 31773 35358 31807
rect 35392 31773 35404 31807
rect 35346 31767 35404 31773
rect 35434 31764 35440 31816
rect 35492 31764 35498 31816
rect 35544 31813 35572 31844
rect 35986 31832 35992 31844
rect 36044 31832 36050 31884
rect 36354 31832 36360 31884
rect 36412 31832 36418 31884
rect 35529 31807 35587 31813
rect 35529 31773 35541 31807
rect 35575 31773 35587 31807
rect 35529 31767 35587 31773
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31773 35679 31807
rect 35621 31767 35679 31773
rect 35759 31807 35817 31813
rect 35759 31773 35771 31807
rect 35805 31804 35817 31807
rect 36262 31804 36268 31816
rect 35805 31776 36268 31804
rect 35805 31773 35817 31776
rect 35759 31767 35817 31773
rect 29420 31708 29868 31736
rect 29420 31696 29426 31708
rect 32214 31696 32220 31748
rect 32272 31736 32278 31748
rect 32309 31739 32367 31745
rect 32309 31736 32321 31739
rect 32272 31708 32321 31736
rect 32272 31696 32278 31708
rect 32309 31705 32321 31708
rect 32355 31705 32367 31739
rect 35452 31736 35480 31764
rect 35636 31736 35664 31767
rect 36262 31764 36268 31776
rect 36320 31764 36326 31816
rect 35452 31708 35664 31736
rect 36624 31739 36682 31745
rect 32309 31699 32367 31705
rect 36624 31705 36636 31739
rect 36670 31736 36682 31739
rect 36906 31736 36912 31748
rect 36670 31708 36912 31736
rect 36670 31705 36682 31708
rect 36624 31699 36682 31705
rect 36906 31696 36912 31708
rect 36964 31696 36970 31748
rect 31110 31668 31116 31680
rect 29012 31640 31116 31668
rect 24673 31631 24731 31637
rect 31110 31628 31116 31640
rect 31168 31668 31174 31680
rect 31570 31668 31576 31680
rect 31168 31640 31576 31668
rect 31168 31628 31174 31640
rect 31570 31628 31576 31640
rect 31628 31628 31634 31680
rect 32125 31671 32183 31677
rect 32125 31637 32137 31671
rect 32171 31668 32183 31671
rect 32398 31668 32404 31680
rect 32171 31640 32404 31668
rect 32171 31637 32183 31640
rect 32125 31631 32183 31637
rect 32398 31628 32404 31640
rect 32456 31628 32462 31680
rect 35894 31628 35900 31680
rect 35952 31628 35958 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 5994 31464 6000 31476
rect 5684 31436 6000 31464
rect 5684 31424 5690 31436
rect 5994 31424 6000 31436
rect 6052 31424 6058 31476
rect 6638 31424 6644 31476
rect 6696 31464 6702 31476
rect 6696 31436 8340 31464
rect 6696 31424 6702 31436
rect 5460 31368 6592 31396
rect 5460 31340 5488 31368
rect 6564 31340 6592 31368
rect 7374 31356 7380 31408
rect 7432 31356 7438 31408
rect 8202 31356 8208 31408
rect 8260 31356 8266 31408
rect 8312 31396 8340 31436
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 10229 31467 10287 31473
rect 10229 31464 10241 31467
rect 9732 31436 10241 31464
rect 9732 31424 9738 31436
rect 10229 31433 10241 31436
rect 10275 31464 10287 31467
rect 11606 31464 11612 31476
rect 10275 31436 11612 31464
rect 10275 31433 10287 31436
rect 10229 31427 10287 31433
rect 11606 31424 11612 31436
rect 11664 31464 11670 31476
rect 12253 31467 12311 31473
rect 11664 31436 12112 31464
rect 11664 31424 11670 31436
rect 8312 31368 10180 31396
rect 4801 31331 4859 31337
rect 4801 31297 4813 31331
rect 4847 31328 4859 31331
rect 4890 31328 4896 31340
rect 4847 31300 4896 31328
rect 4847 31297 4859 31300
rect 4801 31291 4859 31297
rect 4890 31288 4896 31300
rect 4948 31288 4954 31340
rect 4982 31288 4988 31340
rect 5040 31328 5046 31340
rect 5442 31328 5448 31340
rect 5040 31300 5448 31328
rect 5040 31288 5046 31300
rect 5442 31288 5448 31300
rect 5500 31288 5506 31340
rect 5810 31288 5816 31340
rect 5868 31288 5874 31340
rect 5997 31331 6055 31337
rect 5997 31297 6009 31331
rect 6043 31328 6055 31331
rect 6086 31328 6092 31340
rect 6043 31300 6092 31328
rect 6043 31297 6055 31300
rect 5997 31291 6055 31297
rect 6086 31288 6092 31300
rect 6144 31288 6150 31340
rect 6546 31288 6552 31340
rect 6604 31288 6610 31340
rect 6733 31331 6791 31337
rect 6733 31297 6745 31331
rect 6779 31328 6791 31331
rect 6822 31328 6828 31340
rect 6779 31300 6828 31328
rect 6779 31297 6791 31300
rect 6733 31291 6791 31297
rect 6822 31288 6828 31300
rect 6880 31288 6886 31340
rect 7190 31288 7196 31340
rect 7248 31328 7254 31340
rect 10152 31337 10180 31368
rect 11790 31356 11796 31408
rect 11848 31396 11854 31408
rect 12084 31405 12112 31436
rect 12253 31433 12265 31467
rect 12299 31464 12311 31467
rect 13538 31464 13544 31476
rect 12299 31436 13544 31464
rect 12299 31433 12311 31436
rect 12253 31427 12311 31433
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 18877 31467 18935 31473
rect 18877 31433 18889 31467
rect 18923 31464 18935 31467
rect 19426 31464 19432 31476
rect 18923 31436 19432 31464
rect 18923 31433 18935 31436
rect 18877 31427 18935 31433
rect 19426 31424 19432 31436
rect 19484 31424 19490 31476
rect 19610 31424 19616 31476
rect 19668 31464 19674 31476
rect 21174 31464 21180 31476
rect 19668 31436 21180 31464
rect 19668 31424 19674 31436
rect 21174 31424 21180 31436
rect 21232 31424 21238 31476
rect 22097 31467 22155 31473
rect 22097 31433 22109 31467
rect 22143 31433 22155 31467
rect 22097 31427 22155 31433
rect 11885 31399 11943 31405
rect 11885 31396 11897 31399
rect 11848 31368 11897 31396
rect 11848 31356 11854 31368
rect 11885 31365 11897 31368
rect 11931 31365 11943 31399
rect 11885 31359 11943 31365
rect 12069 31399 12127 31405
rect 12069 31365 12081 31399
rect 12115 31396 12127 31399
rect 12342 31396 12348 31408
rect 12115 31368 12348 31396
rect 12115 31365 12127 31368
rect 12069 31359 12127 31365
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 13354 31356 13360 31408
rect 13412 31396 13418 31408
rect 13449 31399 13507 31405
rect 13449 31396 13461 31399
rect 13412 31368 13461 31396
rect 13412 31356 13418 31368
rect 13449 31365 13461 31368
rect 13495 31365 13507 31399
rect 15381 31399 15439 31405
rect 15381 31396 15393 31399
rect 13449 31359 13507 31365
rect 13556 31368 15393 31396
rect 8849 31331 8907 31337
rect 8849 31328 8861 31331
rect 7248 31300 8861 31328
rect 7248 31288 7254 31300
rect 8849 31297 8861 31300
rect 8895 31328 8907 31331
rect 9953 31331 10011 31337
rect 8895 31300 9895 31328
rect 8895 31297 8907 31300
rect 8849 31291 8907 31297
rect 5534 31220 5540 31272
rect 5592 31260 5598 31272
rect 6641 31263 6699 31269
rect 6641 31260 6653 31263
rect 5592 31232 6653 31260
rect 5592 31220 5598 31232
rect 6641 31229 6653 31232
rect 6687 31229 6699 31263
rect 9033 31263 9091 31269
rect 9033 31260 9045 31263
rect 6641 31223 6699 31229
rect 6748 31232 9045 31260
rect 6748 31204 6776 31232
rect 9033 31229 9045 31232
rect 9079 31229 9091 31263
rect 9033 31223 9091 31229
rect 9125 31263 9183 31269
rect 9125 31229 9137 31263
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 6730 31152 6736 31204
rect 6788 31152 6794 31204
rect 7282 31152 7288 31204
rect 7340 31192 7346 31204
rect 9140 31192 9168 31223
rect 9306 31192 9312 31204
rect 7340 31164 9312 31192
rect 7340 31152 7346 31164
rect 9306 31152 9312 31164
rect 9364 31152 9370 31204
rect 5169 31127 5227 31133
rect 5169 31093 5181 31127
rect 5215 31124 5227 31127
rect 5626 31124 5632 31136
rect 5215 31096 5632 31124
rect 5215 31093 5227 31096
rect 5169 31087 5227 31093
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 5721 31127 5779 31133
rect 5721 31093 5733 31127
rect 5767 31124 5779 31127
rect 7190 31124 7196 31136
rect 5767 31096 7196 31124
rect 5767 31093 5779 31096
rect 5721 31087 5779 31093
rect 7190 31084 7196 31096
rect 7248 31084 7254 31136
rect 7834 31084 7840 31136
rect 7892 31124 7898 31136
rect 8665 31127 8723 31133
rect 8665 31124 8677 31127
rect 7892 31096 8677 31124
rect 7892 31084 7898 31096
rect 8665 31093 8677 31096
rect 8711 31093 8723 31127
rect 9867 31124 9895 31300
rect 9953 31297 9965 31331
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 10137 31331 10195 31337
rect 10137 31297 10149 31331
rect 10183 31328 10195 31331
rect 10226 31328 10232 31340
rect 10183 31300 10232 31328
rect 10183 31297 10195 31300
rect 10137 31291 10195 31297
rect 9968 31260 9996 31291
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 12250 31288 12256 31340
rect 12308 31328 12314 31340
rect 12713 31331 12771 31337
rect 12713 31328 12725 31331
rect 12308 31300 12725 31328
rect 12308 31288 12314 31300
rect 12713 31297 12725 31300
rect 12759 31297 12771 31331
rect 12713 31291 12771 31297
rect 12897 31331 12955 31337
rect 12897 31297 12909 31331
rect 12943 31328 12955 31331
rect 12986 31328 12992 31340
rect 12943 31300 12992 31328
rect 12943 31297 12955 31300
rect 12897 31291 12955 31297
rect 12986 31288 12992 31300
rect 13044 31328 13050 31340
rect 13556 31328 13584 31368
rect 15381 31365 15393 31368
rect 15427 31365 15439 31399
rect 15381 31359 15439 31365
rect 13044 31300 13584 31328
rect 13044 31288 13050 31300
rect 13630 31288 13636 31340
rect 13688 31328 13694 31340
rect 14274 31328 14280 31340
rect 13688 31300 14280 31328
rect 13688 31288 13694 31300
rect 14274 31288 14280 31300
rect 14332 31288 14338 31340
rect 15396 31328 15424 31359
rect 15746 31356 15752 31408
rect 15804 31356 15810 31408
rect 16850 31356 16856 31408
rect 16908 31396 16914 31408
rect 19628 31396 19656 31424
rect 16908 31368 19656 31396
rect 16908 31356 16914 31368
rect 15838 31328 15844 31340
rect 15396 31300 15844 31328
rect 15838 31288 15844 31300
rect 15896 31288 15902 31340
rect 16960 31337 16988 31368
rect 20254 31356 20260 31408
rect 20312 31396 20318 31408
rect 22112 31396 22140 31427
rect 23014 31424 23020 31476
rect 23072 31464 23078 31476
rect 23842 31464 23848 31476
rect 23072 31436 23848 31464
rect 23072 31424 23078 31436
rect 23842 31424 23848 31436
rect 23900 31424 23906 31476
rect 24762 31424 24768 31476
rect 24820 31464 24826 31476
rect 25041 31467 25099 31473
rect 25041 31464 25053 31467
rect 24820 31436 25053 31464
rect 24820 31424 24826 31436
rect 25041 31433 25053 31436
rect 25087 31433 25099 31467
rect 25041 31427 25099 31433
rect 25682 31424 25688 31476
rect 25740 31464 25746 31476
rect 25866 31464 25872 31476
rect 25740 31436 25872 31464
rect 25740 31424 25746 31436
rect 25866 31424 25872 31436
rect 25924 31424 25930 31476
rect 25958 31424 25964 31476
rect 26016 31464 26022 31476
rect 26016 31436 26188 31464
rect 26016 31424 26022 31436
rect 20312 31368 22140 31396
rect 23676 31368 24900 31396
rect 20312 31356 20318 31368
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 18138 31328 18144 31340
rect 16945 31291 17003 31297
rect 17236 31300 18144 31328
rect 10502 31260 10508 31272
rect 9968 31232 10508 31260
rect 10502 31220 10508 31232
rect 10560 31220 10566 31272
rect 13722 31220 13728 31272
rect 13780 31260 13786 31272
rect 17236 31260 17264 31300
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 18233 31331 18291 31337
rect 18233 31297 18245 31331
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 13780 31232 17264 31260
rect 13780 31220 13786 31232
rect 17310 31220 17316 31272
rect 17368 31220 17374 31272
rect 17405 31263 17463 31269
rect 17405 31229 17417 31263
rect 17451 31260 17463 31263
rect 17494 31260 17500 31272
rect 17451 31232 17500 31260
rect 17451 31229 17463 31232
rect 17405 31223 17463 31229
rect 17494 31220 17500 31232
rect 17552 31260 17558 31272
rect 17770 31260 17776 31272
rect 17552 31232 17776 31260
rect 17552 31220 17558 31232
rect 17770 31220 17776 31232
rect 17828 31220 17834 31272
rect 18248 31260 18276 31291
rect 18506 31288 18512 31340
rect 18564 31288 18570 31340
rect 18690 31288 18696 31340
rect 18748 31288 18754 31340
rect 19150 31288 19156 31340
rect 19208 31328 19214 31340
rect 19613 31331 19671 31337
rect 19613 31328 19625 31331
rect 19208 31300 19625 31328
rect 19208 31288 19214 31300
rect 19613 31297 19625 31300
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31328 19855 31331
rect 20162 31328 20168 31340
rect 19843 31300 20168 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 21266 31288 21272 31340
rect 21324 31288 21330 31340
rect 21453 31331 21511 31337
rect 21453 31297 21465 31331
rect 21499 31328 21511 31331
rect 22097 31331 22155 31337
rect 22097 31328 22109 31331
rect 21499 31300 22109 31328
rect 21499 31297 21511 31300
rect 21453 31291 21511 31297
rect 22097 31297 22109 31300
rect 22143 31328 22155 31331
rect 22278 31328 22284 31340
rect 22143 31300 22284 31328
rect 22143 31297 22155 31300
rect 22097 31291 22155 31297
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22370 31288 22376 31340
rect 22428 31328 22434 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22428 31300 22477 31328
rect 22428 31288 22434 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 23382 31288 23388 31340
rect 23440 31288 23446 31340
rect 23676 31337 23704 31368
rect 24872 31340 24900 31368
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31297 23719 31331
rect 23661 31291 23719 31297
rect 24486 31288 24492 31340
rect 24544 31328 24550 31340
rect 24581 31331 24639 31337
rect 24581 31328 24593 31331
rect 24544 31300 24593 31328
rect 24544 31288 24550 31300
rect 24581 31297 24593 31300
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 24854 31288 24860 31340
rect 24912 31328 24918 31340
rect 25682 31328 25688 31340
rect 24912 31300 25688 31328
rect 24912 31288 24918 31300
rect 25682 31288 25688 31300
rect 25740 31288 25746 31340
rect 26160 31337 26188 31436
rect 28258 31424 28264 31476
rect 28316 31464 28322 31476
rect 28445 31467 28503 31473
rect 28445 31464 28457 31467
rect 28316 31436 28457 31464
rect 28316 31424 28322 31436
rect 28445 31433 28457 31436
rect 28491 31433 28503 31467
rect 28445 31427 28503 31433
rect 31297 31467 31355 31473
rect 31297 31433 31309 31467
rect 31343 31464 31355 31467
rect 32214 31464 32220 31476
rect 31343 31436 32220 31464
rect 31343 31433 31355 31436
rect 31297 31427 31355 31433
rect 28460 31396 28488 31427
rect 32214 31424 32220 31436
rect 32272 31464 32278 31476
rect 32493 31467 32551 31473
rect 32493 31464 32505 31467
rect 32272 31436 32505 31464
rect 32272 31424 32278 31436
rect 32493 31433 32505 31436
rect 32539 31433 32551 31467
rect 32493 31427 32551 31433
rect 32677 31467 32735 31473
rect 32677 31433 32689 31467
rect 32723 31464 32735 31467
rect 32950 31464 32956 31476
rect 32723 31436 32956 31464
rect 32723 31433 32735 31436
rect 32677 31427 32735 31433
rect 32950 31424 32956 31436
rect 33008 31424 33014 31476
rect 34885 31467 34943 31473
rect 34885 31433 34897 31467
rect 34931 31464 34943 31467
rect 35250 31464 35256 31476
rect 34931 31436 35256 31464
rect 34931 31433 34943 31436
rect 34885 31427 34943 31433
rect 35250 31424 35256 31436
rect 35308 31424 35314 31476
rect 36538 31424 36544 31476
rect 36596 31424 36602 31476
rect 36906 31424 36912 31476
rect 36964 31424 36970 31476
rect 28460 31368 29408 31396
rect 26053 31331 26111 31337
rect 26048 31297 26065 31331
rect 26099 31297 26111 31331
rect 26048 31291 26111 31297
rect 26145 31331 26203 31337
rect 26145 31297 26157 31331
rect 26191 31297 26203 31331
rect 26145 31291 26203 31297
rect 19429 31263 19487 31269
rect 19429 31260 19441 31263
rect 18248 31232 19441 31260
rect 19429 31229 19441 31232
rect 19475 31229 19487 31263
rect 19429 31223 19487 31229
rect 19705 31263 19763 31269
rect 19705 31229 19717 31263
rect 19751 31229 19763 31263
rect 19705 31223 19763 31229
rect 19889 31263 19947 31269
rect 19889 31229 19901 31263
rect 19935 31260 19947 31263
rect 20254 31260 20260 31272
rect 19935 31232 20260 31260
rect 19935 31229 19947 31232
rect 19889 31223 19947 31229
rect 16666 31152 16672 31204
rect 16724 31192 16730 31204
rect 19720 31192 19748 31223
rect 20254 31220 20260 31232
rect 20312 31260 20318 31272
rect 20806 31260 20812 31272
rect 20312 31232 20812 31260
rect 20312 31220 20318 31232
rect 20806 31220 20812 31232
rect 20864 31220 20870 31272
rect 23474 31220 23480 31272
rect 23532 31260 23538 31272
rect 23532 31232 23612 31260
rect 23532 31220 23538 31232
rect 20346 31192 20352 31204
rect 16724 31164 18460 31192
rect 19720 31164 20352 31192
rect 16724 31152 16730 31164
rect 11790 31124 11796 31136
rect 9867 31096 11796 31124
rect 8665 31087 8723 31093
rect 11790 31084 11796 31096
rect 11848 31084 11854 31136
rect 12713 31127 12771 31133
rect 12713 31093 12725 31127
rect 12759 31124 12771 31127
rect 14182 31124 14188 31136
rect 12759 31096 14188 31124
rect 12759 31093 12771 31096
rect 12713 31087 12771 31093
rect 14182 31084 14188 31096
rect 14240 31084 14246 31136
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 16206 31124 16212 31136
rect 15344 31096 16212 31124
rect 15344 31084 15350 31096
rect 16206 31084 16212 31096
rect 16264 31084 16270 31136
rect 17770 31084 17776 31136
rect 17828 31124 17834 31136
rect 18325 31127 18383 31133
rect 18325 31124 18337 31127
rect 17828 31096 18337 31124
rect 17828 31084 17834 31096
rect 18325 31093 18337 31096
rect 18371 31093 18383 31127
rect 18432 31124 18460 31164
rect 20346 31152 20352 31164
rect 20404 31152 20410 31204
rect 23382 31192 23388 31204
rect 20456 31164 23388 31192
rect 20456 31124 20484 31164
rect 23382 31152 23388 31164
rect 23440 31152 23446 31204
rect 23584 31192 23612 31232
rect 23750 31220 23756 31272
rect 23808 31260 23814 31272
rect 23845 31263 23903 31269
rect 23845 31260 23857 31263
rect 23808 31232 23857 31260
rect 23808 31220 23814 31232
rect 23845 31229 23857 31232
rect 23891 31229 23903 31263
rect 23845 31223 23903 31229
rect 23934 31220 23940 31272
rect 23992 31260 23998 31272
rect 24394 31260 24400 31272
rect 23992 31232 24400 31260
rect 23992 31220 23998 31232
rect 24394 31220 24400 31232
rect 24452 31260 24458 31272
rect 26048 31260 26076 31291
rect 26234 31288 26240 31340
rect 26292 31288 26298 31340
rect 26326 31288 26332 31340
rect 26384 31328 26390 31340
rect 26421 31331 26479 31337
rect 26421 31328 26433 31331
rect 26384 31300 26433 31328
rect 26384 31288 26390 31300
rect 26421 31297 26433 31300
rect 26467 31297 26479 31331
rect 26421 31291 26479 31297
rect 26970 31288 26976 31340
rect 27028 31328 27034 31340
rect 27246 31328 27252 31340
rect 27028 31300 27252 31328
rect 27028 31288 27034 31300
rect 27246 31288 27252 31300
rect 27304 31288 27310 31340
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 27816 31260 27844 31291
rect 27982 31288 27988 31340
rect 28040 31328 28046 31340
rect 28353 31331 28411 31337
rect 28353 31328 28365 31331
rect 28040 31300 28365 31328
rect 28040 31288 28046 31300
rect 28353 31297 28365 31300
rect 28399 31297 28411 31331
rect 28353 31291 28411 31297
rect 28626 31288 28632 31340
rect 28684 31288 28690 31340
rect 29178 31288 29184 31340
rect 29236 31288 29242 31340
rect 29380 31337 29408 31368
rect 30926 31356 30932 31408
rect 30984 31356 30990 31408
rect 31021 31399 31079 31405
rect 31021 31365 31033 31399
rect 31067 31396 31079 31399
rect 31202 31396 31208 31408
rect 31067 31368 31208 31396
rect 31067 31365 31079 31368
rect 31021 31359 31079 31365
rect 31202 31356 31208 31368
rect 31260 31356 31266 31408
rect 32306 31356 32312 31408
rect 32364 31356 32370 31408
rect 38102 31356 38108 31408
rect 38160 31356 38166 31408
rect 29365 31331 29423 31337
rect 29365 31297 29377 31331
rect 29411 31297 29423 31331
rect 29365 31291 29423 31297
rect 30650 31288 30656 31340
rect 30708 31288 30714 31340
rect 30742 31288 30748 31340
rect 30800 31328 30806 31340
rect 30800 31300 30972 31328
rect 30800 31288 30806 31300
rect 28994 31260 29000 31272
rect 24452 31232 29000 31260
rect 24452 31220 24458 31232
rect 28994 31220 29000 31232
rect 29052 31220 29058 31272
rect 30944 31260 30972 31300
rect 31110 31288 31116 31340
rect 31168 31337 31174 31340
rect 31168 31328 31176 31337
rect 31168 31300 31213 31328
rect 31168 31291 31176 31300
rect 31168 31288 31174 31291
rect 34330 31288 34336 31340
rect 34388 31288 34394 31340
rect 34514 31288 34520 31340
rect 34572 31288 34578 31340
rect 34609 31331 34667 31337
rect 34609 31297 34621 31331
rect 34655 31297 34667 31331
rect 34609 31291 34667 31297
rect 34146 31260 34152 31272
rect 30944 31232 34152 31260
rect 34146 31220 34152 31232
rect 34204 31220 34210 31272
rect 24673 31195 24731 31201
rect 24673 31192 24685 31195
rect 23584 31164 24685 31192
rect 24673 31161 24685 31164
rect 24719 31161 24731 31195
rect 24673 31155 24731 31161
rect 31294 31152 31300 31204
rect 31352 31192 31358 31204
rect 34624 31192 34652 31291
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 35342 31328 35348 31340
rect 34756 31300 35348 31328
rect 34756 31288 34762 31300
rect 35342 31288 35348 31300
rect 35400 31288 35406 31340
rect 35894 31288 35900 31340
rect 35952 31328 35958 31340
rect 36449 31331 36507 31337
rect 36449 31328 36461 31331
rect 35952 31300 36461 31328
rect 35952 31288 35958 31300
rect 36449 31297 36461 31300
rect 36495 31328 36507 31331
rect 37829 31331 37887 31337
rect 37829 31328 37841 31331
rect 36495 31300 37841 31328
rect 36495 31297 36507 31300
rect 36449 31291 36507 31297
rect 37829 31297 37841 31300
rect 37875 31297 37887 31331
rect 37829 31291 37887 31297
rect 36357 31263 36415 31269
rect 36357 31229 36369 31263
rect 36403 31260 36415 31263
rect 38010 31260 38016 31272
rect 36403 31232 38016 31260
rect 36403 31229 36415 31232
rect 36357 31223 36415 31229
rect 38010 31220 38016 31232
rect 38068 31220 38074 31272
rect 31352 31164 34652 31192
rect 31352 31152 31358 31164
rect 18432 31096 20484 31124
rect 21453 31127 21511 31133
rect 18325 31087 18383 31093
rect 21453 31093 21465 31127
rect 21499 31124 21511 31127
rect 22554 31124 22560 31136
rect 21499 31096 22560 31124
rect 21499 31093 21511 31096
rect 21453 31087 21511 31093
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 22738 31084 22744 31136
rect 22796 31124 22802 31136
rect 25222 31124 25228 31136
rect 22796 31096 25228 31124
rect 22796 31084 22802 31096
rect 25222 31084 25228 31096
rect 25280 31084 25286 31136
rect 25774 31084 25780 31136
rect 25832 31084 25838 31136
rect 27798 31084 27804 31136
rect 27856 31124 27862 31136
rect 29181 31127 29239 31133
rect 29181 31124 29193 31127
rect 27856 31096 29193 31124
rect 27856 31084 27862 31096
rect 29181 31093 29193 31096
rect 29227 31093 29239 31127
rect 29181 31087 29239 31093
rect 32030 31084 32036 31136
rect 32088 31124 32094 31136
rect 32493 31127 32551 31133
rect 32493 31124 32505 31127
rect 32088 31096 32505 31124
rect 32088 31084 32094 31096
rect 32493 31093 32505 31096
rect 32539 31093 32551 31127
rect 32493 31087 32551 31093
rect 34146 31084 34152 31136
rect 34204 31124 34210 31136
rect 35986 31124 35992 31136
rect 34204 31096 35992 31124
rect 34204 31084 34210 31096
rect 35986 31084 35992 31096
rect 36044 31084 36050 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 5258 30880 5264 30932
rect 5316 30920 5322 30932
rect 6730 30920 6736 30932
rect 5316 30892 6736 30920
rect 5316 30880 5322 30892
rect 6730 30880 6736 30892
rect 6788 30880 6794 30932
rect 7006 30880 7012 30932
rect 7064 30880 7070 30932
rect 8205 30923 8263 30929
rect 8205 30889 8217 30923
rect 8251 30920 8263 30923
rect 11882 30920 11888 30932
rect 8251 30892 11888 30920
rect 8251 30889 8263 30892
rect 8205 30883 8263 30889
rect 11882 30880 11888 30892
rect 11940 30880 11946 30932
rect 12158 30880 12164 30932
rect 12216 30920 12222 30932
rect 12437 30923 12495 30929
rect 12437 30920 12449 30923
rect 12216 30892 12449 30920
rect 12216 30880 12222 30892
rect 12437 30889 12449 30892
rect 12483 30889 12495 30923
rect 12437 30883 12495 30889
rect 14550 30880 14556 30932
rect 14608 30880 14614 30932
rect 14642 30880 14648 30932
rect 14700 30920 14706 30932
rect 14737 30923 14795 30929
rect 14737 30920 14749 30923
rect 14700 30892 14749 30920
rect 14700 30880 14706 30892
rect 14737 30889 14749 30892
rect 14783 30889 14795 30923
rect 14737 30883 14795 30889
rect 18049 30923 18107 30929
rect 18049 30889 18061 30923
rect 18095 30920 18107 30923
rect 19518 30920 19524 30932
rect 18095 30892 19524 30920
rect 18095 30889 18107 30892
rect 18049 30883 18107 30889
rect 19518 30880 19524 30892
rect 19576 30880 19582 30932
rect 19889 30923 19947 30929
rect 19889 30889 19901 30923
rect 19935 30920 19947 30923
rect 19978 30920 19984 30932
rect 19935 30892 19984 30920
rect 19935 30889 19947 30892
rect 19889 30883 19947 30889
rect 19978 30880 19984 30892
rect 20036 30880 20042 30932
rect 20438 30880 20444 30932
rect 20496 30880 20502 30932
rect 20806 30880 20812 30932
rect 20864 30920 20870 30932
rect 21085 30923 21143 30929
rect 21085 30920 21097 30923
rect 20864 30892 21097 30920
rect 20864 30880 20870 30892
rect 21085 30889 21097 30892
rect 21131 30889 21143 30923
rect 21085 30883 21143 30889
rect 22094 30880 22100 30932
rect 22152 30920 22158 30932
rect 23290 30920 23296 30932
rect 22152 30892 23296 30920
rect 22152 30880 22158 30892
rect 23290 30880 23296 30892
rect 23348 30880 23354 30932
rect 24029 30923 24087 30929
rect 24029 30889 24041 30923
rect 24075 30920 24087 30923
rect 25133 30923 25191 30929
rect 25133 30920 25145 30923
rect 24075 30892 25145 30920
rect 24075 30889 24087 30892
rect 24029 30883 24087 30889
rect 25133 30889 25145 30892
rect 25179 30920 25191 30923
rect 25406 30920 25412 30932
rect 25179 30892 25412 30920
rect 25179 30889 25191 30892
rect 25133 30883 25191 30889
rect 25406 30880 25412 30892
rect 25464 30880 25470 30932
rect 25866 30880 25872 30932
rect 25924 30920 25930 30932
rect 25961 30923 26019 30929
rect 25961 30920 25973 30923
rect 25924 30892 25973 30920
rect 25924 30880 25930 30892
rect 25961 30889 25973 30892
rect 26007 30889 26019 30923
rect 25961 30883 26019 30889
rect 26326 30880 26332 30932
rect 26384 30880 26390 30932
rect 28445 30923 28503 30929
rect 28445 30889 28457 30923
rect 28491 30920 28503 30923
rect 29730 30920 29736 30932
rect 28491 30892 29736 30920
rect 28491 30889 28503 30892
rect 28445 30883 28503 30889
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 36722 30920 36728 30932
rect 30024 30892 36728 30920
rect 4798 30812 4804 30864
rect 4856 30852 4862 30864
rect 4893 30855 4951 30861
rect 4893 30852 4905 30855
rect 4856 30824 4905 30852
rect 4856 30812 4862 30824
rect 4893 30821 4905 30824
rect 4939 30852 4951 30855
rect 5810 30852 5816 30864
rect 4939 30824 5816 30852
rect 4939 30821 4951 30824
rect 4893 30815 4951 30821
rect 5810 30812 5816 30824
rect 5868 30812 5874 30864
rect 6089 30855 6147 30861
rect 6089 30821 6101 30855
rect 6135 30852 6147 30855
rect 6135 30824 7788 30852
rect 6135 30821 6147 30824
rect 6089 30815 6147 30821
rect 6454 30784 6460 30796
rect 5092 30756 6460 30784
rect 5092 30657 5120 30756
rect 6454 30744 6460 30756
rect 6512 30744 6518 30796
rect 6546 30744 6552 30796
rect 6604 30784 6610 30796
rect 6641 30787 6699 30793
rect 6641 30784 6653 30787
rect 6604 30756 6653 30784
rect 6604 30744 6610 30756
rect 6641 30753 6653 30756
rect 6687 30753 6699 30787
rect 7760 30784 7788 30824
rect 7834 30812 7840 30864
rect 7892 30812 7898 30864
rect 7929 30855 7987 30861
rect 7929 30821 7941 30855
rect 7975 30852 7987 30855
rect 8110 30852 8116 30864
rect 7975 30824 8116 30852
rect 7975 30821 7987 30824
rect 7929 30815 7987 30821
rect 8110 30812 8116 30824
rect 8168 30812 8174 30864
rect 9306 30812 9312 30864
rect 9364 30852 9370 30864
rect 9401 30855 9459 30861
rect 9401 30852 9413 30855
rect 9364 30824 9413 30852
rect 9364 30812 9370 30824
rect 9401 30821 9413 30824
rect 9447 30821 9459 30855
rect 9401 30815 9459 30821
rect 9582 30812 9588 30864
rect 9640 30852 9646 30864
rect 9640 30824 15700 30852
rect 9640 30812 9646 30824
rect 9674 30784 9680 30796
rect 7760 30756 9680 30784
rect 6641 30747 6699 30753
rect 9674 30744 9680 30756
rect 9732 30744 9738 30796
rect 11606 30744 11612 30796
rect 11664 30784 11670 30796
rect 11701 30787 11759 30793
rect 11701 30784 11713 30787
rect 11664 30756 11713 30784
rect 11664 30744 11670 30756
rect 11701 30753 11713 30756
rect 11747 30753 11759 30787
rect 13541 30787 13599 30793
rect 13541 30784 13553 30787
rect 11701 30747 11759 30753
rect 11992 30756 13553 30784
rect 11992 30728 12020 30756
rect 13541 30753 13553 30756
rect 13587 30753 13599 30787
rect 13541 30747 13599 30753
rect 13722 30744 13728 30796
rect 13780 30744 13786 30796
rect 14461 30787 14519 30793
rect 14461 30753 14473 30787
rect 14507 30784 14519 30787
rect 15470 30784 15476 30796
rect 14507 30756 15476 30784
rect 14507 30753 14519 30756
rect 14461 30747 14519 30753
rect 15470 30744 15476 30756
rect 15528 30744 15534 30796
rect 15672 30793 15700 30824
rect 15746 30812 15752 30864
rect 15804 30852 15810 30864
rect 19429 30855 19487 30861
rect 19429 30852 19441 30855
rect 15804 30824 19441 30852
rect 15804 30812 15810 30824
rect 19429 30821 19441 30824
rect 19475 30821 19487 30855
rect 25774 30852 25780 30864
rect 19429 30815 19487 30821
rect 19812 30824 25780 30852
rect 15657 30787 15715 30793
rect 15657 30753 15669 30787
rect 15703 30753 15715 30787
rect 15657 30747 15715 30753
rect 15948 30756 19196 30784
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30716 5779 30719
rect 5810 30716 5816 30728
rect 5767 30688 5816 30716
rect 5767 30685 5779 30688
rect 5721 30679 5779 30685
rect 5810 30676 5816 30688
rect 5868 30716 5874 30728
rect 6825 30719 6883 30725
rect 5868 30688 6684 30716
rect 5868 30676 5874 30688
rect 5077 30651 5135 30657
rect 5077 30617 5089 30651
rect 5123 30617 5135 30651
rect 5077 30611 5135 30617
rect 5258 30608 5264 30660
rect 5316 30608 5322 30660
rect 5902 30608 5908 30660
rect 5960 30608 5966 30660
rect 6546 30608 6552 30660
rect 6604 30608 6610 30660
rect 6656 30648 6684 30688
rect 6825 30685 6837 30719
rect 6871 30716 6883 30719
rect 7282 30716 7288 30728
rect 6871 30688 7288 30716
rect 6871 30685 6883 30688
rect 6825 30679 6883 30685
rect 7282 30676 7288 30688
rect 7340 30676 7346 30728
rect 7742 30676 7748 30728
rect 7800 30676 7806 30728
rect 7834 30676 7840 30728
rect 7892 30716 7898 30728
rect 8021 30719 8079 30725
rect 8021 30716 8033 30719
rect 7892 30688 8033 30716
rect 7892 30676 7898 30688
rect 8021 30685 8033 30688
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 9398 30676 9404 30728
rect 9456 30676 9462 30728
rect 10413 30719 10471 30725
rect 10413 30685 10425 30719
rect 10459 30716 10471 30719
rect 11054 30716 11060 30728
rect 10459 30688 11060 30716
rect 10459 30685 10471 30688
rect 10413 30679 10471 30685
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 11790 30676 11796 30728
rect 11848 30676 11854 30728
rect 11974 30676 11980 30728
rect 12032 30676 12038 30728
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30716 12219 30719
rect 12250 30716 12256 30728
rect 12207 30688 12256 30716
rect 12207 30685 12219 30688
rect 12161 30679 12219 30685
rect 7006 30648 7012 30660
rect 6656 30620 7012 30648
rect 7006 30608 7012 30620
rect 7064 30608 7070 30660
rect 11606 30608 11612 30660
rect 11664 30648 11670 30660
rect 12176 30648 12204 30679
rect 12250 30676 12256 30688
rect 12308 30676 12314 30728
rect 12986 30676 12992 30728
rect 13044 30716 13050 30728
rect 13449 30719 13507 30725
rect 13449 30716 13461 30719
rect 13044 30688 13461 30716
rect 13044 30676 13050 30688
rect 13449 30685 13461 30688
rect 13495 30685 13507 30719
rect 13449 30679 13507 30685
rect 14182 30676 14188 30728
rect 14240 30716 14246 30728
rect 14277 30719 14335 30725
rect 14277 30716 14289 30719
rect 14240 30688 14289 30716
rect 14240 30676 14246 30688
rect 14277 30685 14289 30688
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 14553 30719 14611 30725
rect 14553 30685 14565 30719
rect 14599 30716 14611 30719
rect 15102 30716 15108 30728
rect 14599 30688 15108 30716
rect 14599 30685 14611 30688
rect 14553 30679 14611 30685
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15381 30719 15439 30725
rect 15381 30685 15393 30719
rect 15427 30685 15439 30719
rect 15381 30679 15439 30685
rect 11664 30620 12204 30648
rect 11664 30608 11670 30620
rect 4982 30540 4988 30592
rect 5040 30580 5046 30592
rect 5276 30580 5304 30608
rect 5040 30552 5304 30580
rect 5040 30540 5046 30552
rect 5626 30540 5632 30592
rect 5684 30580 5690 30592
rect 7742 30580 7748 30592
rect 5684 30552 7748 30580
rect 5684 30540 5690 30552
rect 7742 30540 7748 30552
rect 7800 30540 7806 30592
rect 11974 30540 11980 30592
rect 12032 30580 12038 30592
rect 12069 30583 12127 30589
rect 12069 30580 12081 30583
rect 12032 30552 12081 30580
rect 12032 30540 12038 30552
rect 12069 30549 12081 30552
rect 12115 30549 12127 30583
rect 12069 30543 12127 30549
rect 13725 30583 13783 30589
rect 13725 30549 13737 30583
rect 13771 30580 13783 30583
rect 13814 30580 13820 30592
rect 13771 30552 13820 30580
rect 13771 30549 13783 30552
rect 13725 30543 13783 30549
rect 13814 30540 13820 30552
rect 13872 30580 13878 30592
rect 14734 30580 14740 30592
rect 13872 30552 14740 30580
rect 13872 30540 13878 30552
rect 14734 30540 14740 30552
rect 14792 30540 14798 30592
rect 15194 30540 15200 30592
rect 15252 30540 15258 30592
rect 15396 30580 15424 30679
rect 15562 30676 15568 30728
rect 15620 30676 15626 30728
rect 15749 30719 15807 30725
rect 15749 30685 15761 30719
rect 15795 30716 15807 30719
rect 15838 30716 15844 30728
rect 15795 30688 15844 30716
rect 15795 30685 15807 30688
rect 15749 30679 15807 30685
rect 15838 30676 15844 30688
rect 15896 30676 15902 30728
rect 15948 30725 15976 30756
rect 15933 30719 15991 30725
rect 15933 30685 15945 30719
rect 15979 30685 15991 30719
rect 15933 30679 15991 30685
rect 16298 30676 16304 30728
rect 16356 30716 16362 30728
rect 16485 30719 16543 30725
rect 16485 30716 16497 30719
rect 16356 30688 16497 30716
rect 16356 30676 16362 30688
rect 16485 30685 16497 30688
rect 16531 30685 16543 30719
rect 16485 30679 16543 30685
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30716 16911 30719
rect 17678 30716 17684 30728
rect 16899 30688 17684 30716
rect 16899 30685 16911 30688
rect 16853 30679 16911 30685
rect 17678 30676 17684 30688
rect 17736 30676 17742 30728
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 17773 30679 17831 30685
rect 17034 30608 17040 30660
rect 17092 30648 17098 30660
rect 17788 30648 17816 30679
rect 17862 30676 17868 30728
rect 17920 30676 17926 30728
rect 17092 30620 17816 30648
rect 17092 30608 17098 30620
rect 18046 30608 18052 30660
rect 18104 30648 18110 30660
rect 18598 30648 18604 30660
rect 18104 30620 18604 30648
rect 18104 30608 18110 30620
rect 18598 30608 18604 30620
rect 18656 30608 18662 30660
rect 19168 30648 19196 30756
rect 19334 30744 19340 30796
rect 19392 30784 19398 30796
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19392 30756 19717 30784
rect 19392 30744 19398 30756
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 19610 30676 19616 30728
rect 19668 30676 19674 30728
rect 19812 30648 19840 30824
rect 25774 30812 25780 30824
rect 25832 30812 25838 30864
rect 26234 30812 26240 30864
rect 26292 30852 26298 30864
rect 26789 30855 26847 30861
rect 26789 30852 26801 30855
rect 26292 30824 26801 30852
rect 26292 30812 26298 30824
rect 26789 30821 26801 30824
rect 26835 30852 26847 30855
rect 27522 30852 27528 30864
rect 26835 30824 27528 30852
rect 26835 30821 26847 30824
rect 26789 30815 26847 30821
rect 27522 30812 27528 30824
rect 27580 30812 27586 30864
rect 30024 30861 30052 30892
rect 36722 30880 36728 30892
rect 36780 30880 36786 30932
rect 30009 30855 30067 30861
rect 30009 30821 30021 30855
rect 30055 30821 30067 30855
rect 30009 30815 30067 30821
rect 31389 30855 31447 30861
rect 31389 30821 31401 30855
rect 31435 30852 31447 30855
rect 32030 30852 32036 30864
rect 31435 30824 32036 30852
rect 31435 30821 31447 30824
rect 31389 30815 31447 30821
rect 32030 30812 32036 30824
rect 32088 30852 32094 30864
rect 32088 30824 32260 30852
rect 32088 30812 32094 30824
rect 20438 30744 20444 30796
rect 20496 30784 20502 30796
rect 20625 30787 20683 30793
rect 20625 30784 20637 30787
rect 20496 30756 20637 30784
rect 20496 30744 20502 30756
rect 20625 30753 20637 30756
rect 20671 30753 20683 30787
rect 22738 30784 22744 30796
rect 20625 30747 20683 30753
rect 22480 30756 22744 30784
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30716 20407 30719
rect 20530 30716 20536 30728
rect 20395 30688 20536 30716
rect 20395 30685 20407 30688
rect 20349 30679 20407 30685
rect 20530 30676 20536 30688
rect 20588 30676 20594 30728
rect 21082 30676 21088 30728
rect 21140 30676 21146 30728
rect 21266 30676 21272 30728
rect 21324 30716 21330 30728
rect 22480 30725 22508 30756
rect 22738 30744 22744 30756
rect 22796 30744 22802 30796
rect 25041 30787 25099 30793
rect 25041 30784 25053 30787
rect 23584 30756 25053 30784
rect 23584 30728 23612 30756
rect 25041 30753 25053 30756
rect 25087 30753 25099 30787
rect 25041 30747 25099 30753
rect 25130 30744 25136 30796
rect 25188 30784 25194 30796
rect 25188 30756 26004 30784
rect 25188 30744 25194 30756
rect 22465 30719 22523 30725
rect 22465 30716 22477 30719
rect 21324 30688 22477 30716
rect 21324 30676 21330 30688
rect 22465 30685 22477 30688
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 22646 30676 22652 30728
rect 22704 30676 22710 30728
rect 23382 30676 23388 30728
rect 23440 30716 23446 30728
rect 23566 30716 23572 30728
rect 23440 30688 23572 30716
rect 23440 30676 23446 30688
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 23842 30676 23848 30728
rect 23900 30676 23906 30728
rect 24029 30719 24087 30725
rect 24029 30685 24041 30719
rect 24075 30716 24087 30719
rect 24210 30716 24216 30728
rect 24075 30688 24216 30716
rect 24075 30685 24087 30688
rect 24029 30679 24087 30685
rect 24210 30676 24216 30688
rect 24268 30676 24274 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30685 25375 30719
rect 25317 30679 25375 30685
rect 19168 30620 19840 30648
rect 19889 30651 19947 30657
rect 19889 30617 19901 30651
rect 19935 30617 19947 30651
rect 19889 30611 19947 30617
rect 16298 30580 16304 30592
rect 15396 30552 16304 30580
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 17589 30583 17647 30589
rect 17589 30549 17601 30583
rect 17635 30580 17647 30583
rect 17862 30580 17868 30592
rect 17635 30552 17868 30580
rect 17635 30549 17647 30552
rect 17589 30543 17647 30549
rect 17862 30540 17868 30552
rect 17920 30540 17926 30592
rect 18138 30540 18144 30592
rect 18196 30580 18202 30592
rect 19426 30580 19432 30592
rect 18196 30552 19432 30580
rect 18196 30540 18202 30552
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 19904 30580 19932 30611
rect 22738 30608 22744 30660
rect 22796 30648 22802 30660
rect 25332 30648 25360 30679
rect 25498 30676 25504 30728
rect 25556 30716 25562 30728
rect 25774 30716 25780 30728
rect 25556 30688 25780 30716
rect 25556 30676 25562 30688
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 25976 30725 26004 30756
rect 31110 30744 31116 30796
rect 31168 30744 31174 30796
rect 32232 30793 32260 30824
rect 32217 30787 32275 30793
rect 32217 30753 32229 30787
rect 32263 30753 32275 30787
rect 32217 30747 32275 30753
rect 32677 30787 32735 30793
rect 32677 30753 32689 30787
rect 32723 30784 32735 30787
rect 33870 30784 33876 30796
rect 32723 30756 33876 30784
rect 32723 30753 32735 30756
rect 32677 30747 32735 30753
rect 33870 30744 33876 30756
rect 33928 30744 33934 30796
rect 25961 30719 26019 30725
rect 25961 30685 25973 30719
rect 26007 30685 26019 30719
rect 25961 30679 26019 30685
rect 26050 30676 26056 30728
rect 26108 30676 26114 30728
rect 27062 30676 27068 30728
rect 27120 30716 27126 30728
rect 27157 30719 27215 30725
rect 27157 30716 27169 30719
rect 27120 30688 27169 30716
rect 27120 30676 27126 30688
rect 27157 30685 27169 30688
rect 27203 30685 27215 30719
rect 27157 30679 27215 30685
rect 27522 30676 27528 30728
rect 27580 30716 27586 30728
rect 27617 30719 27675 30725
rect 27617 30716 27629 30719
rect 27580 30688 27629 30716
rect 27580 30676 27586 30688
rect 27617 30685 27629 30688
rect 27663 30685 27675 30719
rect 27617 30679 27675 30685
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30716 27859 30719
rect 28166 30716 28172 30728
rect 27847 30688 28172 30716
rect 27847 30685 27859 30688
rect 27801 30679 27859 30685
rect 28166 30676 28172 30688
rect 28224 30676 28230 30728
rect 28258 30676 28264 30728
rect 28316 30676 28322 30728
rect 28445 30719 28503 30725
rect 28445 30685 28457 30719
rect 28491 30716 28503 30719
rect 29178 30716 29184 30728
rect 28491 30688 29184 30716
rect 28491 30685 28503 30688
rect 28445 30679 28503 30685
rect 29178 30676 29184 30688
rect 29236 30676 29242 30728
rect 29822 30676 29828 30728
rect 29880 30676 29886 30728
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30685 29975 30719
rect 29917 30679 29975 30685
rect 22796 30620 25360 30648
rect 22796 30608 22802 30620
rect 26694 30608 26700 30660
rect 26752 30648 26758 30660
rect 26973 30651 27031 30657
rect 26973 30648 26985 30651
rect 26752 30620 26985 30648
rect 26752 30608 26758 30620
rect 26973 30617 26985 30620
rect 27019 30648 27031 30651
rect 27246 30648 27252 30660
rect 27019 30620 27252 30648
rect 27019 30617 27031 30620
rect 26973 30611 27031 30617
rect 27246 30608 27252 30620
rect 27304 30608 27310 30660
rect 29932 30648 29960 30679
rect 30742 30676 30748 30728
rect 30800 30676 30806 30728
rect 30838 30719 30896 30725
rect 30838 30685 30850 30719
rect 30884 30685 30896 30719
rect 30838 30679 30896 30685
rect 27448 30620 29960 30648
rect 20625 30583 20683 30589
rect 20625 30580 20637 30583
rect 19904 30552 20637 30580
rect 20625 30549 20637 30552
rect 20671 30580 20683 30583
rect 20898 30580 20904 30592
rect 20671 30552 20904 30580
rect 20671 30549 20683 30552
rect 20625 30543 20683 30549
rect 20898 30540 20904 30552
rect 20956 30540 20962 30592
rect 22830 30540 22836 30592
rect 22888 30540 22894 30592
rect 25501 30583 25559 30589
rect 25501 30549 25513 30583
rect 25547 30580 25559 30583
rect 27448 30580 27476 30620
rect 30466 30608 30472 30660
rect 30524 30648 30530 30660
rect 30852 30648 30880 30679
rect 30926 30676 30932 30728
rect 30984 30716 30990 30728
rect 31021 30719 31079 30725
rect 31021 30716 31033 30719
rect 30984 30688 31033 30716
rect 30984 30676 30990 30688
rect 31021 30685 31033 30688
rect 31067 30685 31079 30719
rect 31128 30716 31156 30744
rect 31210 30719 31268 30725
rect 31210 30716 31222 30719
rect 31128 30688 31222 30716
rect 31021 30679 31079 30685
rect 31210 30685 31222 30688
rect 31256 30716 31268 30719
rect 31478 30716 31484 30728
rect 31256 30688 31484 30716
rect 31256 30685 31268 30688
rect 31210 30679 31268 30685
rect 30524 30620 30880 30648
rect 30524 30608 30530 30620
rect 25547 30552 27476 30580
rect 25547 30549 25559 30552
rect 25501 30543 25559 30549
rect 27522 30540 27528 30592
rect 27580 30580 27586 30592
rect 27709 30583 27767 30589
rect 27709 30580 27721 30583
rect 27580 30552 27721 30580
rect 27580 30540 27586 30552
rect 27709 30549 27721 30552
rect 27755 30549 27767 30583
rect 27709 30543 27767 30549
rect 28629 30583 28687 30589
rect 28629 30549 28641 30583
rect 28675 30580 28687 30583
rect 28902 30580 28908 30592
rect 28675 30552 28908 30580
rect 28675 30549 28687 30552
rect 28629 30543 28687 30549
rect 28902 30540 28908 30552
rect 28960 30540 28966 30592
rect 31036 30580 31064 30679
rect 31478 30676 31484 30688
rect 31536 30676 31542 30728
rect 32306 30676 32312 30728
rect 32364 30676 32370 30728
rect 37826 30676 37832 30728
rect 37884 30676 37890 30728
rect 31110 30608 31116 30660
rect 31168 30608 31174 30660
rect 32324 30648 32352 30676
rect 32674 30648 32680 30660
rect 32324 30620 32680 30648
rect 32674 30608 32680 30620
rect 32732 30608 32738 30660
rect 38105 30651 38163 30657
rect 38105 30617 38117 30651
rect 38151 30648 38163 30651
rect 39022 30648 39028 30660
rect 38151 30620 39028 30648
rect 38151 30617 38163 30620
rect 38105 30611 38163 30617
rect 39022 30608 39028 30620
rect 39080 30608 39086 30660
rect 31294 30580 31300 30592
rect 31036 30552 31300 30580
rect 31294 30540 31300 30552
rect 31352 30540 31358 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 5902 30336 5908 30388
rect 5960 30376 5966 30388
rect 13173 30379 13231 30385
rect 5960 30348 9812 30376
rect 5960 30336 5966 30348
rect 7374 30308 7380 30320
rect 2792 30280 7380 30308
rect 2792 30252 2820 30280
rect 7374 30268 7380 30280
rect 7432 30308 7438 30320
rect 8386 30308 8392 30320
rect 7432 30280 8392 30308
rect 7432 30268 7438 30280
rect 8386 30268 8392 30280
rect 8444 30268 8450 30320
rect 9398 30308 9404 30320
rect 8588 30280 9404 30308
rect 2774 30200 2780 30252
rect 2832 30200 2838 30252
rect 3044 30243 3102 30249
rect 3044 30209 3056 30243
rect 3090 30240 3102 30243
rect 3970 30240 3976 30252
rect 3090 30212 3976 30240
rect 3090 30209 3102 30212
rect 3044 30203 3102 30209
rect 3970 30200 3976 30212
rect 4028 30200 4034 30252
rect 4798 30200 4804 30252
rect 4856 30200 4862 30252
rect 4985 30243 5043 30249
rect 4985 30209 4997 30243
rect 5031 30240 5043 30243
rect 5074 30240 5080 30252
rect 5031 30212 5080 30240
rect 5031 30209 5043 30212
rect 4985 30203 5043 30209
rect 5074 30200 5080 30212
rect 5132 30200 5138 30252
rect 5534 30200 5540 30252
rect 5592 30200 5598 30252
rect 5810 30200 5816 30252
rect 5868 30200 5874 30252
rect 6454 30200 6460 30252
rect 6512 30240 6518 30252
rect 7193 30243 7251 30249
rect 7193 30240 7205 30243
rect 6512 30212 7205 30240
rect 6512 30200 6518 30212
rect 7193 30209 7205 30212
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 4890 30132 4896 30184
rect 4948 30172 4954 30184
rect 5629 30175 5687 30181
rect 5629 30172 5641 30175
rect 4948 30144 5641 30172
rect 4948 30132 4954 30144
rect 5629 30141 5641 30144
rect 5675 30141 5687 30175
rect 5629 30135 5687 30141
rect 5721 30175 5779 30181
rect 5721 30141 5733 30175
rect 5767 30141 5779 30175
rect 7098 30172 7104 30184
rect 5721 30135 5779 30141
rect 6472 30144 7104 30172
rect 5736 30104 5764 30135
rect 6472 30104 6500 30144
rect 7098 30132 7104 30144
rect 7156 30132 7162 30184
rect 7208 30172 7236 30203
rect 7466 30200 7472 30252
rect 7524 30240 7530 30252
rect 8588 30249 8616 30280
rect 9398 30268 9404 30280
rect 9456 30268 9462 30320
rect 7745 30243 7803 30249
rect 7745 30240 7757 30243
rect 7524 30212 7757 30240
rect 7524 30200 7530 30212
rect 7745 30209 7757 30212
rect 7791 30240 7803 30243
rect 8573 30243 8631 30249
rect 7791 30212 8432 30240
rect 7791 30209 7803 30212
rect 7745 30203 7803 30209
rect 7650 30172 7656 30184
rect 7208 30144 7656 30172
rect 7650 30132 7656 30144
rect 7708 30132 7714 30184
rect 8404 30181 8432 30212
rect 8573 30209 8585 30243
rect 8619 30209 8631 30243
rect 8573 30203 8631 30209
rect 8754 30200 8760 30252
rect 8812 30240 8818 30252
rect 9030 30240 9036 30252
rect 8812 30212 9036 30240
rect 8812 30200 8818 30212
rect 9030 30200 9036 30212
rect 9088 30200 9094 30252
rect 9674 30200 9680 30252
rect 9732 30200 9738 30252
rect 9784 30240 9812 30348
rect 13173 30345 13185 30379
rect 13219 30376 13231 30379
rect 14366 30376 14372 30388
rect 13219 30348 14372 30376
rect 13219 30345 13231 30348
rect 13173 30339 13231 30345
rect 14366 30336 14372 30348
rect 14424 30336 14430 30388
rect 15562 30336 15568 30388
rect 15620 30376 15626 30388
rect 16117 30379 16175 30385
rect 16117 30376 16129 30379
rect 15620 30348 16129 30376
rect 15620 30336 15626 30348
rect 16117 30345 16129 30348
rect 16163 30345 16175 30379
rect 16117 30339 16175 30345
rect 18322 30336 18328 30388
rect 18380 30336 18386 30388
rect 20346 30336 20352 30388
rect 20404 30376 20410 30388
rect 24210 30376 24216 30388
rect 20404 30348 24216 30376
rect 20404 30336 20410 30348
rect 24210 30336 24216 30348
rect 24268 30376 24274 30388
rect 25958 30376 25964 30388
rect 24268 30348 25964 30376
rect 24268 30336 24274 30348
rect 9858 30268 9864 30320
rect 9916 30268 9922 30320
rect 10318 30268 10324 30320
rect 10376 30268 10382 30320
rect 10686 30308 10692 30320
rect 10520 30280 10692 30308
rect 10520 30249 10548 30280
rect 10686 30268 10692 30280
rect 10744 30308 10750 30320
rect 15105 30311 15163 30317
rect 10744 30280 11744 30308
rect 10744 30268 10750 30280
rect 11716 30249 11744 30280
rect 15105 30277 15117 30311
rect 15151 30308 15163 30311
rect 15746 30308 15752 30320
rect 15151 30280 15752 30308
rect 15151 30277 15163 30280
rect 15105 30271 15163 30277
rect 15746 30268 15752 30280
rect 15804 30268 15810 30320
rect 16482 30268 16488 30320
rect 16540 30308 16546 30320
rect 18138 30308 18144 30320
rect 16540 30280 18144 30308
rect 16540 30268 16546 30280
rect 18138 30268 18144 30280
rect 18196 30308 18202 30320
rect 18340 30308 18368 30336
rect 18196 30280 18368 30308
rect 18524 30280 24440 30308
rect 18196 30268 18202 30280
rect 10505 30243 10563 30249
rect 10505 30240 10517 30243
rect 9784 30212 10517 30240
rect 10505 30209 10517 30212
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 10597 30243 10655 30249
rect 10597 30209 10609 30243
rect 10643 30209 10655 30243
rect 10597 30203 10655 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 11701 30203 11759 30209
rect 8389 30175 8447 30181
rect 8389 30141 8401 30175
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9401 30175 9459 30181
rect 9401 30172 9413 30175
rect 9364 30144 9413 30172
rect 9364 30132 9370 30144
rect 9401 30141 9413 30144
rect 9447 30141 9459 30175
rect 10612 30172 10640 30203
rect 11790 30200 11796 30252
rect 11848 30200 11854 30252
rect 13081 30243 13139 30249
rect 13081 30240 13093 30243
rect 12406 30212 13093 30240
rect 9401 30135 9459 30141
rect 10520 30144 10640 30172
rect 5736 30076 6500 30104
rect 9416 30104 9444 30135
rect 10520 30116 10548 30144
rect 9416 30076 10364 30104
rect 4157 30039 4215 30045
rect 4157 30005 4169 30039
rect 4203 30036 4215 30039
rect 4614 30036 4620 30048
rect 4203 30008 4620 30036
rect 4203 30005 4215 30008
rect 4157 29999 4215 30005
rect 4614 29996 4620 30008
rect 4672 29996 4678 30048
rect 4798 29996 4804 30048
rect 4856 29996 4862 30048
rect 5994 29996 6000 30048
rect 6052 29996 6058 30048
rect 6086 29996 6092 30048
rect 6144 30036 6150 30048
rect 9030 30036 9036 30048
rect 6144 30008 9036 30036
rect 6144 29996 6150 30008
rect 9030 29996 9036 30008
rect 9088 30036 9094 30048
rect 10336 30045 10364 30076
rect 10502 30064 10508 30116
rect 10560 30064 10566 30116
rect 10781 30107 10839 30113
rect 10781 30073 10793 30107
rect 10827 30104 10839 30107
rect 11606 30104 11612 30116
rect 10827 30076 11612 30104
rect 10827 30073 10839 30076
rect 10781 30067 10839 30073
rect 11606 30064 11612 30076
rect 11664 30064 11670 30116
rect 11882 30064 11888 30116
rect 11940 30104 11946 30116
rect 12069 30107 12127 30113
rect 12069 30104 12081 30107
rect 11940 30076 12081 30104
rect 11940 30064 11946 30076
rect 12069 30073 12081 30076
rect 12115 30104 12127 30107
rect 12406 30104 12434 30212
rect 13081 30209 13093 30212
rect 13127 30209 13139 30243
rect 13081 30203 13139 30209
rect 13265 30243 13323 30249
rect 13265 30209 13277 30243
rect 13311 30209 13323 30243
rect 13265 30203 13323 30209
rect 14553 30243 14611 30249
rect 14553 30209 14565 30243
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 12986 30132 12992 30184
rect 13044 30172 13050 30184
rect 13280 30172 13308 30203
rect 13044 30144 13308 30172
rect 13044 30132 13050 30144
rect 12115 30076 12434 30104
rect 14568 30104 14596 30203
rect 15378 30200 15384 30252
rect 15436 30200 15442 30252
rect 16209 30243 16267 30249
rect 16209 30209 16221 30243
rect 16255 30240 16267 30243
rect 16666 30240 16672 30252
rect 16255 30212 16672 30240
rect 16255 30209 16267 30212
rect 16209 30203 16267 30209
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 17770 30200 17776 30252
rect 17828 30200 17834 30252
rect 17862 30200 17868 30252
rect 17920 30200 17926 30252
rect 18322 30200 18328 30252
rect 18380 30200 18386 30252
rect 18524 30249 18552 30280
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30209 18567 30243
rect 18509 30203 18567 30209
rect 20165 30243 20223 30249
rect 20165 30209 20177 30243
rect 20211 30240 20223 30243
rect 20254 30240 20260 30252
rect 20211 30212 20260 30240
rect 20211 30209 20223 30212
rect 20165 30203 20223 30209
rect 20254 30200 20260 30212
rect 20312 30200 20318 30252
rect 20346 30200 20352 30252
rect 20404 30200 20410 30252
rect 22649 30243 22707 30249
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 23198 30240 23204 30252
rect 22695 30212 23204 30240
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 23198 30200 23204 30212
rect 23256 30200 23262 30252
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30240 23443 30243
rect 23566 30240 23572 30252
rect 23431 30212 23572 30240
rect 23431 30209 23443 30212
rect 23385 30203 23443 30209
rect 23566 30200 23572 30212
rect 23624 30200 23630 30252
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 24029 30243 24087 30249
rect 24029 30209 24041 30243
rect 24075 30240 24087 30243
rect 24302 30240 24308 30252
rect 24075 30212 24308 30240
rect 24075 30209 24087 30212
rect 24029 30203 24087 30209
rect 14734 30132 14740 30184
rect 14792 30172 14798 30184
rect 15197 30175 15255 30181
rect 15197 30172 15209 30175
rect 14792 30144 15209 30172
rect 14792 30132 14798 30144
rect 15197 30141 15209 30144
rect 15243 30141 15255 30175
rect 15197 30135 15255 30141
rect 18598 30132 18604 30184
rect 18656 30172 18662 30184
rect 21450 30172 21456 30184
rect 18656 30144 21456 30172
rect 18656 30132 18662 30144
rect 21450 30132 21456 30144
rect 21508 30132 21514 30184
rect 23017 30175 23075 30181
rect 23017 30141 23029 30175
rect 23063 30172 23075 30175
rect 23290 30172 23296 30184
rect 23063 30144 23296 30172
rect 23063 30141 23075 30144
rect 23017 30135 23075 30141
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 15286 30104 15292 30116
rect 14568 30076 15292 30104
rect 12115 30073 12127 30076
rect 12069 30067 12127 30073
rect 15286 30064 15292 30076
rect 15344 30064 15350 30116
rect 15565 30107 15623 30113
rect 15565 30073 15577 30107
rect 15611 30104 15623 30107
rect 15654 30104 15660 30116
rect 15611 30076 15660 30104
rect 15611 30073 15623 30076
rect 15565 30067 15623 30073
rect 15654 30064 15660 30076
rect 15712 30064 15718 30116
rect 17402 30064 17408 30116
rect 17460 30104 17466 30116
rect 17497 30107 17555 30113
rect 17497 30104 17509 30107
rect 17460 30076 17509 30104
rect 17460 30064 17466 30076
rect 17497 30073 17509 30076
rect 17543 30073 17555 30107
rect 17497 30067 17555 30073
rect 17770 30064 17776 30116
rect 17828 30104 17834 30116
rect 22814 30107 22872 30113
rect 17828 30076 22508 30104
rect 17828 30064 17834 30076
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 9088 30008 9505 30036
rect 9088 29996 9094 30008
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 10321 30039 10379 30045
rect 10321 30005 10333 30039
rect 10367 30036 10379 30039
rect 11701 30039 11759 30045
rect 11701 30036 11713 30039
rect 10367 30008 11713 30036
rect 10367 30005 10379 30008
rect 10321 29999 10379 30005
rect 11701 30005 11713 30008
rect 11747 30036 11759 30039
rect 12526 30036 12532 30048
rect 11747 30008 12532 30036
rect 11747 30005 11759 30008
rect 11701 29999 11759 30005
rect 12526 29996 12532 30008
rect 12584 29996 12590 30048
rect 14458 29996 14464 30048
rect 14516 29996 14522 30048
rect 14550 29996 14556 30048
rect 14608 30036 14614 30048
rect 15105 30039 15163 30045
rect 15105 30036 15117 30039
rect 14608 30008 15117 30036
rect 14608 29996 14614 30008
rect 15105 30005 15117 30008
rect 15151 30005 15163 30039
rect 15105 29999 15163 30005
rect 17586 29996 17592 30048
rect 17644 30036 17650 30048
rect 17681 30039 17739 30045
rect 17681 30036 17693 30039
rect 17644 30008 17693 30036
rect 17644 29996 17650 30008
rect 17681 30005 17693 30008
rect 17727 30005 17739 30039
rect 17681 29999 17739 30005
rect 18506 29996 18512 30048
rect 18564 29996 18570 30048
rect 19981 30039 20039 30045
rect 19981 30005 19993 30039
rect 20027 30036 20039 30039
rect 20714 30036 20720 30048
rect 20027 30008 20720 30036
rect 20027 30005 20039 30008
rect 19981 29999 20039 30005
rect 20714 29996 20720 30008
rect 20772 29996 20778 30048
rect 22480 30036 22508 30076
rect 22814 30073 22826 30107
rect 22860 30104 22872 30107
rect 22860 30073 22876 30104
rect 22814 30067 22876 30073
rect 22646 30036 22652 30048
rect 22480 30008 22652 30036
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22848 30036 22876 30067
rect 22922 30064 22928 30116
rect 22980 30064 22986 30116
rect 23106 30036 23112 30048
rect 22848 30008 23112 30036
rect 23106 29996 23112 30008
rect 23164 29996 23170 30048
rect 23860 30036 23888 30203
rect 24302 30200 24308 30212
rect 24360 30200 24366 30252
rect 24412 30172 24440 30280
rect 24486 30268 24492 30320
rect 24544 30308 24550 30320
rect 24581 30311 24639 30317
rect 24581 30308 24593 30311
rect 24544 30280 24593 30308
rect 24544 30268 24550 30280
rect 24581 30277 24593 30280
rect 24627 30277 24639 30311
rect 24581 30271 24639 30277
rect 24688 30240 24716 30348
rect 25958 30336 25964 30348
rect 26016 30336 26022 30388
rect 27246 30336 27252 30388
rect 27304 30376 27310 30388
rect 27706 30376 27712 30388
rect 27304 30348 27712 30376
rect 27304 30336 27310 30348
rect 27706 30336 27712 30348
rect 27764 30376 27770 30388
rect 29362 30376 29368 30388
rect 27764 30348 29368 30376
rect 27764 30336 27770 30348
rect 29362 30336 29368 30348
rect 29420 30336 29426 30388
rect 30377 30379 30435 30385
rect 30377 30345 30389 30379
rect 30423 30376 30435 30379
rect 30650 30376 30656 30388
rect 30423 30348 30656 30376
rect 30423 30345 30435 30348
rect 30377 30339 30435 30345
rect 30650 30336 30656 30348
rect 30708 30336 30714 30388
rect 34977 30379 35035 30385
rect 33704 30348 34008 30376
rect 24765 30311 24823 30317
rect 24765 30277 24777 30311
rect 24811 30308 24823 30311
rect 25498 30308 25504 30320
rect 24811 30280 25504 30308
rect 24811 30277 24823 30280
rect 24765 30271 24823 30277
rect 25498 30268 25504 30280
rect 25556 30268 25562 30320
rect 27430 30268 27436 30320
rect 27488 30308 27494 30320
rect 27488 30280 29040 30308
rect 27488 30268 27494 30280
rect 24949 30243 25007 30249
rect 24949 30240 24961 30243
rect 24688 30212 24961 30240
rect 24949 30209 24961 30212
rect 24995 30209 25007 30243
rect 24949 30203 25007 30209
rect 25406 30200 25412 30252
rect 25464 30200 25470 30252
rect 25590 30200 25596 30252
rect 25648 30200 25654 30252
rect 25958 30200 25964 30252
rect 26016 30200 26022 30252
rect 27614 30200 27620 30252
rect 27672 30200 27678 30252
rect 29012 30249 29040 30280
rect 29086 30268 29092 30320
rect 29144 30268 29150 30320
rect 30006 30268 30012 30320
rect 30064 30268 30070 30320
rect 30466 30268 30472 30320
rect 30524 30308 30530 30320
rect 33704 30308 33732 30348
rect 33870 30317 33876 30320
rect 33864 30308 33876 30317
rect 30524 30280 33732 30308
rect 33831 30280 33876 30308
rect 30524 30268 30530 30280
rect 33864 30271 33876 30280
rect 33870 30268 33876 30271
rect 33928 30268 33934 30320
rect 33980 30308 34008 30348
rect 34977 30345 34989 30379
rect 35023 30345 35035 30379
rect 35894 30376 35900 30388
rect 34977 30339 35035 30345
rect 35728 30348 35900 30376
rect 34992 30308 35020 30339
rect 35728 30308 35756 30348
rect 35894 30336 35900 30348
rect 35952 30336 35958 30388
rect 37829 30311 37887 30317
rect 37829 30308 37841 30311
rect 33980 30280 35756 30308
rect 35820 30280 37841 30308
rect 28997 30243 29055 30249
rect 28997 30209 29009 30243
rect 29043 30209 29055 30243
rect 29104 30240 29132 30268
rect 29181 30243 29239 30249
rect 29181 30240 29193 30243
rect 29104 30212 29193 30240
rect 28997 30203 29055 30209
rect 29181 30209 29193 30212
rect 29227 30209 29239 30243
rect 29181 30203 29239 30209
rect 29730 30200 29736 30252
rect 29788 30200 29794 30252
rect 29826 30243 29884 30249
rect 29826 30209 29838 30243
rect 29872 30209 29884 30243
rect 29826 30203 29884 30209
rect 24762 30172 24768 30184
rect 24412 30144 24768 30172
rect 24762 30132 24768 30144
rect 24820 30172 24826 30184
rect 25314 30172 25320 30184
rect 24820 30144 25320 30172
rect 24820 30132 24826 30144
rect 25314 30132 25320 30144
rect 25372 30132 25378 30184
rect 26053 30175 26111 30181
rect 26053 30141 26065 30175
rect 26099 30172 26111 30175
rect 26142 30172 26148 30184
rect 26099 30144 26148 30172
rect 26099 30141 26111 30144
rect 26053 30135 26111 30141
rect 26142 30132 26148 30144
rect 26200 30132 26206 30184
rect 27430 30132 27436 30184
rect 27488 30172 27494 30184
rect 27893 30175 27951 30181
rect 27893 30172 27905 30175
rect 27488 30144 27905 30172
rect 27488 30132 27494 30144
rect 27893 30141 27905 30144
rect 27939 30141 27951 30175
rect 27893 30135 27951 30141
rect 29086 30132 29092 30184
rect 29144 30172 29150 30184
rect 29840 30172 29868 30203
rect 30098 30200 30104 30252
rect 30156 30200 30162 30252
rect 30282 30249 30288 30252
rect 30239 30243 30288 30249
rect 30239 30209 30251 30243
rect 30285 30209 30288 30243
rect 30239 30203 30288 30209
rect 30282 30200 30288 30203
rect 30340 30200 30346 30252
rect 32490 30200 32496 30252
rect 32548 30200 32554 30252
rect 32674 30200 32680 30252
rect 32732 30200 32738 30252
rect 33244 30212 35389 30240
rect 33244 30172 33272 30212
rect 29144 30144 33272 30172
rect 29144 30132 29150 30144
rect 33318 30132 33324 30184
rect 33376 30172 33382 30184
rect 33597 30175 33655 30181
rect 33597 30172 33609 30175
rect 33376 30144 33609 30172
rect 33376 30132 33382 30144
rect 33597 30141 33609 30144
rect 33643 30141 33655 30175
rect 35361 30172 35389 30212
rect 35434 30200 35440 30252
rect 35492 30240 35498 30252
rect 35621 30243 35679 30249
rect 35621 30240 35633 30243
rect 35492 30212 35633 30240
rect 35492 30200 35498 30212
rect 35621 30209 35633 30212
rect 35667 30209 35679 30243
rect 35621 30203 35679 30209
rect 35714 30243 35772 30249
rect 35714 30209 35726 30243
rect 35760 30240 35772 30243
rect 35820 30240 35848 30280
rect 37829 30277 37841 30280
rect 37875 30308 37887 30311
rect 38194 30308 38200 30320
rect 37875 30280 38200 30308
rect 37875 30277 37887 30280
rect 37829 30271 37887 30277
rect 38194 30268 38200 30280
rect 38252 30268 38258 30320
rect 35760 30212 35848 30240
rect 35897 30243 35955 30249
rect 35760 30209 35772 30212
rect 35714 30203 35772 30209
rect 35897 30209 35909 30243
rect 35943 30209 35955 30243
rect 35897 30203 35955 30209
rect 35728 30172 35756 30203
rect 35361 30144 35756 30172
rect 35912 30172 35940 30203
rect 35986 30200 35992 30252
rect 36044 30200 36050 30252
rect 36127 30243 36185 30249
rect 36127 30209 36139 30243
rect 36173 30240 36185 30243
rect 36262 30240 36268 30252
rect 36173 30212 36268 30240
rect 36173 30209 36185 30212
rect 36127 30203 36185 30209
rect 36262 30200 36268 30212
rect 36320 30200 36326 30252
rect 37921 30175 37979 30181
rect 35912 30144 36032 30172
rect 33597 30135 33655 30141
rect 24029 30107 24087 30113
rect 24029 30073 24041 30107
rect 24075 30104 24087 30107
rect 25406 30104 25412 30116
rect 24075 30076 25412 30104
rect 24075 30073 24087 30076
rect 24029 30067 24087 30073
rect 25406 30064 25412 30076
rect 25464 30064 25470 30116
rect 27448 30104 27476 30132
rect 36004 30116 36032 30144
rect 37921 30141 37933 30175
rect 37967 30141 37979 30175
rect 37921 30135 37979 30141
rect 25516 30076 27476 30104
rect 28920 30076 29868 30104
rect 25516 30036 25544 30076
rect 23860 30008 25544 30036
rect 26513 30039 26571 30045
rect 26513 30005 26525 30039
rect 26559 30036 26571 30039
rect 28920 30036 28948 30076
rect 26559 30008 28948 30036
rect 26559 30005 26571 30008
rect 26513 29999 26571 30005
rect 28994 29996 29000 30048
rect 29052 29996 29058 30048
rect 29840 30036 29868 30076
rect 30098 30064 30104 30116
rect 30156 30104 30162 30116
rect 33410 30104 33416 30116
rect 30156 30076 33416 30104
rect 30156 30064 30162 30076
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 35986 30064 35992 30116
rect 36044 30064 36050 30116
rect 36265 30107 36323 30113
rect 36265 30073 36277 30107
rect 36311 30104 36323 30107
rect 37826 30104 37832 30116
rect 36311 30076 37832 30104
rect 36311 30073 36323 30076
rect 36265 30067 36323 30073
rect 37826 30064 37832 30076
rect 37884 30104 37890 30116
rect 37936 30104 37964 30135
rect 38010 30132 38016 30184
rect 38068 30132 38074 30184
rect 37884 30076 37964 30104
rect 37884 30064 37890 30076
rect 31018 30036 31024 30048
rect 29840 30008 31024 30036
rect 31018 29996 31024 30008
rect 31076 29996 31082 30048
rect 32493 30039 32551 30045
rect 32493 30005 32505 30039
rect 32539 30036 32551 30039
rect 33134 30036 33140 30048
rect 32539 30008 33140 30036
rect 32539 30005 32551 30008
rect 32493 29999 32551 30005
rect 33134 29996 33140 30008
rect 33192 29996 33198 30048
rect 37458 29996 37464 30048
rect 37516 29996 37522 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 3970 29792 3976 29844
rect 4028 29792 4034 29844
rect 10134 29832 10140 29844
rect 4632 29804 10140 29832
rect 3418 29656 3424 29708
rect 3476 29656 3482 29708
rect 4632 29705 4660 29804
rect 10134 29792 10140 29804
rect 10192 29792 10198 29844
rect 11146 29792 11152 29844
rect 11204 29832 11210 29844
rect 11885 29835 11943 29841
rect 11885 29832 11897 29835
rect 11204 29804 11897 29832
rect 11204 29792 11210 29804
rect 11885 29801 11897 29804
rect 11931 29801 11943 29835
rect 11885 29795 11943 29801
rect 12066 29792 12072 29844
rect 12124 29792 12130 29844
rect 17218 29792 17224 29844
rect 17276 29792 17282 29844
rect 17405 29835 17463 29841
rect 17405 29801 17417 29835
rect 17451 29801 17463 29835
rect 17405 29795 17463 29801
rect 5994 29724 6000 29776
rect 6052 29764 6058 29776
rect 11517 29767 11575 29773
rect 11517 29764 11529 29767
rect 6052 29736 11529 29764
rect 6052 29724 6058 29736
rect 11517 29733 11529 29736
rect 11563 29764 11575 29767
rect 13814 29764 13820 29776
rect 11563 29736 13820 29764
rect 11563 29733 11575 29736
rect 11517 29727 11575 29733
rect 13814 29724 13820 29736
rect 13872 29724 13878 29776
rect 16206 29724 16212 29776
rect 16264 29764 16270 29776
rect 17420 29764 17448 29795
rect 19978 29792 19984 29844
rect 20036 29832 20042 29844
rect 20717 29835 20775 29841
rect 20717 29832 20729 29835
rect 20036 29804 20729 29832
rect 20036 29792 20042 29804
rect 20717 29801 20729 29804
rect 20763 29801 20775 29835
rect 20717 29795 20775 29801
rect 20824 29804 21680 29832
rect 16264 29736 17448 29764
rect 16264 29724 16270 29736
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 20824 29764 20852 29804
rect 21545 29767 21603 29773
rect 21545 29764 21557 29767
rect 17644 29736 20852 29764
rect 21100 29736 21557 29764
rect 17644 29724 17650 29736
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29665 4675 29699
rect 13262 29696 13268 29708
rect 4617 29659 4675 29665
rect 5552 29668 13268 29696
rect 3142 29588 3148 29640
rect 3200 29588 3206 29640
rect 3326 29588 3332 29640
rect 3384 29588 3390 29640
rect 5552 29628 5580 29668
rect 13262 29656 13268 29668
rect 13320 29656 13326 29708
rect 15470 29656 15476 29708
rect 15528 29696 15534 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 15528 29668 17509 29696
rect 15528 29656 15534 29668
rect 17497 29665 17509 29668
rect 17543 29696 17555 29699
rect 18506 29696 18512 29708
rect 17543 29668 18512 29696
rect 17543 29665 17555 29668
rect 17497 29659 17555 29665
rect 18506 29656 18512 29668
rect 18564 29656 18570 29708
rect 19426 29656 19432 29708
rect 19484 29696 19490 29708
rect 19484 29668 20484 29696
rect 19484 29656 19490 29668
rect 4816 29600 5580 29628
rect 2961 29563 3019 29569
rect 2961 29529 2973 29563
rect 3007 29560 3019 29563
rect 4433 29563 4491 29569
rect 4433 29560 4445 29563
rect 3007 29532 4445 29560
rect 3007 29529 3019 29532
rect 2961 29523 3019 29529
rect 4433 29529 4445 29532
rect 4479 29529 4491 29563
rect 4433 29523 4491 29529
rect 4341 29495 4399 29501
rect 4341 29461 4353 29495
rect 4387 29492 4399 29495
rect 4614 29492 4620 29504
rect 4387 29464 4620 29492
rect 4387 29461 4399 29464
rect 4341 29455 4399 29461
rect 4614 29452 4620 29464
rect 4672 29492 4678 29504
rect 4816 29492 4844 29600
rect 5626 29588 5632 29640
rect 5684 29628 5690 29640
rect 5997 29631 6055 29637
rect 5997 29628 6009 29631
rect 5684 29600 6009 29628
rect 5684 29588 5690 29600
rect 5997 29597 6009 29600
rect 6043 29597 6055 29631
rect 5997 29591 6055 29597
rect 7190 29588 7196 29640
rect 7248 29588 7254 29640
rect 7285 29631 7343 29637
rect 7285 29597 7297 29631
rect 7331 29597 7343 29631
rect 7285 29591 7343 29597
rect 5721 29563 5779 29569
rect 5721 29529 5733 29563
rect 5767 29560 5779 29563
rect 7300 29560 7328 29591
rect 7374 29588 7380 29640
rect 7432 29628 7438 29640
rect 7558 29628 7564 29640
rect 7432 29600 7564 29628
rect 7432 29588 7438 29600
rect 7558 29588 7564 29600
rect 7616 29588 7622 29640
rect 7650 29588 7656 29640
rect 7708 29628 7714 29640
rect 7745 29631 7803 29637
rect 7745 29628 7757 29631
rect 7708 29600 7757 29628
rect 7708 29588 7714 29600
rect 7745 29597 7757 29600
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 9309 29631 9367 29637
rect 9309 29597 9321 29631
rect 9355 29628 9367 29631
rect 9398 29628 9404 29640
rect 9355 29600 9404 29628
rect 9355 29597 9367 29600
rect 9309 29591 9367 29597
rect 9398 29588 9404 29600
rect 9456 29588 9462 29640
rect 14090 29588 14096 29640
rect 14148 29628 14154 29640
rect 15013 29631 15071 29637
rect 15013 29628 15025 29631
rect 14148 29600 15025 29628
rect 14148 29588 14154 29600
rect 15013 29597 15025 29600
rect 15059 29597 15071 29631
rect 15013 29591 15071 29597
rect 16482 29588 16488 29640
rect 16540 29588 16546 29640
rect 16669 29631 16727 29637
rect 16669 29597 16681 29631
rect 16715 29628 16727 29631
rect 16758 29628 16764 29640
rect 16715 29600 16764 29628
rect 16715 29597 16727 29600
rect 16669 29591 16727 29597
rect 16758 29588 16764 29600
rect 16816 29588 16822 29640
rect 17402 29588 17408 29640
rect 17460 29628 17466 29640
rect 17862 29628 17868 29640
rect 17460 29600 17868 29628
rect 17460 29588 17466 29600
rect 17862 29588 17868 29600
rect 17920 29588 17926 29640
rect 20254 29588 20260 29640
rect 20312 29628 20318 29640
rect 20456 29637 20484 29668
rect 20349 29631 20407 29637
rect 20349 29628 20361 29631
rect 20312 29600 20361 29628
rect 20312 29588 20318 29600
rect 20349 29597 20361 29600
rect 20395 29597 20407 29631
rect 20349 29591 20407 29597
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29597 20499 29631
rect 20441 29591 20499 29597
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 21100 29628 21128 29736
rect 21545 29733 21557 29736
rect 21591 29733 21603 29767
rect 21652 29764 21680 29804
rect 21726 29792 21732 29844
rect 21784 29832 21790 29844
rect 22281 29835 22339 29841
rect 22281 29832 22293 29835
rect 21784 29804 22293 29832
rect 21784 29792 21790 29804
rect 22281 29801 22293 29804
rect 22327 29801 22339 29835
rect 22281 29795 22339 29801
rect 22462 29792 22468 29844
rect 22520 29832 22526 29844
rect 22520 29804 22968 29832
rect 22520 29792 22526 29804
rect 22738 29764 22744 29776
rect 21652 29736 22744 29764
rect 21545 29727 21603 29733
rect 22738 29724 22744 29736
rect 22796 29724 22802 29776
rect 22833 29767 22891 29773
rect 22833 29733 22845 29767
rect 22879 29733 22891 29767
rect 22940 29764 22968 29804
rect 23014 29792 23020 29844
rect 23072 29832 23078 29844
rect 23290 29832 23296 29844
rect 23072 29804 23296 29832
rect 23072 29792 23078 29804
rect 23290 29792 23296 29804
rect 23348 29792 23354 29844
rect 23382 29792 23388 29844
rect 23440 29792 23446 29844
rect 25774 29792 25780 29844
rect 25832 29832 25838 29844
rect 26053 29835 26111 29841
rect 26053 29832 26065 29835
rect 25832 29804 26065 29832
rect 25832 29792 25838 29804
rect 26053 29801 26065 29804
rect 26099 29801 26111 29835
rect 26053 29795 26111 29801
rect 28610 29835 28668 29841
rect 28610 29801 28622 29835
rect 28656 29832 28668 29835
rect 28994 29832 29000 29844
rect 28656 29804 29000 29832
rect 28656 29801 28668 29804
rect 28610 29795 28668 29801
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 30377 29835 30435 29841
rect 30377 29801 30389 29835
rect 30423 29832 30435 29835
rect 30742 29832 30748 29844
rect 30423 29804 30748 29832
rect 30423 29801 30435 29804
rect 30377 29795 30435 29801
rect 30742 29792 30748 29804
rect 30800 29792 30806 29844
rect 31018 29792 31024 29844
rect 31076 29832 31082 29844
rect 31662 29832 31668 29844
rect 31076 29804 31668 29832
rect 31076 29792 31082 29804
rect 31662 29792 31668 29804
rect 31720 29792 31726 29844
rect 32125 29835 32183 29841
rect 32125 29801 32137 29835
rect 32171 29832 32183 29835
rect 32490 29832 32496 29844
rect 32171 29804 32496 29832
rect 32171 29801 32183 29804
rect 32125 29795 32183 29801
rect 32490 29792 32496 29804
rect 32548 29792 32554 29844
rect 34241 29835 34299 29841
rect 34241 29832 34253 29835
rect 32876 29804 34253 29832
rect 24026 29764 24032 29776
rect 22940 29736 24032 29764
rect 22833 29727 22891 29733
rect 21453 29699 21511 29705
rect 21453 29665 21465 29699
rect 21499 29665 21511 29699
rect 21453 29659 21511 29665
rect 20855 29600 21128 29628
rect 21468 29628 21496 29659
rect 21634 29656 21640 29708
rect 21692 29656 21698 29708
rect 22848 29696 22876 29727
rect 24026 29724 24032 29736
rect 24084 29724 24090 29776
rect 26237 29767 26295 29773
rect 26237 29733 26249 29767
rect 26283 29764 26295 29767
rect 26418 29764 26424 29776
rect 26283 29736 26424 29764
rect 26283 29733 26295 29736
rect 26237 29727 26295 29733
rect 26418 29724 26424 29736
rect 26476 29724 26482 29776
rect 28721 29767 28779 29773
rect 28721 29733 28733 29767
rect 28767 29764 28779 29767
rect 28902 29764 28908 29776
rect 28767 29736 28908 29764
rect 28767 29733 28779 29736
rect 28721 29727 28779 29733
rect 28902 29724 28908 29736
rect 28960 29764 28966 29776
rect 32876 29764 32904 29804
rect 34241 29801 34253 29804
rect 34287 29832 34299 29835
rect 34606 29832 34612 29844
rect 34287 29804 34612 29832
rect 34287 29801 34299 29804
rect 34241 29795 34299 29801
rect 34606 29792 34612 29804
rect 34664 29792 34670 29844
rect 35434 29792 35440 29844
rect 35492 29792 35498 29844
rect 36262 29792 36268 29844
rect 36320 29792 36326 29844
rect 38194 29792 38200 29844
rect 38252 29792 38258 29844
rect 28960 29736 30788 29764
rect 28960 29724 28966 29736
rect 30760 29708 30788 29736
rect 31220 29736 32904 29764
rect 22848 29668 28488 29696
rect 21468 29600 21680 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 8202 29560 8208 29572
rect 5767 29532 8208 29560
rect 5767 29529 5779 29532
rect 5721 29523 5779 29529
rect 4672 29464 4844 29492
rect 4672 29452 4678 29464
rect 5074 29452 5080 29504
rect 5132 29492 5138 29504
rect 5626 29492 5632 29504
rect 5132 29464 5632 29492
rect 5132 29452 5138 29464
rect 5626 29452 5632 29464
rect 5684 29492 5690 29504
rect 5736 29492 5764 29523
rect 8202 29520 8208 29532
rect 8260 29520 8266 29572
rect 10134 29520 10140 29572
rect 10192 29520 10198 29572
rect 10873 29563 10931 29569
rect 10873 29529 10885 29563
rect 10919 29560 10931 29563
rect 11790 29560 11796 29572
rect 10919 29532 11796 29560
rect 10919 29529 10931 29532
rect 10873 29523 10931 29529
rect 11790 29520 11796 29532
rect 11848 29520 11854 29572
rect 11882 29520 11888 29572
rect 11940 29520 11946 29572
rect 12342 29520 12348 29572
rect 12400 29560 12406 29572
rect 12621 29563 12679 29569
rect 12621 29560 12633 29563
rect 12400 29532 12633 29560
rect 12400 29520 12406 29532
rect 12621 29529 12633 29532
rect 12667 29529 12679 29563
rect 12621 29523 12679 29529
rect 13449 29563 13507 29569
rect 13449 29529 13461 29563
rect 13495 29560 13507 29563
rect 14182 29560 14188 29572
rect 13495 29532 14188 29560
rect 13495 29529 13507 29532
rect 13449 29523 13507 29529
rect 14182 29520 14188 29532
rect 14240 29520 14246 29572
rect 14277 29563 14335 29569
rect 14277 29529 14289 29563
rect 14323 29560 14335 29563
rect 14458 29560 14464 29572
rect 14323 29532 14464 29560
rect 14323 29529 14335 29532
rect 14277 29523 14335 29529
rect 14458 29520 14464 29532
rect 14516 29560 14522 29572
rect 16114 29560 16120 29572
rect 14516 29532 16120 29560
rect 14516 29520 14522 29532
rect 16114 29520 16120 29532
rect 16172 29520 16178 29572
rect 17678 29520 17684 29572
rect 17736 29520 17742 29572
rect 5684 29464 5764 29492
rect 5684 29452 5690 29464
rect 7558 29452 7564 29504
rect 7616 29452 7622 29504
rect 10152 29492 10180 29520
rect 11698 29492 11704 29504
rect 10152 29464 11704 29492
rect 11698 29452 11704 29464
rect 11756 29492 11762 29504
rect 14090 29492 14096 29504
rect 11756 29464 14096 29492
rect 11756 29452 11762 29464
rect 14090 29452 14096 29464
rect 14148 29452 14154 29504
rect 16574 29452 16580 29504
rect 16632 29452 16638 29504
rect 20346 29452 20352 29504
rect 20404 29492 20410 29504
rect 20456 29492 20484 29591
rect 21652 29560 21680 29600
rect 21726 29588 21732 29640
rect 21784 29628 21790 29640
rect 21910 29628 21916 29640
rect 21784 29600 21916 29628
rect 21784 29588 21790 29600
rect 21910 29588 21916 29600
rect 21968 29588 21974 29640
rect 22465 29631 22523 29637
rect 22465 29597 22477 29631
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 22186 29560 22192 29572
rect 21008 29532 21588 29560
rect 21652 29532 22192 29560
rect 21008 29501 21036 29532
rect 20404 29464 20484 29492
rect 20993 29495 21051 29501
rect 20404 29452 20410 29464
rect 20993 29461 21005 29495
rect 21039 29461 21051 29495
rect 21560 29492 21588 29532
rect 22186 29520 22192 29532
rect 22244 29520 22250 29572
rect 22480 29560 22508 29591
rect 22554 29588 22560 29640
rect 22612 29628 22618 29640
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 22612 29600 22661 29628
rect 22612 29588 22618 29600
rect 22649 29597 22661 29600
rect 22695 29628 22707 29631
rect 23106 29628 23112 29640
rect 22695 29600 23112 29628
rect 22695 29597 22707 29600
rect 22649 29591 22707 29597
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 23290 29588 23296 29640
rect 23348 29588 23354 29640
rect 23382 29588 23388 29640
rect 23440 29628 23446 29640
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 23440 29600 23489 29628
rect 23440 29588 23446 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 26234 29628 26240 29640
rect 23477 29591 23535 29597
rect 26084 29600 26240 29628
rect 26084 29597 26157 29600
rect 22480 29532 23520 29560
rect 22646 29492 22652 29504
rect 21560 29464 22652 29492
rect 20993 29455 21051 29461
rect 22646 29452 22652 29464
rect 22704 29452 22710 29504
rect 23492 29492 23520 29532
rect 23750 29520 23756 29572
rect 23808 29560 23814 29572
rect 25869 29563 25927 29569
rect 26084 29566 26111 29597
rect 25869 29560 25881 29563
rect 23808 29532 25881 29560
rect 23808 29520 23814 29532
rect 25869 29529 25881 29532
rect 25915 29529 25927 29563
rect 26099 29563 26111 29566
rect 26145 29563 26157 29597
rect 26234 29588 26240 29600
rect 26292 29588 26298 29640
rect 26973 29631 27031 29637
rect 26973 29597 26985 29631
rect 27019 29597 27031 29631
rect 26973 29591 27031 29597
rect 26099 29557 26157 29563
rect 26988 29560 27016 29591
rect 27430 29588 27436 29640
rect 27488 29588 27494 29640
rect 28460 29637 28488 29668
rect 28810 29656 28816 29708
rect 28868 29656 28874 29708
rect 30742 29656 30748 29708
rect 30800 29656 30806 29708
rect 28445 29631 28503 29637
rect 28445 29597 28457 29631
rect 28491 29597 28503 29631
rect 29270 29628 29276 29640
rect 28445 29591 28503 29597
rect 28966 29600 29276 29628
rect 27246 29560 27252 29572
rect 25869 29523 25927 29529
rect 26206 29532 27252 29560
rect 25130 29492 25136 29504
rect 23492 29464 25136 29492
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 25884 29492 25912 29523
rect 26206 29492 26234 29532
rect 27246 29520 27252 29532
rect 27304 29520 27310 29572
rect 28966 29560 28994 29600
rect 29270 29588 29276 29600
rect 29328 29588 29334 29640
rect 29730 29588 29736 29640
rect 29788 29588 29794 29640
rect 29914 29637 29920 29640
rect 29881 29631 29920 29637
rect 29881 29597 29893 29631
rect 29881 29591 29920 29597
rect 29914 29588 29920 29591
rect 29972 29588 29978 29640
rect 30006 29588 30012 29640
rect 30064 29588 30070 29640
rect 30282 29637 30288 29640
rect 30239 29631 30288 29637
rect 30239 29597 30251 29631
rect 30285 29597 30288 29631
rect 30239 29591 30288 29597
rect 30282 29588 30288 29591
rect 30340 29588 30346 29640
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 31021 29631 31079 29637
rect 31021 29628 31033 29631
rect 30432 29600 31033 29628
rect 30432 29588 30438 29600
rect 31021 29597 31033 29600
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 31114 29631 31172 29637
rect 31114 29597 31126 29631
rect 31160 29628 31172 29631
rect 31220 29628 31248 29736
rect 36354 29656 36360 29708
rect 36412 29696 36418 29708
rect 36817 29699 36875 29705
rect 36817 29696 36829 29699
rect 36412 29668 36829 29696
rect 36412 29656 36418 29668
rect 36817 29665 36829 29668
rect 36863 29665 36875 29699
rect 36817 29659 36875 29665
rect 31160 29600 31248 29628
rect 31160 29597 31172 29600
rect 31114 29591 31172 29597
rect 28368 29532 28994 29560
rect 29181 29563 29239 29569
rect 25884 29464 26234 29492
rect 27062 29452 27068 29504
rect 27120 29492 27126 29504
rect 28368 29492 28396 29532
rect 29181 29529 29193 29563
rect 29227 29560 29239 29563
rect 29638 29560 29644 29572
rect 29227 29532 29644 29560
rect 29227 29529 29239 29532
rect 29181 29523 29239 29529
rect 29638 29520 29644 29532
rect 29696 29520 29702 29572
rect 30098 29520 30104 29572
rect 30156 29520 30162 29572
rect 27120 29464 28396 29492
rect 27120 29452 27126 29464
rect 28442 29452 28448 29504
rect 28500 29492 28506 29504
rect 31128 29492 31156 29591
rect 31478 29588 31484 29640
rect 31536 29637 31542 29640
rect 31536 29628 31544 29637
rect 31536 29600 31581 29628
rect 31536 29591 31544 29600
rect 31536 29588 31542 29591
rect 32398 29588 32404 29640
rect 32456 29588 32462 29640
rect 32861 29631 32919 29637
rect 32861 29597 32873 29631
rect 32907 29628 32919 29631
rect 32907 29600 33364 29628
rect 32907 29597 32919 29600
rect 32861 29591 32919 29597
rect 33336 29572 33364 29600
rect 33410 29588 33416 29640
rect 33468 29628 33474 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 33468 29600 34897 29628
rect 33468 29588 33474 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29628 35311 29631
rect 35434 29628 35440 29640
rect 35299 29600 35440 29628
rect 35299 29597 35311 29600
rect 35253 29591 35311 29597
rect 35434 29588 35440 29600
rect 35492 29588 35498 29640
rect 36078 29588 36084 29640
rect 36136 29588 36142 29640
rect 37084 29631 37142 29637
rect 37084 29597 37096 29631
rect 37130 29628 37142 29631
rect 37458 29628 37464 29640
rect 37130 29600 37464 29628
rect 37130 29597 37142 29600
rect 37084 29591 37142 29597
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 31294 29520 31300 29572
rect 31352 29520 31358 29572
rect 31389 29563 31447 29569
rect 31389 29529 31401 29563
rect 31435 29529 31447 29563
rect 32125 29563 32183 29569
rect 32125 29560 32137 29563
rect 31389 29523 31447 29529
rect 31680 29532 32137 29560
rect 28500 29464 31156 29492
rect 31404 29492 31432 29523
rect 31478 29492 31484 29504
rect 31404 29464 31484 29492
rect 28500 29452 28506 29464
rect 31478 29452 31484 29464
rect 31536 29452 31542 29504
rect 31680 29501 31708 29532
rect 32125 29529 32137 29532
rect 32171 29560 32183 29563
rect 32490 29560 32496 29572
rect 32171 29532 32496 29560
rect 32171 29529 32183 29532
rect 32125 29523 32183 29529
rect 32490 29520 32496 29532
rect 32548 29520 32554 29572
rect 33134 29569 33140 29572
rect 33128 29560 33140 29569
rect 33095 29532 33140 29560
rect 33128 29523 33140 29532
rect 33134 29520 33140 29523
rect 33192 29520 33198 29572
rect 33318 29520 33324 29572
rect 33376 29520 33382 29572
rect 34514 29520 34520 29572
rect 34572 29560 34578 29572
rect 35066 29560 35072 29572
rect 34572 29532 35072 29560
rect 34572 29520 34578 29532
rect 35066 29520 35072 29532
rect 35124 29520 35130 29572
rect 35158 29520 35164 29572
rect 35216 29520 35222 29572
rect 31665 29495 31723 29501
rect 31665 29461 31677 29495
rect 31711 29461 31723 29495
rect 31665 29455 31723 29461
rect 32306 29452 32312 29504
rect 32364 29452 32370 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5810 29248 5816 29300
rect 5868 29288 5874 29300
rect 9401 29291 9459 29297
rect 5868 29260 9260 29288
rect 5868 29248 5874 29260
rect 3326 29180 3332 29232
rect 3384 29220 3390 29232
rect 3970 29220 3976 29232
rect 3384 29192 3976 29220
rect 3384 29180 3390 29192
rect 3970 29180 3976 29192
rect 4028 29220 4034 29232
rect 4341 29223 4399 29229
rect 4341 29220 4353 29223
rect 4028 29192 4353 29220
rect 4028 29180 4034 29192
rect 4341 29189 4353 29192
rect 4387 29189 4399 29223
rect 4341 29183 4399 29189
rect 4433 29223 4491 29229
rect 4433 29189 4445 29223
rect 4479 29220 4491 29223
rect 4798 29220 4804 29232
rect 4479 29192 4804 29220
rect 4479 29189 4491 29192
rect 4433 29183 4491 29189
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 6733 29223 6791 29229
rect 5276 29192 6684 29220
rect 5276 29164 5304 29192
rect 3142 29112 3148 29164
rect 3200 29152 3206 29164
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 3200 29124 4261 29152
rect 3200 29112 3206 29124
rect 4249 29121 4261 29124
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29152 4675 29155
rect 4890 29152 4896 29164
rect 4663 29124 4896 29152
rect 4663 29121 4675 29124
rect 4617 29115 4675 29121
rect 4264 29084 4292 29115
rect 4890 29112 4896 29124
rect 4948 29112 4954 29164
rect 5258 29112 5264 29164
rect 5316 29112 5322 29164
rect 5537 29155 5595 29161
rect 5537 29121 5549 29155
rect 5583 29152 5595 29155
rect 5994 29152 6000 29164
rect 5583 29124 6000 29152
rect 5583 29121 5595 29124
rect 5537 29115 5595 29121
rect 5994 29112 6000 29124
rect 6052 29112 6058 29164
rect 6656 29152 6684 29192
rect 6733 29189 6745 29223
rect 6779 29220 6791 29223
rect 6822 29220 6828 29232
rect 6779 29192 6828 29220
rect 6779 29189 6791 29192
rect 6733 29183 6791 29189
rect 6822 29180 6828 29192
rect 6880 29180 6886 29232
rect 6914 29180 6920 29232
rect 6972 29180 6978 29232
rect 7006 29180 7012 29232
rect 7064 29220 7070 29232
rect 8941 29223 8999 29229
rect 8941 29220 8953 29223
rect 7064 29192 8953 29220
rect 7064 29180 7070 29192
rect 8941 29189 8953 29192
rect 8987 29189 8999 29223
rect 8941 29183 8999 29189
rect 7466 29152 7472 29164
rect 6656 29124 7472 29152
rect 7466 29112 7472 29124
rect 7524 29112 7530 29164
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29121 8171 29155
rect 8113 29115 8171 29121
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 8754 29152 8760 29164
rect 8435 29124 8760 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 5166 29084 5172 29096
rect 4264 29056 5172 29084
rect 5166 29044 5172 29056
rect 5224 29044 5230 29096
rect 5442 29044 5448 29096
rect 5500 29044 5506 29096
rect 6012 29084 6040 29112
rect 8128 29084 8156 29115
rect 8754 29112 8760 29124
rect 8812 29112 8818 29164
rect 9232 29161 9260 29260
rect 9401 29257 9413 29291
rect 9447 29257 9459 29291
rect 9401 29251 9459 29257
rect 9416 29220 9444 29251
rect 11146 29248 11152 29300
rect 11204 29248 11210 29300
rect 11974 29288 11980 29300
rect 11348 29260 11980 29288
rect 11348 29220 11376 29260
rect 11974 29248 11980 29260
rect 12032 29288 12038 29300
rect 14645 29291 14703 29297
rect 12032 29260 12664 29288
rect 12032 29248 12038 29260
rect 9416 29192 11376 29220
rect 11698 29180 11704 29232
rect 11756 29180 11762 29232
rect 11885 29223 11943 29229
rect 11885 29220 11897 29223
rect 11808 29192 11897 29220
rect 9217 29155 9275 29161
rect 9217 29121 9229 29155
rect 9263 29152 9275 29155
rect 9490 29152 9496 29164
rect 9263 29124 9496 29152
rect 9263 29121 9275 29124
rect 9217 29115 9275 29121
rect 9490 29112 9496 29124
rect 9548 29112 9554 29164
rect 9950 29112 9956 29164
rect 10008 29112 10014 29164
rect 10042 29112 10048 29164
rect 10100 29112 10106 29164
rect 10965 29155 11023 29161
rect 10965 29121 10977 29155
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 6012 29056 8156 29084
rect 8202 29044 8208 29096
rect 8260 29084 8266 29096
rect 9033 29087 9091 29093
rect 9033 29084 9045 29087
rect 8260 29056 9045 29084
rect 8260 29044 8266 29056
rect 9033 29053 9045 29056
rect 9079 29053 9091 29087
rect 9033 29047 9091 29053
rect 4065 29019 4123 29025
rect 4065 28985 4077 29019
rect 4111 29016 4123 29019
rect 4614 29016 4620 29028
rect 4111 28988 4620 29016
rect 4111 28985 4123 28988
rect 4065 28979 4123 28985
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 5074 28976 5080 29028
rect 5132 28976 5138 29028
rect 7742 28976 7748 29028
rect 7800 29016 7806 29028
rect 8113 29019 8171 29025
rect 8113 29016 8125 29019
rect 7800 28988 8125 29016
rect 7800 28976 7806 28988
rect 8113 28985 8125 28988
rect 8159 28985 8171 29019
rect 9048 29016 9076 29047
rect 9582 29044 9588 29096
rect 9640 29084 9646 29096
rect 10980 29084 11008 29115
rect 11146 29112 11152 29164
rect 11204 29112 11210 29164
rect 9640 29056 11008 29084
rect 9640 29044 9646 29056
rect 9674 29016 9680 29028
rect 9048 28988 9680 29016
rect 8113 28979 8171 28985
rect 9674 28976 9680 28988
rect 9732 29016 9738 29028
rect 10502 29016 10508 29028
rect 9732 28988 10508 29016
rect 9732 28976 9738 28988
rect 10502 28976 10508 28988
rect 10560 28976 10566 29028
rect 10980 29016 11008 29056
rect 11808 29016 11836 29192
rect 11885 29189 11897 29192
rect 11931 29189 11943 29223
rect 11885 29183 11943 29189
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 12434 29152 12440 29164
rect 12207 29124 12440 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 12434 29112 12440 29124
rect 12492 29112 12498 29164
rect 12636 29161 12664 29260
rect 14645 29257 14657 29291
rect 14691 29288 14703 29291
rect 14826 29288 14832 29300
rect 14691 29260 14832 29288
rect 14691 29257 14703 29260
rect 14645 29251 14703 29257
rect 14826 29248 14832 29260
rect 14884 29248 14890 29300
rect 16206 29248 16212 29300
rect 16264 29288 16270 29300
rect 16301 29291 16359 29297
rect 16301 29288 16313 29291
rect 16264 29260 16313 29288
rect 16264 29248 16270 29260
rect 16301 29257 16313 29260
rect 16347 29257 16359 29291
rect 16301 29251 16359 29257
rect 18414 29248 18420 29300
rect 18472 29288 18478 29300
rect 19245 29291 19303 29297
rect 19245 29288 19257 29291
rect 18472 29260 19257 29288
rect 18472 29248 18478 29260
rect 19245 29257 19257 29260
rect 19291 29257 19303 29291
rect 19245 29251 19303 29257
rect 19334 29248 19340 29300
rect 19392 29288 19398 29300
rect 19392 29260 22692 29288
rect 19392 29248 19398 29260
rect 13814 29180 13820 29232
rect 13872 29220 13878 29232
rect 14277 29223 14335 29229
rect 14277 29220 14289 29223
rect 13872 29192 14289 29220
rect 13872 29180 13878 29192
rect 14277 29189 14289 29192
rect 14323 29189 14335 29223
rect 14277 29183 14335 29189
rect 14369 29223 14427 29229
rect 14369 29189 14381 29223
rect 14415 29220 14427 29223
rect 16574 29220 16580 29232
rect 14415 29192 16580 29220
rect 14415 29189 14427 29192
rect 14369 29183 14427 29189
rect 16574 29180 16580 29192
rect 16632 29220 16638 29232
rect 17405 29223 17463 29229
rect 16632 29192 17080 29220
rect 16632 29180 16638 29192
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 12805 29155 12863 29161
rect 12805 29121 12817 29155
rect 12851 29152 12863 29155
rect 12986 29152 12992 29164
rect 12851 29124 12992 29152
rect 12851 29121 12863 29124
rect 12805 29115 12863 29121
rect 12986 29112 12992 29124
rect 13044 29112 13050 29164
rect 13262 29112 13268 29164
rect 13320 29112 13326 29164
rect 13449 29155 13507 29161
rect 13449 29121 13461 29155
rect 13495 29152 13507 29155
rect 13906 29152 13912 29164
rect 13495 29124 13912 29152
rect 13495 29121 13507 29124
rect 13449 29115 13507 29121
rect 13906 29112 13912 29124
rect 13964 29112 13970 29164
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 14461 29155 14519 29161
rect 14461 29121 14473 29155
rect 14507 29121 14519 29155
rect 14461 29115 14519 29121
rect 16117 29155 16175 29161
rect 16117 29121 16129 29155
rect 16163 29152 16175 29155
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16163 29124 16865 29152
rect 16163 29121 16175 29124
rect 16117 29115 16175 29121
rect 16853 29121 16865 29124
rect 16899 29152 16911 29155
rect 16942 29152 16948 29164
rect 16899 29124 16948 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 13280 29084 13308 29112
rect 14476 29084 14504 29115
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 17052 29161 17080 29192
rect 17405 29189 17417 29223
rect 17451 29220 17463 29223
rect 20162 29220 20168 29232
rect 17451 29192 20168 29220
rect 17451 29189 17463 29192
rect 17405 29183 17463 29189
rect 20162 29180 20168 29192
rect 20220 29180 20226 29232
rect 20438 29220 20444 29232
rect 20272 29192 20444 29220
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17586 29152 17592 29164
rect 17037 29115 17095 29121
rect 17144 29124 17592 29152
rect 13280 29056 13584 29084
rect 10980 28988 11836 29016
rect 5350 28908 5356 28960
rect 5408 28948 5414 28960
rect 5902 28948 5908 28960
rect 5408 28920 5908 28948
rect 5408 28908 5414 28920
rect 5902 28908 5908 28920
rect 5960 28908 5966 28960
rect 6638 28908 6644 28960
rect 6696 28908 6702 28960
rect 6822 28908 6828 28960
rect 6880 28948 6886 28960
rect 8941 28951 8999 28957
rect 8941 28948 8953 28951
rect 6880 28920 8953 28948
rect 6880 28908 6886 28920
rect 8941 28917 8953 28920
rect 8987 28948 8999 28951
rect 9122 28948 9128 28960
rect 8987 28920 9128 28948
rect 8987 28917 8999 28920
rect 8941 28911 8999 28917
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 9953 28951 10011 28957
rect 9953 28917 9965 28951
rect 9999 28948 10011 28951
rect 10134 28948 10140 28960
rect 9999 28920 10140 28948
rect 9999 28917 10011 28920
rect 9953 28911 10011 28917
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 11146 28908 11152 28960
rect 11204 28948 11210 28960
rect 11885 28951 11943 28957
rect 11885 28948 11897 28951
rect 11204 28920 11897 28948
rect 11204 28908 11210 28920
rect 11885 28917 11897 28920
rect 11931 28948 11943 28951
rect 11974 28948 11980 28960
rect 11931 28920 11980 28948
rect 11931 28917 11943 28920
rect 11885 28911 11943 28917
rect 11974 28908 11980 28920
rect 12032 28908 12038 28960
rect 12621 28951 12679 28957
rect 12621 28917 12633 28951
rect 12667 28948 12679 28951
rect 13170 28948 13176 28960
rect 12667 28920 13176 28948
rect 12667 28917 12679 28920
rect 12621 28911 12679 28917
rect 13170 28908 13176 28920
rect 13228 28908 13234 28960
rect 13446 28908 13452 28960
rect 13504 28908 13510 28960
rect 13556 28948 13584 29056
rect 13648 29056 14504 29084
rect 13648 29025 13676 29056
rect 14734 29044 14740 29096
rect 14792 29084 14798 29096
rect 15838 29084 15844 29096
rect 14792 29056 15844 29084
rect 14792 29044 14798 29056
rect 15838 29044 15844 29056
rect 15896 29044 15902 29096
rect 15933 29087 15991 29093
rect 15933 29053 15945 29087
rect 15979 29084 15991 29087
rect 17144 29084 17172 29124
rect 17586 29112 17592 29124
rect 17644 29112 17650 29164
rect 17865 29155 17923 29161
rect 17865 29121 17877 29155
rect 17911 29152 17923 29155
rect 17954 29152 17960 29164
rect 17911 29124 17960 29152
rect 17911 29121 17923 29124
rect 17865 29115 17923 29121
rect 17954 29112 17960 29124
rect 18012 29152 18018 29164
rect 18785 29155 18843 29161
rect 18012 29124 18460 29152
rect 18012 29112 18018 29124
rect 15979 29056 17172 29084
rect 15979 29053 15991 29056
rect 15933 29047 15991 29053
rect 13633 29019 13691 29025
rect 13633 28985 13645 29019
rect 13679 28985 13691 29019
rect 13633 28979 13691 28985
rect 13906 28976 13912 29028
rect 13964 29016 13970 29028
rect 14752 29016 14780 29044
rect 13964 28988 14780 29016
rect 13964 28976 13970 28988
rect 15102 28976 15108 29028
rect 15160 29016 15166 29028
rect 15948 29016 15976 29047
rect 17494 29044 17500 29096
rect 17552 29084 17558 29096
rect 18233 29087 18291 29093
rect 18233 29084 18245 29087
rect 17552 29056 18245 29084
rect 17552 29044 17558 29056
rect 18233 29053 18245 29056
rect 18279 29053 18291 29087
rect 18432 29084 18460 29124
rect 18785 29121 18797 29155
rect 18831 29152 18843 29155
rect 18966 29152 18972 29164
rect 18831 29124 18972 29152
rect 18831 29121 18843 29124
rect 18785 29115 18843 29121
rect 18966 29112 18972 29124
rect 19024 29152 19030 29164
rect 19521 29155 19579 29161
rect 19521 29152 19533 29155
rect 19024 29124 19533 29152
rect 19024 29112 19030 29124
rect 19521 29121 19533 29124
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 19610 29112 19616 29164
rect 19668 29112 19674 29164
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 20272 29152 20300 29192
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 19935 29124 20300 29152
rect 20349 29155 20407 29161
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 20349 29121 20361 29155
rect 20395 29152 20407 29155
rect 20990 29152 20996 29164
rect 20395 29124 20996 29152
rect 20395 29121 20407 29124
rect 20349 29115 20407 29121
rect 18506 29084 18512 29096
rect 18432 29056 18512 29084
rect 18233 29047 18291 29053
rect 18506 29044 18512 29056
rect 18564 29084 18570 29096
rect 19150 29084 19156 29096
rect 18564 29056 19156 29084
rect 18564 29044 18570 29056
rect 19150 29044 19156 29056
rect 19208 29044 19214 29096
rect 19242 29044 19248 29096
rect 19300 29084 19306 29096
rect 19720 29084 19748 29115
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 22186 29112 22192 29164
rect 22244 29152 22250 29164
rect 22557 29155 22615 29161
rect 22557 29152 22569 29155
rect 22244 29124 22569 29152
rect 22244 29112 22250 29124
rect 22557 29121 22569 29124
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 19300 29056 19748 29084
rect 19300 29044 19306 29056
rect 19794 29044 19800 29096
rect 19852 29084 19858 29096
rect 20254 29084 20260 29096
rect 19852 29056 20260 29084
rect 19852 29044 19858 29056
rect 20254 29044 20260 29056
rect 20312 29084 20318 29096
rect 20625 29087 20683 29093
rect 20625 29084 20637 29087
rect 20312 29056 20637 29084
rect 20312 29044 20318 29056
rect 20625 29053 20637 29056
rect 20671 29053 20683 29087
rect 20625 29047 20683 29053
rect 20809 29087 20867 29093
rect 20809 29053 20821 29087
rect 20855 29084 20867 29087
rect 22462 29084 22468 29096
rect 20855 29056 22468 29084
rect 20855 29053 20867 29056
rect 20809 29047 20867 29053
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 22664 29084 22692 29260
rect 23382 29248 23388 29300
rect 23440 29248 23446 29300
rect 23658 29288 23664 29300
rect 23584 29260 23664 29288
rect 22741 29155 22799 29161
rect 22741 29121 22753 29155
rect 22787 29152 22799 29155
rect 23400 29152 23428 29248
rect 23584 29161 23612 29260
rect 23658 29248 23664 29260
rect 23716 29248 23722 29300
rect 24946 29248 24952 29300
rect 25004 29248 25010 29300
rect 25682 29288 25688 29300
rect 25056 29260 25688 29288
rect 24302 29220 24308 29232
rect 23676 29192 24308 29220
rect 23676 29161 23704 29192
rect 24302 29180 24308 29192
rect 24360 29180 24366 29232
rect 25056 29220 25084 29260
rect 25682 29248 25688 29260
rect 25740 29288 25746 29300
rect 27154 29288 27160 29300
rect 25740 29260 27160 29288
rect 25740 29248 25746 29260
rect 27154 29248 27160 29260
rect 27212 29248 27218 29300
rect 30098 29248 30104 29300
rect 30156 29288 30162 29300
rect 30156 29260 31800 29288
rect 30156 29248 30162 29260
rect 24872 29192 25084 29220
rect 22787 29124 23428 29152
rect 23569 29155 23627 29161
rect 22787 29121 22799 29124
rect 22741 29115 22799 29121
rect 23569 29121 23581 29155
rect 23615 29121 23627 29155
rect 23569 29115 23627 29121
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29121 23719 29155
rect 23661 29115 23719 29121
rect 23750 29112 23756 29164
rect 23808 29112 23814 29164
rect 23842 29112 23848 29164
rect 23900 29152 23906 29164
rect 24872 29152 24900 29192
rect 25314 29180 25320 29232
rect 25372 29220 25378 29232
rect 27062 29220 27068 29232
rect 25372 29192 27068 29220
rect 25372 29180 25378 29192
rect 27062 29180 27068 29192
rect 27120 29220 27126 29232
rect 27982 29220 27988 29232
rect 27120 29192 27988 29220
rect 27120 29180 27126 29192
rect 27982 29180 27988 29192
rect 28040 29180 28046 29232
rect 28258 29180 28264 29232
rect 28316 29220 28322 29232
rect 28445 29223 28503 29229
rect 28445 29220 28457 29223
rect 28316 29192 28457 29220
rect 28316 29180 28322 29192
rect 28445 29189 28457 29192
rect 28491 29189 28503 29223
rect 28445 29183 28503 29189
rect 28537 29223 28595 29229
rect 28537 29189 28549 29223
rect 28583 29220 28595 29223
rect 28626 29220 28632 29232
rect 28583 29192 28632 29220
rect 28583 29189 28595 29192
rect 28537 29183 28595 29189
rect 28626 29180 28632 29192
rect 28684 29220 28690 29232
rect 31665 29223 31723 29229
rect 31665 29220 31677 29223
rect 28684 29192 30328 29220
rect 28684 29180 28690 29192
rect 23900 29124 24900 29152
rect 23900 29112 23906 29124
rect 24946 29112 24952 29164
rect 25004 29152 25010 29164
rect 25498 29152 25504 29164
rect 25004 29124 25504 29152
rect 25004 29112 25010 29124
rect 25498 29112 25504 29124
rect 25556 29152 25562 29164
rect 25961 29155 26019 29161
rect 25961 29152 25973 29155
rect 25556 29124 25973 29152
rect 25556 29112 25562 29124
rect 25961 29121 25973 29124
rect 26007 29121 26019 29155
rect 25961 29115 26019 29121
rect 27154 29112 27160 29164
rect 27212 29112 27218 29164
rect 27246 29112 27252 29164
rect 27304 29152 27310 29164
rect 27525 29155 27583 29161
rect 27525 29152 27537 29155
rect 27304 29124 27537 29152
rect 27304 29112 27310 29124
rect 27525 29121 27537 29124
rect 27571 29121 27583 29155
rect 27525 29115 27583 29121
rect 28353 29155 28411 29161
rect 28353 29121 28365 29155
rect 28399 29121 28411 29155
rect 28353 29115 28411 29121
rect 28721 29155 28779 29161
rect 28721 29121 28733 29155
rect 28767 29152 28779 29155
rect 29086 29152 29092 29164
rect 28767 29124 29092 29152
rect 28767 29121 28779 29124
rect 28721 29115 28779 29121
rect 23382 29084 23388 29096
rect 22664 29056 23388 29084
rect 23382 29044 23388 29056
rect 23440 29084 23446 29096
rect 25038 29084 25044 29096
rect 23440 29056 25044 29084
rect 23440 29044 23446 29056
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 25133 29087 25191 29093
rect 25133 29053 25145 29087
rect 25179 29053 25191 29087
rect 25133 29047 25191 29053
rect 15160 28988 15976 29016
rect 18325 29019 18383 29025
rect 15160 28976 15166 28988
rect 18325 28985 18337 29019
rect 18371 29016 18383 29019
rect 18874 29016 18880 29028
rect 18371 28988 18880 29016
rect 18371 28985 18383 28988
rect 18325 28979 18383 28985
rect 18874 28976 18880 28988
rect 18932 28976 18938 29028
rect 19610 28976 19616 29028
rect 19668 29016 19674 29028
rect 20441 29019 20499 29025
rect 20441 29016 20453 29019
rect 19668 28988 20453 29016
rect 19668 28976 19674 28988
rect 20441 28985 20453 28988
rect 20487 29016 20499 29019
rect 20714 29016 20720 29028
rect 20487 28988 20720 29016
rect 20487 28985 20499 28988
rect 20441 28979 20499 28985
rect 20714 28976 20720 28988
rect 20772 29016 20778 29028
rect 21450 29016 21456 29028
rect 20772 28988 21456 29016
rect 20772 28976 20778 28988
rect 21450 28976 21456 28988
rect 21508 28976 21514 29028
rect 22094 28976 22100 29028
rect 22152 29016 22158 29028
rect 22925 29019 22983 29025
rect 22925 29016 22937 29019
rect 22152 28988 22937 29016
rect 22152 28976 22158 28988
rect 22925 28985 22937 28988
rect 22971 28985 22983 29019
rect 22925 28979 22983 28985
rect 23014 28976 23020 29028
rect 23072 29016 23078 29028
rect 24854 29016 24860 29028
rect 23072 28988 24860 29016
rect 23072 28976 23078 28988
rect 24854 28976 24860 28988
rect 24912 28976 24918 29028
rect 25148 29016 25176 29047
rect 25222 29044 25228 29096
rect 25280 29044 25286 29096
rect 25314 29044 25320 29096
rect 25372 29044 25378 29096
rect 25409 29087 25467 29093
rect 25409 29053 25421 29087
rect 25455 29084 25467 29087
rect 25682 29084 25688 29096
rect 25455 29056 25688 29084
rect 25455 29053 25467 29056
rect 25409 29047 25467 29053
rect 25682 29044 25688 29056
rect 25740 29044 25746 29096
rect 26050 29044 26056 29096
rect 26108 29044 26114 29096
rect 26970 29044 26976 29096
rect 27028 29084 27034 29096
rect 27341 29087 27399 29093
rect 27341 29084 27353 29087
rect 27028 29056 27353 29084
rect 27028 29044 27034 29056
rect 27341 29053 27353 29056
rect 27387 29053 27399 29087
rect 27341 29047 27399 29053
rect 28258 29044 28264 29096
rect 28316 29084 28322 29096
rect 28368 29084 28396 29115
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 29181 29155 29239 29161
rect 29181 29121 29193 29155
rect 29227 29121 29239 29155
rect 29181 29115 29239 29121
rect 28316 29056 28396 29084
rect 28316 29044 28322 29056
rect 28994 29044 29000 29096
rect 29052 29084 29058 29096
rect 29196 29084 29224 29115
rect 29052 29056 29224 29084
rect 29365 29087 29423 29093
rect 29052 29044 29058 29056
rect 29365 29053 29377 29087
rect 29411 29053 29423 29087
rect 30300 29084 30328 29192
rect 30944 29192 31677 29220
rect 30944 29164 30972 29192
rect 31665 29189 31677 29192
rect 31711 29189 31723 29223
rect 31665 29183 31723 29189
rect 30377 29155 30435 29161
rect 30377 29121 30389 29155
rect 30423 29152 30435 29155
rect 30650 29152 30656 29164
rect 30423 29124 30656 29152
rect 30423 29121 30435 29124
rect 30377 29115 30435 29121
rect 30650 29112 30656 29124
rect 30708 29112 30714 29164
rect 30745 29155 30803 29161
rect 30745 29121 30757 29155
rect 30791 29152 30803 29155
rect 30926 29152 30932 29164
rect 30791 29124 30932 29152
rect 30791 29121 30803 29124
rect 30745 29115 30803 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31297 29155 31355 29161
rect 31297 29121 31309 29155
rect 31343 29152 31355 29155
rect 31386 29152 31392 29164
rect 31343 29124 31392 29152
rect 31343 29121 31355 29124
rect 31297 29115 31355 29121
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31478 29112 31484 29164
rect 31536 29112 31542 29164
rect 31772 29152 31800 29260
rect 32490 29248 32496 29300
rect 32548 29248 32554 29300
rect 32674 29248 32680 29300
rect 32732 29248 32738 29300
rect 32306 29180 32312 29232
rect 32364 29220 32370 29232
rect 33042 29220 33048 29232
rect 32364 29192 33048 29220
rect 32364 29180 32370 29192
rect 33042 29180 33048 29192
rect 33100 29180 33106 29232
rect 35066 29180 35072 29232
rect 35124 29220 35130 29232
rect 35342 29220 35348 29232
rect 35124 29192 35348 29220
rect 35124 29180 35130 29192
rect 35342 29180 35348 29192
rect 35400 29180 35406 29232
rect 37921 29223 37979 29229
rect 37921 29189 37933 29223
rect 37967 29220 37979 29223
rect 38010 29220 38016 29232
rect 37967 29192 38016 29220
rect 37967 29189 37979 29192
rect 37921 29183 37979 29189
rect 38010 29180 38016 29192
rect 38068 29180 38074 29232
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 31772 29124 34897 29152
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 35161 29155 35219 29161
rect 35161 29121 35173 29155
rect 35207 29121 35219 29155
rect 35161 29115 35219 29121
rect 35253 29155 35311 29161
rect 35253 29121 35265 29155
rect 35299 29152 35311 29155
rect 35434 29152 35440 29164
rect 35299 29124 35440 29152
rect 35299 29121 35311 29124
rect 35253 29115 35311 29121
rect 31496 29084 31524 29112
rect 30300 29056 31524 29084
rect 29365 29047 29423 29053
rect 26234 29016 26240 29028
rect 25148 28988 26240 29016
rect 26234 28976 26240 28988
rect 26292 29016 26298 29028
rect 26329 29019 26387 29025
rect 26329 29016 26341 29019
rect 26292 28988 26341 29016
rect 26292 28976 26298 28988
rect 26329 28985 26341 28988
rect 26375 28985 26387 29019
rect 26329 28979 26387 28985
rect 28166 28976 28172 29028
rect 28224 28976 28230 29028
rect 29086 28976 29092 29028
rect 29144 29016 29150 29028
rect 29380 29016 29408 29047
rect 35176 29016 35204 29115
rect 35434 29112 35440 29124
rect 35492 29112 35498 29164
rect 36170 29112 36176 29164
rect 36228 29152 36234 29164
rect 36449 29155 36507 29161
rect 36449 29152 36461 29155
rect 36228 29124 36461 29152
rect 36228 29112 36234 29124
rect 36449 29121 36461 29124
rect 36495 29121 36507 29155
rect 36449 29115 36507 29121
rect 37550 29112 37556 29164
rect 37608 29112 37614 29164
rect 36725 29087 36783 29093
rect 36725 29053 36737 29087
rect 36771 29084 36783 29087
rect 39022 29084 39028 29096
rect 36771 29056 39028 29084
rect 36771 29053 36783 29056
rect 36725 29047 36783 29053
rect 39022 29044 39028 29056
rect 39080 29044 39086 29096
rect 29144 28988 29408 29016
rect 31726 28994 35204 29016
rect 31680 28988 35204 28994
rect 29144 28976 29150 28988
rect 15120 28948 15148 28976
rect 31680 28966 31754 28988
rect 13556 28920 15148 28948
rect 18417 28951 18475 28957
rect 18417 28917 18429 28951
rect 18463 28948 18475 28951
rect 21082 28948 21088 28960
rect 18463 28920 21088 28948
rect 18463 28917 18475 28920
rect 18417 28911 18475 28917
rect 21082 28908 21088 28920
rect 21140 28908 21146 28960
rect 25038 28908 25044 28960
rect 25096 28948 25102 28960
rect 25590 28948 25596 28960
rect 25096 28920 25596 28948
rect 25096 28908 25102 28920
rect 25590 28908 25596 28920
rect 25648 28948 25654 28960
rect 25961 28951 26019 28957
rect 25961 28948 25973 28951
rect 25648 28920 25973 28948
rect 25648 28908 25654 28920
rect 25961 28917 25973 28920
rect 26007 28917 26019 28951
rect 25961 28911 26019 28917
rect 27249 28951 27307 28957
rect 27249 28917 27261 28951
rect 27295 28948 27307 28951
rect 28902 28948 28908 28960
rect 27295 28920 28908 28948
rect 27295 28917 27307 28920
rect 27249 28911 27307 28917
rect 28902 28908 28908 28920
rect 28960 28908 28966 28960
rect 31110 28908 31116 28960
rect 31168 28948 31174 28960
rect 31680 28948 31708 28966
rect 31168 28920 31708 28948
rect 31168 28908 31174 28920
rect 32398 28908 32404 28960
rect 32456 28948 32462 28960
rect 32493 28951 32551 28957
rect 32493 28948 32505 28951
rect 32456 28920 32505 28948
rect 32456 28908 32462 28920
rect 32493 28917 32505 28920
rect 32539 28917 32551 28951
rect 32493 28911 32551 28917
rect 35437 28951 35495 28957
rect 35437 28917 35449 28951
rect 35483 28948 35495 28951
rect 35526 28948 35532 28960
rect 35483 28920 35532 28948
rect 35483 28917 35495 28920
rect 35437 28911 35495 28917
rect 35526 28908 35532 28920
rect 35584 28908 35590 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 3970 28704 3976 28756
rect 4028 28744 4034 28756
rect 4617 28747 4675 28753
rect 4617 28744 4629 28747
rect 4028 28716 4629 28744
rect 4028 28704 4034 28716
rect 4617 28713 4629 28716
rect 4663 28713 4675 28747
rect 4617 28707 4675 28713
rect 4982 28704 4988 28756
rect 5040 28744 5046 28756
rect 5350 28744 5356 28756
rect 5040 28716 5356 28744
rect 5040 28704 5046 28716
rect 5350 28704 5356 28716
rect 5408 28704 5414 28756
rect 9214 28704 9220 28756
rect 9272 28744 9278 28756
rect 10321 28747 10379 28753
rect 10321 28744 10333 28747
rect 9272 28716 10333 28744
rect 9272 28704 9278 28716
rect 10321 28713 10333 28716
rect 10367 28713 10379 28747
rect 10321 28707 10379 28713
rect 10520 28716 10732 28744
rect 7469 28679 7527 28685
rect 7469 28676 7481 28679
rect 6932 28648 7481 28676
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28540 4767 28543
rect 4755 28512 5304 28540
rect 4755 28509 4767 28512
rect 4709 28503 4767 28509
rect 5276 28413 5304 28512
rect 5442 28500 5448 28552
rect 5500 28500 5506 28552
rect 6638 28500 6644 28552
rect 6696 28500 6702 28552
rect 6932 28549 6960 28648
rect 7469 28645 7481 28648
rect 7515 28676 7527 28679
rect 9306 28676 9312 28688
rect 7515 28648 9312 28676
rect 7515 28645 7527 28648
rect 7469 28639 7527 28645
rect 9306 28636 9312 28648
rect 9364 28636 9370 28688
rect 9490 28636 9496 28688
rect 9548 28676 9554 28688
rect 10520 28676 10548 28716
rect 9548 28648 10548 28676
rect 9548 28636 9554 28648
rect 10594 28636 10600 28688
rect 10652 28636 10658 28688
rect 10704 28676 10732 28716
rect 11054 28704 11060 28756
rect 11112 28744 11118 28756
rect 11882 28744 11888 28756
rect 11112 28716 11888 28744
rect 11112 28704 11118 28716
rect 11882 28704 11888 28716
rect 11940 28704 11946 28756
rect 11974 28704 11980 28756
rect 12032 28744 12038 28756
rect 12529 28747 12587 28753
rect 12529 28744 12541 28747
rect 12032 28716 12541 28744
rect 12032 28704 12038 28716
rect 12529 28713 12541 28716
rect 12575 28713 12587 28747
rect 12529 28707 12587 28713
rect 15105 28747 15163 28753
rect 15105 28713 15117 28747
rect 15151 28744 15163 28747
rect 15378 28744 15384 28756
rect 15151 28716 15384 28744
rect 15151 28713 15163 28716
rect 15105 28707 15163 28713
rect 15378 28704 15384 28716
rect 15436 28704 15442 28756
rect 16482 28744 16488 28756
rect 16408 28716 16488 28744
rect 10704 28648 12756 28676
rect 8018 28568 8024 28620
rect 8076 28608 8082 28620
rect 10413 28611 10471 28617
rect 8076 28580 9720 28608
rect 8076 28568 8082 28580
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28509 6975 28543
rect 6917 28503 6975 28509
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 7377 28543 7435 28549
rect 7377 28540 7389 28543
rect 7248 28512 7389 28540
rect 7248 28500 7254 28512
rect 7377 28509 7389 28512
rect 7423 28509 7435 28543
rect 7377 28503 7435 28509
rect 7466 28500 7472 28552
rect 7524 28540 7530 28552
rect 7561 28543 7619 28549
rect 7561 28540 7573 28543
rect 7524 28512 7573 28540
rect 7524 28500 7530 28512
rect 7561 28509 7573 28512
rect 7607 28509 7619 28543
rect 7561 28503 7619 28509
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9692 28540 9720 28580
rect 10413 28577 10425 28611
rect 10459 28608 10471 28611
rect 10612 28608 10640 28636
rect 10459 28580 10640 28608
rect 10459 28577 10471 28580
rect 10413 28571 10471 28577
rect 9692 28512 10456 28540
rect 9585 28503 9643 28509
rect 5629 28475 5687 28481
rect 5629 28441 5641 28475
rect 5675 28441 5687 28475
rect 5629 28435 5687 28441
rect 5261 28407 5319 28413
rect 5261 28373 5273 28407
rect 5307 28404 5319 28407
rect 5350 28404 5356 28416
rect 5307 28376 5356 28404
rect 5307 28373 5319 28376
rect 5261 28367 5319 28373
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 5644 28404 5672 28435
rect 6546 28432 6552 28484
rect 6604 28432 6610 28484
rect 9600 28472 9628 28503
rect 9674 28472 9680 28484
rect 9600 28444 9680 28472
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 10134 28432 10140 28484
rect 10192 28472 10198 28484
rect 10321 28475 10379 28481
rect 10321 28472 10333 28475
rect 10192 28444 10333 28472
rect 10192 28432 10198 28444
rect 10321 28441 10333 28444
rect 10367 28441 10379 28475
rect 10428 28472 10456 28512
rect 10502 28500 10508 28552
rect 10560 28540 10566 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 10560 28512 10609 28540
rect 10560 28500 10566 28512
rect 10597 28509 10609 28512
rect 10643 28540 10655 28543
rect 11514 28540 11520 28552
rect 10643 28512 11520 28540
rect 10643 28509 10655 28512
rect 10597 28503 10655 28509
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 11624 28512 12434 28540
rect 11624 28472 11652 28512
rect 10428 28444 11652 28472
rect 10321 28435 10379 28441
rect 11790 28432 11796 28484
rect 11848 28472 11854 28484
rect 12069 28475 12127 28481
rect 12069 28472 12081 28475
rect 11848 28444 12081 28472
rect 11848 28432 11854 28444
rect 12069 28441 12081 28444
rect 12115 28441 12127 28475
rect 12406 28472 12434 28512
rect 12526 28500 12532 28552
rect 12584 28500 12590 28552
rect 12728 28549 12756 28648
rect 13446 28636 13452 28688
rect 13504 28676 13510 28688
rect 16408 28685 16436 28716
rect 16482 28704 16488 28716
rect 16540 28704 16546 28756
rect 17678 28704 17684 28756
rect 17736 28704 17742 28756
rect 19794 28704 19800 28756
rect 19852 28704 19858 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 21560 28716 27077 28744
rect 16393 28679 16451 28685
rect 13504 28648 16344 28676
rect 13504 28636 13510 28648
rect 15013 28611 15071 28617
rect 15013 28577 15025 28611
rect 15059 28608 15071 28611
rect 16117 28611 16175 28617
rect 16117 28608 16129 28611
rect 15059 28580 16129 28608
rect 15059 28577 15071 28580
rect 15013 28571 15071 28577
rect 16117 28577 16129 28580
rect 16163 28577 16175 28611
rect 16117 28571 16175 28577
rect 16316 28552 16344 28648
rect 16393 28645 16405 28679
rect 16439 28645 16451 28679
rect 16393 28639 16451 28645
rect 16758 28636 16764 28688
rect 16816 28636 16822 28688
rect 16485 28611 16543 28617
rect 16485 28577 16497 28611
rect 16531 28608 16543 28611
rect 16776 28608 16804 28636
rect 17954 28608 17960 28620
rect 16531 28580 16804 28608
rect 17512 28580 17960 28608
rect 16531 28577 16543 28580
rect 16485 28571 16543 28577
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 14734 28500 14740 28552
rect 14792 28500 14798 28552
rect 14875 28543 14933 28549
rect 14875 28509 14887 28543
rect 14921 28540 14933 28543
rect 15102 28540 15108 28552
rect 14921 28512 15108 28540
rect 14921 28509 14933 28512
rect 14875 28503 14933 28509
rect 15102 28500 15108 28512
rect 15160 28500 15166 28552
rect 15194 28500 15200 28552
rect 15252 28500 15258 28552
rect 16298 28500 16304 28552
rect 16356 28500 16362 28552
rect 16574 28500 16580 28552
rect 16632 28500 16638 28552
rect 16761 28543 16819 28549
rect 16761 28509 16773 28543
rect 16807 28540 16819 28543
rect 16850 28540 16856 28552
rect 16807 28512 16856 28540
rect 16807 28509 16819 28512
rect 16761 28503 16819 28509
rect 16850 28500 16856 28512
rect 16908 28540 16914 28552
rect 17512 28540 17540 28580
rect 17954 28568 17960 28580
rect 18012 28568 18018 28620
rect 21450 28568 21456 28620
rect 21508 28568 21514 28620
rect 16908 28512 17540 28540
rect 17589 28543 17647 28549
rect 16908 28500 16914 28512
rect 17589 28509 17601 28543
rect 17635 28509 17647 28543
rect 17589 28503 17647 28509
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28540 17831 28543
rect 17862 28540 17868 28552
rect 17819 28512 17868 28540
rect 17819 28509 17831 28512
rect 17773 28503 17831 28509
rect 12406 28444 13308 28472
rect 12069 28435 12127 28441
rect 5810 28404 5816 28416
rect 5644 28376 5816 28404
rect 5810 28364 5816 28376
rect 5868 28404 5874 28416
rect 7374 28404 7380 28416
rect 5868 28376 7380 28404
rect 5868 28364 5874 28376
rect 7374 28364 7380 28376
rect 7432 28364 7438 28416
rect 7834 28364 7840 28416
rect 7892 28404 7898 28416
rect 9217 28407 9275 28413
rect 9217 28404 9229 28407
rect 7892 28376 9229 28404
rect 7892 28364 7898 28376
rect 9217 28373 9229 28376
rect 9263 28404 9275 28407
rect 9582 28404 9588 28416
rect 9263 28376 9588 28404
rect 9263 28373 9275 28376
rect 9217 28367 9275 28373
rect 9582 28364 9588 28376
rect 9640 28364 9646 28416
rect 10778 28364 10784 28416
rect 10836 28364 10842 28416
rect 11698 28364 11704 28416
rect 11756 28364 11762 28416
rect 11885 28407 11943 28413
rect 11885 28373 11897 28407
rect 11931 28404 11943 28407
rect 12618 28404 12624 28416
rect 11931 28376 12624 28404
rect 11931 28373 11943 28376
rect 11885 28367 11943 28373
rect 12618 28364 12624 28376
rect 12676 28364 12682 28416
rect 13280 28404 13308 28444
rect 13354 28432 13360 28484
rect 13412 28472 13418 28484
rect 17604 28472 17632 28503
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 18230 28500 18236 28552
rect 18288 28540 18294 28552
rect 19429 28543 19487 28549
rect 19429 28540 19441 28543
rect 18288 28512 19441 28540
rect 18288 28500 18294 28512
rect 19429 28509 19441 28512
rect 19475 28509 19487 28543
rect 19429 28503 19487 28509
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28540 21235 28543
rect 21358 28540 21364 28552
rect 21223 28512 21364 28540
rect 21223 28509 21235 28512
rect 21177 28503 21235 28509
rect 21358 28500 21364 28512
rect 21416 28500 21422 28552
rect 19242 28472 19248 28484
rect 13412 28444 19248 28472
rect 13412 28432 13418 28444
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 19613 28475 19671 28481
rect 19613 28441 19625 28475
rect 19659 28472 19671 28475
rect 19978 28472 19984 28484
rect 19659 28444 19984 28472
rect 19659 28441 19671 28444
rect 19613 28435 19671 28441
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 20438 28432 20444 28484
rect 20496 28472 20502 28484
rect 21560 28481 21588 28716
rect 27065 28713 27077 28716
rect 27111 28744 27123 28747
rect 27154 28744 27160 28756
rect 27111 28716 27160 28744
rect 27111 28713 27123 28716
rect 27065 28707 27123 28713
rect 27154 28704 27160 28716
rect 27212 28704 27218 28756
rect 31113 28747 31171 28753
rect 31113 28713 31125 28747
rect 31159 28744 31171 28747
rect 31294 28744 31300 28756
rect 31159 28716 31300 28744
rect 31159 28713 31171 28716
rect 31113 28707 31171 28713
rect 31294 28704 31300 28716
rect 31352 28704 31358 28756
rect 31386 28704 31392 28756
rect 31444 28744 31450 28756
rect 32309 28747 32367 28753
rect 31444 28716 32076 28744
rect 31444 28704 31450 28716
rect 23842 28676 23848 28688
rect 23400 28648 23848 28676
rect 23106 28500 23112 28552
rect 23164 28500 23170 28552
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23400 28540 23428 28648
rect 23842 28636 23848 28648
rect 23900 28636 23906 28688
rect 24946 28636 24952 28688
rect 25004 28636 25010 28688
rect 25038 28636 25044 28688
rect 25096 28636 25102 28688
rect 25133 28611 25191 28617
rect 25133 28608 25145 28611
rect 23768 28580 25145 28608
rect 23247 28512 23428 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 23474 28500 23480 28552
rect 23532 28500 23538 28552
rect 23768 28549 23796 28580
rect 25133 28577 25145 28580
rect 25179 28608 25191 28611
rect 26050 28608 26056 28620
rect 25179 28580 26056 28608
rect 25179 28577 25191 28580
rect 25133 28571 25191 28577
rect 26050 28568 26056 28580
rect 26108 28568 26114 28620
rect 27890 28608 27896 28620
rect 26160 28580 27896 28608
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28540 24087 28543
rect 24118 28540 24124 28552
rect 24075 28512 24124 28540
rect 24075 28509 24087 28512
rect 24029 28503 24087 28509
rect 24118 28500 24124 28512
rect 24176 28540 24182 28552
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 24176 28512 24593 28540
rect 24176 28500 24182 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 26160 28540 26188 28580
rect 27890 28568 27896 28580
rect 27948 28568 27954 28620
rect 31110 28608 31116 28620
rect 28368 28580 31116 28608
rect 24581 28503 24639 28509
rect 24688 28512 26188 28540
rect 21545 28475 21603 28481
rect 21545 28472 21557 28475
rect 20496 28444 21557 28472
rect 20496 28432 20502 28444
rect 21545 28441 21557 28444
rect 21591 28441 21603 28475
rect 21545 28435 21603 28441
rect 21662 28475 21720 28481
rect 21662 28441 21674 28475
rect 21708 28472 21720 28475
rect 21910 28472 21916 28484
rect 21708 28444 21916 28472
rect 21708 28441 21720 28444
rect 21662 28435 21720 28441
rect 21910 28432 21916 28444
rect 21968 28432 21974 28484
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 23290 28472 23296 28484
rect 22612 28444 23296 28472
rect 22612 28432 22618 28444
rect 23290 28432 23296 28444
rect 23348 28432 23354 28484
rect 14826 28404 14832 28416
rect 13280 28376 14832 28404
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 14918 28364 14924 28416
rect 14976 28404 14982 28416
rect 21450 28404 21456 28416
rect 14976 28376 21456 28404
rect 14976 28364 14982 28376
rect 21450 28364 21456 28376
rect 21508 28364 21514 28416
rect 21818 28364 21824 28416
rect 21876 28364 21882 28416
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 22830 28404 22836 28416
rect 22336 28376 22836 28404
rect 22336 28364 22342 28376
rect 22830 28364 22836 28376
rect 22888 28404 22894 28416
rect 24688 28404 24716 28512
rect 27062 28500 27068 28552
rect 27120 28540 27126 28552
rect 27341 28543 27399 28549
rect 27341 28540 27353 28543
rect 27120 28512 27353 28540
rect 27120 28500 27126 28512
rect 27341 28509 27353 28512
rect 27387 28509 27399 28543
rect 27341 28503 27399 28509
rect 27982 28500 27988 28552
rect 28040 28540 28046 28552
rect 28258 28540 28264 28552
rect 28040 28512 28264 28540
rect 28040 28500 28046 28512
rect 28258 28500 28264 28512
rect 28316 28500 28322 28552
rect 24762 28432 24768 28484
rect 24820 28472 24826 28484
rect 27157 28475 27215 28481
rect 24820 28444 27108 28472
rect 24820 28432 24826 28444
rect 22888 28376 24716 28404
rect 22888 28364 22894 28376
rect 25038 28364 25044 28416
rect 25096 28404 25102 28416
rect 25409 28407 25467 28413
rect 25409 28404 25421 28407
rect 25096 28376 25421 28404
rect 25096 28364 25102 28376
rect 25409 28373 25421 28376
rect 25455 28373 25467 28407
rect 27080 28404 27108 28444
rect 27157 28441 27169 28475
rect 27203 28472 27215 28475
rect 27246 28472 27252 28484
rect 27203 28444 27252 28472
rect 27203 28441 27215 28444
rect 27157 28435 27215 28441
rect 27246 28432 27252 28444
rect 27304 28472 27310 28484
rect 27430 28472 27436 28484
rect 27304 28444 27436 28472
rect 27304 28432 27310 28444
rect 27430 28432 27436 28444
rect 27488 28432 27494 28484
rect 28368 28481 28396 28580
rect 31110 28568 31116 28580
rect 31168 28568 31174 28620
rect 31312 28608 31340 28704
rect 31312 28580 31984 28608
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28540 28687 28543
rect 29914 28540 29920 28552
rect 28675 28512 29920 28540
rect 28675 28509 28687 28512
rect 28629 28503 28687 28509
rect 29914 28500 29920 28512
rect 29972 28500 29978 28552
rect 30653 28543 30711 28549
rect 30653 28509 30665 28543
rect 30699 28509 30711 28543
rect 30653 28503 30711 28509
rect 28353 28475 28411 28481
rect 28353 28472 28365 28475
rect 27540 28444 28365 28472
rect 27540 28404 27568 28444
rect 28353 28441 28365 28444
rect 28399 28441 28411 28475
rect 28353 28435 28411 28441
rect 28445 28475 28503 28481
rect 28445 28441 28457 28475
rect 28491 28441 28503 28475
rect 30668 28472 30696 28503
rect 31202 28500 31208 28552
rect 31260 28500 31266 28552
rect 31662 28500 31668 28552
rect 31720 28500 31726 28552
rect 31754 28500 31760 28552
rect 31812 28540 31818 28552
rect 31956 28549 31984 28580
rect 31941 28543 31999 28549
rect 31812 28512 31857 28540
rect 31812 28500 31818 28512
rect 31941 28509 31953 28543
rect 31987 28509 31999 28543
rect 32048 28540 32076 28716
rect 32309 28713 32321 28747
rect 32355 28744 32367 28747
rect 32398 28744 32404 28756
rect 32355 28716 32404 28744
rect 32355 28713 32367 28716
rect 32309 28707 32367 28713
rect 32398 28704 32404 28716
rect 32456 28704 32462 28756
rect 32416 28608 32444 28704
rect 35986 28676 35992 28688
rect 35820 28648 35992 28676
rect 32953 28611 33011 28617
rect 32953 28608 32965 28611
rect 32416 28580 32965 28608
rect 32953 28577 32965 28580
rect 32999 28577 33011 28611
rect 32953 28571 33011 28577
rect 33410 28568 33416 28620
rect 33468 28568 33474 28620
rect 33870 28568 33876 28620
rect 33928 28608 33934 28620
rect 35820 28608 35848 28648
rect 35986 28636 35992 28648
rect 36044 28636 36050 28688
rect 33928 28580 35848 28608
rect 33928 28568 33934 28580
rect 32130 28543 32188 28549
rect 32130 28540 32142 28543
rect 32048 28512 32142 28540
rect 31941 28503 31999 28509
rect 32130 28509 32142 28512
rect 32176 28509 32188 28543
rect 32130 28503 32188 28509
rect 33042 28500 33048 28552
rect 33100 28500 33106 28552
rect 35526 28500 35532 28552
rect 35584 28500 35590 28552
rect 35820 28549 35848 28580
rect 36354 28568 36360 28620
rect 36412 28608 36418 28620
rect 36633 28611 36691 28617
rect 36633 28608 36645 28611
rect 36412 28580 36645 28608
rect 36412 28568 36418 28580
rect 36633 28577 36645 28580
rect 36679 28577 36691 28611
rect 36633 28571 36691 28577
rect 35622 28543 35680 28549
rect 35622 28509 35634 28543
rect 35668 28509 35680 28543
rect 35622 28503 35680 28509
rect 35805 28543 35863 28549
rect 35805 28509 35817 28543
rect 35851 28509 35863 28543
rect 35805 28503 35863 28509
rect 31386 28472 31392 28484
rect 30668 28444 31392 28472
rect 28445 28435 28503 28441
rect 27080 28376 27568 28404
rect 25409 28367 25467 28373
rect 27614 28364 27620 28416
rect 27672 28404 27678 28416
rect 28077 28407 28135 28413
rect 28077 28404 28089 28407
rect 27672 28376 28089 28404
rect 27672 28364 27678 28376
rect 28077 28373 28089 28376
rect 28123 28373 28135 28407
rect 28460 28404 28488 28435
rect 31386 28432 31392 28444
rect 31444 28432 31450 28484
rect 32030 28432 32036 28484
rect 32088 28432 32094 28484
rect 28626 28404 28632 28416
rect 28460 28376 28632 28404
rect 28077 28367 28135 28373
rect 28626 28364 28632 28376
rect 28684 28364 28690 28416
rect 29914 28364 29920 28416
rect 29972 28404 29978 28416
rect 35636 28404 35664 28503
rect 35894 28500 35900 28552
rect 35952 28500 35958 28552
rect 36035 28543 36093 28549
rect 36035 28509 36047 28543
rect 36081 28540 36093 28543
rect 36262 28540 36268 28552
rect 36081 28512 36268 28540
rect 36081 28509 36093 28512
rect 36035 28503 36093 28509
rect 36262 28500 36268 28512
rect 36320 28500 36326 28552
rect 36900 28475 36958 28481
rect 36004 28444 36308 28472
rect 36004 28404 36032 28444
rect 29972 28376 36032 28404
rect 29972 28364 29978 28376
rect 36170 28364 36176 28416
rect 36228 28364 36234 28416
rect 36280 28404 36308 28444
rect 36900 28441 36912 28475
rect 36946 28472 36958 28475
rect 37458 28472 37464 28484
rect 36946 28444 37464 28472
rect 36946 28441 36958 28444
rect 36900 28435 36958 28441
rect 37458 28432 37464 28444
rect 37516 28432 37522 28484
rect 37826 28404 37832 28416
rect 36280 28376 37832 28404
rect 37826 28364 37832 28376
rect 37884 28404 37890 28416
rect 38013 28407 38071 28413
rect 38013 28404 38025 28407
rect 37884 28376 38025 28404
rect 37884 28364 37890 28376
rect 38013 28373 38025 28376
rect 38059 28373 38071 28407
rect 38013 28367 38071 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 4798 28160 4804 28212
rect 4856 28200 4862 28212
rect 11698 28200 11704 28212
rect 4856 28172 11704 28200
rect 4856 28160 4862 28172
rect 3878 27956 3884 28008
rect 3936 27996 3942 28008
rect 4908 27996 4936 28172
rect 11698 28160 11704 28172
rect 11756 28160 11762 28212
rect 11790 28160 11796 28212
rect 11848 28200 11854 28212
rect 11848 28172 13492 28200
rect 11848 28160 11854 28172
rect 6546 28132 6552 28144
rect 5000 28104 6552 28132
rect 5000 28073 5028 28104
rect 6546 28092 6552 28104
rect 6604 28092 6610 28144
rect 6825 28135 6883 28141
rect 6825 28101 6837 28135
rect 6871 28132 6883 28135
rect 7190 28132 7196 28144
rect 6871 28104 7196 28132
rect 6871 28101 6883 28104
rect 6825 28095 6883 28101
rect 7190 28092 7196 28104
rect 7248 28092 7254 28144
rect 10778 28092 10784 28144
rect 10836 28132 10842 28144
rect 13354 28132 13360 28144
rect 10836 28104 13360 28132
rect 10836 28092 10842 28104
rect 13354 28092 13360 28104
rect 13412 28092 13418 28144
rect 13464 28132 13492 28172
rect 14642 28160 14648 28212
rect 14700 28160 14706 28212
rect 16942 28160 16948 28212
rect 17000 28160 17006 28212
rect 20162 28160 20168 28212
rect 20220 28200 20226 28212
rect 20220 28172 20484 28200
rect 20220 28160 20226 28172
rect 13464 28104 20392 28132
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28033 5043 28067
rect 4985 28027 5043 28033
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28033 5135 28067
rect 5077 28027 5135 28033
rect 5092 27996 5120 28027
rect 5166 28024 5172 28076
rect 5224 28024 5230 28076
rect 5353 28067 5411 28073
rect 5353 28033 5365 28067
rect 5399 28064 5411 28067
rect 5534 28064 5540 28076
rect 5399 28036 5540 28064
rect 5399 28033 5411 28036
rect 5353 28027 5411 28033
rect 5534 28024 5540 28036
rect 5592 28024 5598 28076
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 9309 28067 9367 28073
rect 9309 28064 9321 28067
rect 9272 28036 9321 28064
rect 9272 28024 9278 28036
rect 9309 28033 9321 28036
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 9493 28067 9551 28073
rect 9493 28033 9505 28067
rect 9539 28064 9551 28067
rect 10042 28064 10048 28076
rect 9539 28036 10048 28064
rect 9539 28033 9551 28036
rect 9493 28027 9551 28033
rect 10042 28024 10048 28036
rect 10100 28024 10106 28076
rect 10134 28024 10140 28076
rect 10192 28064 10198 28076
rect 10229 28067 10287 28073
rect 10229 28064 10241 28067
rect 10192 28036 10241 28064
rect 10192 28024 10198 28036
rect 10229 28033 10241 28036
rect 10275 28033 10287 28067
rect 10229 28027 10287 28033
rect 10502 28024 10508 28076
rect 10560 28024 10566 28076
rect 12618 28024 12624 28076
rect 12676 28024 12682 28076
rect 13464 28073 13492 28104
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28033 13507 28067
rect 13449 28027 13507 28033
rect 14093 28067 14151 28073
rect 14093 28033 14105 28067
rect 14139 28033 14151 28067
rect 14093 28027 14151 28033
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 16482 28064 16488 28076
rect 14507 28036 16488 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 3936 27968 5120 27996
rect 3936 27956 3942 27968
rect 5184 27928 5212 28024
rect 7098 27956 7104 28008
rect 7156 27996 7162 28008
rect 7193 27999 7251 28005
rect 7193 27996 7205 27999
rect 7156 27968 7205 27996
rect 7156 27956 7162 27968
rect 7193 27965 7205 27968
rect 7239 27965 7251 27999
rect 7193 27959 7251 27965
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27996 10471 27999
rect 10594 27996 10600 28008
rect 10459 27968 10600 27996
rect 10459 27965 10471 27968
rect 10413 27959 10471 27965
rect 10594 27956 10600 27968
rect 10652 27956 10658 28008
rect 13354 27956 13360 28008
rect 13412 27956 13418 28008
rect 7742 27928 7748 27940
rect 5184 27900 7748 27928
rect 7742 27888 7748 27900
rect 7800 27888 7806 27940
rect 8294 27888 8300 27940
rect 8352 27928 8358 27940
rect 10689 27931 10747 27937
rect 8352 27900 10272 27928
rect 8352 27888 8358 27900
rect 4798 27820 4804 27872
rect 4856 27820 4862 27872
rect 6546 27820 6552 27872
rect 6604 27860 6610 27872
rect 6641 27863 6699 27869
rect 6641 27860 6653 27863
rect 6604 27832 6653 27860
rect 6604 27820 6610 27832
rect 6641 27829 6653 27832
rect 6687 27829 6699 27863
rect 6641 27823 6699 27829
rect 6822 27820 6828 27872
rect 6880 27820 6886 27872
rect 9214 27820 9220 27872
rect 9272 27860 9278 27872
rect 10244 27869 10272 27900
rect 10689 27897 10701 27931
rect 10735 27928 10747 27931
rect 14108 27928 14136 28027
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 16850 28024 16856 28076
rect 16908 28024 16914 28076
rect 17037 28067 17095 28073
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 18322 28064 18328 28076
rect 17083 28036 18328 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 16574 27956 16580 28008
rect 16632 27996 16638 28008
rect 17052 27996 17080 28027
rect 18322 28024 18328 28036
rect 18380 28064 18386 28076
rect 19978 28064 19984 28076
rect 18380 28036 19984 28064
rect 18380 28024 18386 28036
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 20162 28024 20168 28076
rect 20220 28024 20226 28076
rect 16632 27968 17080 27996
rect 16632 27956 16638 27968
rect 20254 27956 20260 28008
rect 20312 27956 20318 28008
rect 20364 27996 20392 28104
rect 20456 28064 20484 28172
rect 20990 28160 20996 28212
rect 21048 28200 21054 28212
rect 24762 28200 24768 28212
rect 21048 28172 24768 28200
rect 21048 28160 21054 28172
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 24854 28160 24860 28212
rect 24912 28200 24918 28212
rect 25958 28200 25964 28212
rect 24912 28172 25964 28200
rect 24912 28160 24918 28172
rect 25958 28160 25964 28172
rect 26016 28160 26022 28212
rect 27890 28160 27896 28212
rect 27948 28200 27954 28212
rect 28537 28203 28595 28209
rect 28537 28200 28549 28203
rect 27948 28172 28549 28200
rect 27948 28160 27954 28172
rect 28537 28169 28549 28172
rect 28583 28200 28595 28203
rect 28626 28200 28632 28212
rect 28583 28172 28632 28200
rect 28583 28169 28595 28172
rect 28537 28163 28595 28169
rect 28626 28160 28632 28172
rect 28684 28160 28690 28212
rect 30374 28160 30380 28212
rect 30432 28160 30438 28212
rect 31754 28200 31760 28212
rect 30484 28172 31760 28200
rect 20530 28092 20536 28144
rect 20588 28132 20594 28144
rect 20588 28104 22416 28132
rect 20588 28092 20594 28104
rect 22278 28064 22284 28076
rect 20456 28036 22284 28064
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22388 28073 22416 28104
rect 22830 28092 22836 28144
rect 22888 28132 22894 28144
rect 23290 28132 23296 28144
rect 22888 28104 23296 28132
rect 22888 28092 22894 28104
rect 23290 28092 23296 28104
rect 23348 28092 23354 28144
rect 24118 28092 24124 28144
rect 24176 28132 24182 28144
rect 25130 28132 25136 28144
rect 24176 28104 25136 28132
rect 24176 28092 24182 28104
rect 25130 28092 25136 28104
rect 25188 28092 25194 28144
rect 25424 28104 27476 28132
rect 25424 28076 25452 28104
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28033 22431 28067
rect 22373 28027 22431 28033
rect 22649 28067 22707 28073
rect 22649 28033 22661 28067
rect 22695 28064 22707 28067
rect 23106 28064 23112 28076
rect 22695 28036 23112 28064
rect 22695 28033 22707 28036
rect 22649 28027 22707 28033
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 23198 28024 23204 28076
rect 23256 28024 23262 28076
rect 24029 28067 24087 28073
rect 24029 28033 24041 28067
rect 24075 28064 24087 28067
rect 25038 28064 25044 28076
rect 24075 28036 25044 28064
rect 24075 28033 24087 28036
rect 24029 28027 24087 28033
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25406 28024 25412 28076
rect 25464 28024 25470 28076
rect 25961 28067 26019 28073
rect 25961 28033 25973 28067
rect 26007 28033 26019 28067
rect 25961 28027 26019 28033
rect 24946 27996 24952 28008
rect 20364 27968 24952 27996
rect 24946 27956 24952 27968
rect 25004 27956 25010 28008
rect 25222 27956 25228 28008
rect 25280 27996 25286 28008
rect 25976 27996 26004 28027
rect 26234 28024 26240 28076
rect 26292 28024 26298 28076
rect 27338 28024 27344 28076
rect 27396 28024 27402 28076
rect 27448 28064 27476 28104
rect 27798 28092 27804 28144
rect 27856 28092 27862 28144
rect 30006 28092 30012 28144
rect 30064 28092 30070 28144
rect 28353 28067 28411 28073
rect 28353 28064 28365 28067
rect 27448 28036 28365 28064
rect 28353 28033 28365 28036
rect 28399 28033 28411 28067
rect 28353 28027 28411 28033
rect 29730 28024 29736 28076
rect 29788 28024 29794 28076
rect 30282 28073 30288 28076
rect 29826 28067 29884 28073
rect 29826 28033 29838 28067
rect 29872 28033 29884 28067
rect 29826 28027 29884 28033
rect 30101 28067 30159 28073
rect 30101 28033 30113 28067
rect 30147 28033 30159 28067
rect 30101 28027 30159 28033
rect 30239 28067 30288 28073
rect 30239 28033 30251 28067
rect 30285 28033 30288 28067
rect 30239 28027 30288 28033
rect 25280 27968 26004 27996
rect 25280 27956 25286 27968
rect 27430 27956 27436 28008
rect 27488 27956 27494 28008
rect 29546 27956 29552 28008
rect 29604 27996 29610 28008
rect 29840 27996 29868 28027
rect 29604 27968 29868 27996
rect 30116 27996 30144 28027
rect 30282 28024 30288 28027
rect 30340 28024 30346 28076
rect 30374 27996 30380 28008
rect 30116 27968 30380 27996
rect 29604 27956 29610 27968
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 10735 27900 14136 27928
rect 10735 27897 10747 27900
rect 10689 27891 10747 27897
rect 14826 27888 14832 27940
rect 14884 27928 14890 27940
rect 19334 27928 19340 27940
rect 14884 27900 19340 27928
rect 14884 27888 14890 27900
rect 19334 27888 19340 27900
rect 19392 27888 19398 27940
rect 19978 27888 19984 27940
rect 20036 27928 20042 27940
rect 22373 27931 22431 27937
rect 20036 27900 22094 27928
rect 20036 27888 20042 27900
rect 9401 27863 9459 27869
rect 9401 27860 9413 27863
rect 9272 27832 9413 27860
rect 9272 27820 9278 27832
rect 9401 27829 9413 27832
rect 9447 27829 9459 27863
rect 9401 27823 9459 27829
rect 10229 27863 10287 27869
rect 10229 27829 10241 27863
rect 10275 27829 10287 27863
rect 10229 27823 10287 27829
rect 13170 27820 13176 27872
rect 13228 27860 13234 27872
rect 14185 27863 14243 27869
rect 14185 27860 14197 27863
rect 13228 27832 14197 27860
rect 13228 27820 13234 27832
rect 14185 27829 14197 27832
rect 14231 27829 14243 27863
rect 14185 27823 14243 27829
rect 20070 27820 20076 27872
rect 20128 27860 20134 27872
rect 20165 27863 20223 27869
rect 20165 27860 20177 27863
rect 20128 27832 20177 27860
rect 20128 27820 20134 27832
rect 20165 27829 20177 27832
rect 20211 27829 20223 27863
rect 20165 27823 20223 27829
rect 20530 27820 20536 27872
rect 20588 27820 20594 27872
rect 22066 27860 22094 27900
rect 22373 27897 22385 27931
rect 22419 27928 22431 27931
rect 22830 27928 22836 27940
rect 22419 27900 22836 27928
rect 22419 27897 22431 27900
rect 22373 27891 22431 27897
rect 22830 27888 22836 27900
rect 22888 27888 22894 27940
rect 24489 27931 24547 27937
rect 24489 27928 24501 27931
rect 23308 27900 24501 27928
rect 23308 27860 23336 27900
rect 24489 27897 24501 27900
rect 24535 27928 24547 27931
rect 26970 27928 26976 27940
rect 24535 27900 26976 27928
rect 24535 27897 24547 27900
rect 24489 27891 24547 27897
rect 26970 27888 26976 27900
rect 27028 27888 27034 27940
rect 27062 27888 27068 27940
rect 27120 27928 27126 27940
rect 30484 27928 30512 28172
rect 31754 28160 31760 28172
rect 31812 28200 31818 28212
rect 34238 28200 34244 28212
rect 31812 28172 32260 28200
rect 31812 28160 31818 28172
rect 31021 28135 31079 28141
rect 31021 28101 31033 28135
rect 31067 28132 31079 28135
rect 31846 28132 31852 28144
rect 31067 28104 31852 28132
rect 31067 28101 31079 28104
rect 31021 28095 31079 28101
rect 31846 28092 31852 28104
rect 31904 28092 31910 28144
rect 31757 28067 31815 28073
rect 31757 28033 31769 28067
rect 31803 28033 31815 28067
rect 31757 28027 31815 28033
rect 27120 27900 30512 27928
rect 31772 27928 31800 28027
rect 32232 27996 32260 28172
rect 32692 28172 34244 28200
rect 32306 28024 32312 28076
rect 32364 28024 32370 28076
rect 32398 28024 32404 28076
rect 32456 28024 32462 28076
rect 32692 28073 32720 28172
rect 34238 28160 34244 28172
rect 34296 28160 34302 28212
rect 37458 28160 37464 28212
rect 37516 28160 37522 28212
rect 37826 28160 37832 28212
rect 37884 28160 37890 28212
rect 33410 28092 33416 28144
rect 33468 28132 33474 28144
rect 34394 28135 34452 28141
rect 34394 28132 34406 28135
rect 33468 28104 34406 28132
rect 33468 28092 33474 28104
rect 34394 28101 34406 28104
rect 34440 28101 34452 28135
rect 34394 28095 34452 28101
rect 36170 28092 36176 28144
rect 36228 28132 36234 28144
rect 37921 28135 37979 28141
rect 37921 28132 37933 28135
rect 36228 28104 37933 28132
rect 36228 28092 36234 28104
rect 37921 28101 37933 28104
rect 37967 28101 37979 28135
rect 37921 28095 37979 28101
rect 32585 28067 32643 28073
rect 32585 28033 32597 28067
rect 32631 28033 32643 28067
rect 32585 28027 32643 28033
rect 32677 28067 32735 28073
rect 32677 28033 32689 28067
rect 32723 28033 32735 28067
rect 32677 28027 32735 28033
rect 32861 28067 32919 28073
rect 32861 28033 32873 28067
rect 32907 28064 32919 28067
rect 33594 28064 33600 28076
rect 32907 28036 33600 28064
rect 32907 28033 32919 28036
rect 32861 28027 32919 28033
rect 32600 27996 32628 28027
rect 33594 28024 33600 28036
rect 33652 28024 33658 28076
rect 32232 27968 32720 27996
rect 32582 27928 32588 27940
rect 31772 27900 32588 27928
rect 27120 27888 27126 27900
rect 32582 27888 32588 27900
rect 32640 27888 32646 27940
rect 22066 27832 23336 27860
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 23474 27860 23480 27872
rect 23431 27832 23480 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 23474 27820 23480 27832
rect 23532 27860 23538 27872
rect 26418 27860 26424 27872
rect 23532 27832 26424 27860
rect 23532 27820 23538 27832
rect 26418 27820 26424 27832
rect 26476 27820 26482 27872
rect 27154 27820 27160 27872
rect 27212 27820 27218 27872
rect 27522 27820 27528 27872
rect 27580 27820 27586 27872
rect 32692 27860 32720 27968
rect 33318 27956 33324 28008
rect 33376 27996 33382 28008
rect 34149 27999 34207 28005
rect 34149 27996 34161 27999
rect 33376 27968 34161 27996
rect 33376 27956 33382 27968
rect 34149 27965 34161 27968
rect 34195 27965 34207 27999
rect 34149 27959 34207 27965
rect 38010 27956 38016 28008
rect 38068 27956 38074 28008
rect 35529 27863 35587 27869
rect 35529 27860 35541 27863
rect 32692 27832 35541 27860
rect 35529 27829 35541 27832
rect 35575 27829 35587 27863
rect 35529 27823 35587 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 18693 27659 18751 27665
rect 4540 27628 4752 27656
rect 4249 27591 4307 27597
rect 4249 27557 4261 27591
rect 4295 27588 4307 27591
rect 4540 27588 4568 27628
rect 4295 27560 4568 27588
rect 4295 27557 4307 27560
rect 4249 27551 4307 27557
rect 4614 27548 4620 27600
rect 4672 27548 4678 27600
rect 4724 27588 4752 27628
rect 18693 27625 18705 27659
rect 18739 27625 18751 27659
rect 18693 27619 18751 27625
rect 5626 27588 5632 27600
rect 4724 27560 5632 27588
rect 5626 27548 5632 27560
rect 5684 27548 5690 27600
rect 7190 27548 7196 27600
rect 7248 27588 7254 27600
rect 7466 27588 7472 27600
rect 7248 27560 7472 27588
rect 7248 27548 7254 27560
rect 4341 27523 4399 27529
rect 4341 27489 4353 27523
rect 4387 27520 4399 27523
rect 4632 27520 4660 27548
rect 4387 27492 4660 27520
rect 4387 27489 4399 27492
rect 4341 27483 4399 27489
rect 5350 27480 5356 27532
rect 5408 27480 5414 27532
rect 7300 27529 7328 27560
rect 7466 27548 7472 27560
rect 7524 27588 7530 27600
rect 7524 27560 8156 27588
rect 7524 27548 7530 27560
rect 7285 27523 7343 27529
rect 7285 27489 7297 27523
rect 7331 27489 7343 27523
rect 7285 27483 7343 27489
rect 7742 27480 7748 27532
rect 7800 27520 7806 27532
rect 7921 27523 7979 27529
rect 7921 27520 7933 27523
rect 7800 27492 7933 27520
rect 7800 27480 7806 27492
rect 7921 27489 7933 27492
rect 7967 27489 7979 27523
rect 7921 27483 7979 27489
rect 8128 27520 8156 27560
rect 9122 27548 9128 27600
rect 9180 27548 9186 27600
rect 10686 27548 10692 27600
rect 10744 27548 10750 27600
rect 16945 27591 17003 27597
rect 16945 27557 16957 27591
rect 16991 27588 17003 27591
rect 17034 27588 17040 27600
rect 16991 27560 17040 27588
rect 16991 27557 17003 27560
rect 16945 27551 17003 27557
rect 17034 27548 17040 27560
rect 17092 27588 17098 27600
rect 17678 27588 17684 27600
rect 17092 27560 17684 27588
rect 17092 27548 17098 27560
rect 17678 27548 17684 27560
rect 17736 27548 17742 27600
rect 18230 27548 18236 27600
rect 18288 27588 18294 27600
rect 18509 27591 18567 27597
rect 18509 27588 18521 27591
rect 18288 27560 18521 27588
rect 18288 27548 18294 27560
rect 18509 27557 18521 27560
rect 18555 27557 18567 27591
rect 18708 27588 18736 27619
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 20990 27656 20996 27668
rect 19392 27628 20996 27656
rect 19392 27616 19398 27628
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 21174 27616 21180 27668
rect 21232 27656 21238 27668
rect 23658 27656 23664 27668
rect 21232 27628 23664 27656
rect 21232 27616 21238 27628
rect 23658 27616 23664 27628
rect 23716 27616 23722 27668
rect 29730 27616 29736 27668
rect 29788 27656 29794 27668
rect 30926 27656 30932 27668
rect 29788 27628 30932 27656
rect 29788 27616 29794 27628
rect 30926 27616 30932 27628
rect 30984 27616 30990 27668
rect 31110 27616 31116 27668
rect 31168 27616 31174 27668
rect 31202 27616 31208 27668
rect 31260 27656 31266 27668
rect 31481 27659 31539 27665
rect 31481 27656 31493 27659
rect 31260 27628 31493 27656
rect 31260 27616 31266 27628
rect 31481 27625 31493 27628
rect 31527 27625 31539 27659
rect 31481 27619 31539 27625
rect 32306 27616 32312 27668
rect 32364 27656 32370 27668
rect 32364 27628 33548 27656
rect 32364 27616 32370 27628
rect 18708 27560 19472 27588
rect 18509 27551 18567 27557
rect 9140 27520 9168 27548
rect 10226 27520 10232 27532
rect 8128 27492 9168 27520
rect 9324 27492 10232 27520
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27421 4215 27455
rect 4157 27415 4215 27421
rect 4172 27384 4200 27415
rect 4430 27412 4436 27464
rect 4488 27412 4494 27464
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27452 4675 27455
rect 4663 27424 5028 27452
rect 4663 27421 4675 27424
rect 4617 27415 4675 27421
rect 4798 27384 4804 27396
rect 4172 27356 4804 27384
rect 4798 27344 4804 27356
rect 4856 27344 4862 27396
rect 5000 27384 5028 27424
rect 5074 27412 5080 27464
rect 5132 27412 5138 27464
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 5276 27384 5304 27415
rect 5442 27412 5448 27464
rect 5500 27412 5506 27464
rect 5629 27455 5687 27461
rect 5629 27421 5641 27455
rect 5675 27452 5687 27455
rect 5718 27452 5724 27464
rect 5675 27424 5724 27452
rect 5675 27421 5687 27424
rect 5629 27415 5687 27421
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 7098 27412 7104 27464
rect 7156 27452 7162 27464
rect 7834 27452 7840 27464
rect 7156 27424 7840 27452
rect 7156 27412 7162 27424
rect 7834 27412 7840 27424
rect 7892 27452 7898 27464
rect 8128 27461 8156 27492
rect 8010 27455 8068 27461
rect 8010 27452 8022 27455
rect 7892 27424 8022 27452
rect 7892 27412 7898 27424
rect 8010 27421 8022 27424
rect 8056 27421 8068 27455
rect 8010 27415 8068 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8113 27415 8171 27421
rect 8205 27455 8263 27461
rect 8205 27421 8217 27455
rect 8251 27421 8263 27455
rect 8205 27415 8263 27421
rect 6178 27384 6184 27396
rect 5000 27356 5120 27384
rect 5276 27356 6184 27384
rect 5092 27328 5120 27356
rect 6178 27344 6184 27356
rect 6236 27344 6242 27396
rect 6270 27344 6276 27396
rect 6328 27384 6334 27396
rect 8220 27384 8248 27415
rect 8294 27412 8300 27464
rect 8352 27452 8358 27464
rect 9324 27461 9352 27492
rect 10226 27480 10232 27492
rect 10284 27520 10290 27532
rect 10704 27520 10732 27548
rect 10284 27492 10732 27520
rect 16853 27523 16911 27529
rect 10284 27480 10290 27492
rect 16853 27489 16865 27523
rect 16899 27520 16911 27523
rect 17954 27520 17960 27532
rect 16899 27492 17960 27520
rect 16899 27489 16911 27492
rect 16853 27483 16911 27489
rect 17954 27480 17960 27492
rect 18012 27520 18018 27532
rect 18598 27520 18604 27532
rect 18012 27492 18604 27520
rect 18012 27480 18018 27492
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 19444 27529 19472 27560
rect 21560 27560 22876 27588
rect 18693 27523 18751 27529
rect 18693 27489 18705 27523
rect 18739 27489 18751 27523
rect 18693 27483 18751 27489
rect 18785 27523 18843 27529
rect 18785 27489 18797 27523
rect 18831 27520 18843 27523
rect 19429 27523 19487 27529
rect 18831 27492 19380 27520
rect 18831 27489 18843 27492
rect 18785 27483 18843 27489
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 8352 27424 9137 27452
rect 8352 27412 8358 27424
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27452 10563 27455
rect 10778 27452 10784 27464
rect 10551 27424 10784 27452
rect 10551 27421 10563 27424
rect 10505 27415 10563 27421
rect 10778 27412 10784 27424
rect 10836 27452 10842 27464
rect 11882 27452 11888 27464
rect 10836 27424 11888 27452
rect 10836 27412 10842 27424
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 12342 27412 12348 27464
rect 12400 27412 12406 27464
rect 16761 27455 16819 27461
rect 16761 27421 16773 27455
rect 16807 27421 16819 27455
rect 16761 27415 16819 27421
rect 17037 27455 17095 27461
rect 17037 27421 17049 27455
rect 17083 27452 17095 27455
rect 17126 27452 17132 27464
rect 17083 27424 17132 27452
rect 17083 27421 17095 27424
rect 17037 27415 17095 27421
rect 6328 27356 8156 27384
rect 8220 27356 9260 27384
rect 6328 27344 6334 27356
rect 3970 27276 3976 27328
rect 4028 27276 4034 27328
rect 5074 27276 5080 27328
rect 5132 27276 5138 27328
rect 5534 27276 5540 27328
rect 5592 27316 5598 27328
rect 5813 27319 5871 27325
rect 5813 27316 5825 27319
rect 5592 27288 5825 27316
rect 5592 27276 5598 27288
rect 5813 27285 5825 27288
rect 5859 27285 5871 27319
rect 5813 27279 5871 27285
rect 5902 27276 5908 27328
rect 5960 27316 5966 27328
rect 6917 27319 6975 27325
rect 6917 27316 6929 27319
rect 5960 27288 6929 27316
rect 5960 27276 5966 27288
rect 6917 27285 6929 27288
rect 6963 27285 6975 27319
rect 6917 27279 6975 27285
rect 7742 27276 7748 27328
rect 7800 27276 7806 27328
rect 8128 27316 8156 27356
rect 9030 27316 9036 27328
rect 8128 27288 9036 27316
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 9232 27325 9260 27356
rect 10318 27344 10324 27396
rect 10376 27344 10382 27396
rect 12612 27387 12670 27393
rect 12612 27353 12624 27387
rect 12658 27384 12670 27387
rect 12802 27384 12808 27396
rect 12658 27356 12808 27384
rect 12658 27353 12670 27356
rect 12612 27347 12670 27353
rect 12802 27344 12808 27356
rect 12860 27344 12866 27396
rect 16776 27384 16804 27415
rect 17126 27412 17132 27424
rect 17184 27412 17190 27464
rect 16776 27356 17080 27384
rect 17052 27328 17080 27356
rect 17402 27344 17408 27396
rect 17460 27384 17466 27396
rect 18708 27384 18736 27483
rect 18877 27455 18935 27461
rect 18877 27421 18889 27455
rect 18923 27452 18935 27455
rect 19058 27452 19064 27464
rect 18923 27424 19064 27452
rect 18923 27421 18935 27424
rect 18877 27415 18935 27421
rect 19058 27412 19064 27424
rect 19116 27412 19122 27464
rect 19352 27452 19380 27492
rect 19429 27489 19441 27523
rect 19475 27489 19487 27523
rect 20438 27520 20444 27532
rect 19429 27483 19487 27489
rect 19996 27492 20444 27520
rect 19996 27452 20024 27492
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 19352 27424 20024 27452
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 21560 27461 21588 27560
rect 22848 27520 22876 27560
rect 22922 27548 22928 27600
rect 22980 27588 22986 27600
rect 23198 27588 23204 27600
rect 22980 27560 23204 27588
rect 22980 27548 22986 27560
rect 23198 27548 23204 27560
rect 23256 27548 23262 27600
rect 23566 27548 23572 27600
rect 23624 27548 23630 27600
rect 23753 27591 23811 27597
rect 23753 27557 23765 27591
rect 23799 27588 23811 27591
rect 24118 27588 24124 27600
rect 23799 27560 24124 27588
rect 23799 27557 23811 27560
rect 23753 27551 23811 27557
rect 24118 27548 24124 27560
rect 24176 27548 24182 27600
rect 27798 27548 27804 27600
rect 27856 27548 27862 27600
rect 23474 27520 23480 27532
rect 22848 27492 23480 27520
rect 23474 27480 23480 27492
rect 23532 27480 23538 27532
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 25774 27520 25780 27532
rect 24912 27492 25780 27520
rect 24912 27480 24918 27492
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 26973 27523 27031 27529
rect 26344 27492 26832 27520
rect 20165 27455 20223 27461
rect 20165 27452 20177 27455
rect 20128 27424 20177 27452
rect 20128 27412 20134 27424
rect 20165 27421 20177 27424
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 21818 27412 21824 27464
rect 21876 27452 21882 27464
rect 22189 27455 22247 27461
rect 22189 27452 22201 27455
rect 21876 27424 22201 27452
rect 21876 27412 21882 27424
rect 22189 27421 22201 27424
rect 22235 27421 22247 27455
rect 22189 27415 22247 27421
rect 22646 27412 22652 27464
rect 22704 27412 22710 27464
rect 25314 27452 25320 27464
rect 23860 27424 25320 27452
rect 19981 27387 20039 27393
rect 17460 27356 19932 27384
rect 17460 27344 17466 27356
rect 19904 27328 19932 27356
rect 19981 27353 19993 27387
rect 20027 27384 20039 27387
rect 20714 27384 20720 27396
rect 20027 27356 20720 27384
rect 20027 27353 20039 27356
rect 19981 27347 20039 27353
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 21082 27344 21088 27396
rect 21140 27344 21146 27396
rect 23860 27384 23888 27424
rect 25314 27412 25320 27424
rect 25372 27452 25378 27464
rect 26142 27452 26148 27464
rect 25372 27424 26148 27452
rect 25372 27412 25378 27424
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 26344 27461 26372 27492
rect 26329 27455 26387 27461
rect 26329 27421 26341 27455
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 22066 27356 23888 27384
rect 9217 27319 9275 27325
rect 9217 27285 9229 27319
rect 9263 27316 9275 27319
rect 9858 27316 9864 27328
rect 9263 27288 9864 27316
rect 9263 27285 9275 27288
rect 9217 27279 9275 27285
rect 9858 27276 9864 27288
rect 9916 27276 9922 27328
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 13446 27316 13452 27328
rect 12492 27288 13452 27316
rect 12492 27276 12498 27288
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 13725 27319 13783 27325
rect 13725 27285 13737 27319
rect 13771 27316 13783 27319
rect 13998 27316 14004 27328
rect 13771 27288 14004 27316
rect 13771 27285 13783 27288
rect 13725 27279 13783 27285
rect 13998 27276 14004 27288
rect 14056 27276 14062 27328
rect 16574 27276 16580 27328
rect 16632 27276 16638 27328
rect 17034 27276 17040 27328
rect 17092 27276 17098 27328
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 19392 27288 19625 27316
rect 19392 27276 19398 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19613 27279 19671 27285
rect 19886 27276 19892 27328
rect 19944 27276 19950 27328
rect 20073 27319 20131 27325
rect 20073 27285 20085 27319
rect 20119 27316 20131 27319
rect 22066 27316 22094 27356
rect 23934 27344 23940 27396
rect 23992 27384 23998 27396
rect 24029 27387 24087 27393
rect 24029 27384 24041 27387
rect 23992 27356 24041 27384
rect 23992 27344 23998 27356
rect 24029 27353 24041 27356
rect 24075 27353 24087 27387
rect 25225 27387 25283 27393
rect 25225 27384 25237 27387
rect 24029 27347 24087 27353
rect 24872 27356 25237 27384
rect 20119 27288 22094 27316
rect 22373 27319 22431 27325
rect 20119 27285 20131 27288
rect 20073 27279 20131 27285
rect 22373 27285 22385 27319
rect 22419 27316 22431 27319
rect 22462 27316 22468 27328
rect 22419 27288 22468 27316
rect 22419 27285 22431 27288
rect 22373 27279 22431 27285
rect 22462 27276 22468 27288
rect 22520 27276 22526 27328
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 24762 27316 24768 27328
rect 23164 27288 24768 27316
rect 23164 27276 23170 27288
rect 24762 27276 24768 27288
rect 24820 27316 24826 27328
rect 24872 27316 24900 27356
rect 25225 27353 25237 27356
rect 25271 27353 25283 27387
rect 25225 27347 25283 27353
rect 24820 27288 24900 27316
rect 25041 27319 25099 27325
rect 24820 27276 24826 27288
rect 25041 27285 25053 27319
rect 25087 27316 25099 27319
rect 25130 27316 25136 27328
rect 25087 27288 25136 27316
rect 25087 27285 25099 27288
rect 25041 27279 25099 27285
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 25240 27316 25268 27347
rect 25406 27344 25412 27396
rect 25464 27344 25470 27396
rect 25498 27344 25504 27396
rect 25556 27384 25562 27396
rect 26528 27384 26556 27415
rect 26602 27412 26608 27464
rect 26660 27412 26666 27464
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27421 26755 27455
rect 26804 27452 26832 27492
rect 26973 27489 26985 27523
rect 27019 27520 27031 27523
rect 27816 27520 27844 27548
rect 27019 27492 27476 27520
rect 27019 27489 27031 27492
rect 26973 27483 27031 27489
rect 27338 27452 27344 27464
rect 26804 27424 27344 27452
rect 26697 27415 26755 27421
rect 25556 27356 26556 27384
rect 25556 27344 25562 27356
rect 26234 27316 26240 27328
rect 25240 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27316 26298 27328
rect 26712 27316 26740 27415
rect 27338 27412 27344 27424
rect 27396 27412 27402 27464
rect 27448 27461 27476 27492
rect 27632 27492 27844 27520
rect 27632 27461 27660 27492
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 27617 27455 27675 27461
rect 27617 27421 27629 27455
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 27706 27412 27712 27464
rect 27764 27412 27770 27464
rect 27801 27455 27859 27461
rect 27801 27421 27813 27455
rect 27847 27421 27859 27455
rect 29748 27452 29776 27616
rect 30282 27548 30288 27600
rect 30340 27548 30346 27600
rect 30469 27591 30527 27597
rect 30469 27557 30481 27591
rect 30515 27588 30527 27591
rect 31662 27588 31668 27600
rect 30515 27560 31668 27588
rect 30515 27557 30527 27560
rect 30469 27551 30527 27557
rect 31662 27548 31668 27560
rect 31720 27548 31726 27600
rect 33520 27597 33548 27628
rect 33505 27591 33563 27597
rect 33505 27557 33517 27591
rect 33551 27557 33563 27591
rect 33505 27551 33563 27557
rect 33686 27548 33692 27600
rect 33744 27588 33750 27600
rect 35434 27588 35440 27600
rect 33744 27560 35440 27588
rect 33744 27548 33750 27560
rect 35434 27548 35440 27560
rect 35492 27548 35498 27600
rect 30300 27520 30328 27548
rect 30300 27492 30512 27520
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29748 27424 29837 27452
rect 27801 27415 27859 27421
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 26786 27344 26792 27396
rect 26844 27384 26850 27396
rect 27816 27384 27844 27415
rect 29914 27412 29920 27464
rect 29972 27452 29978 27464
rect 29972 27424 30017 27452
rect 29972 27412 29978 27424
rect 30098 27412 30104 27464
rect 30156 27412 30162 27464
rect 30331 27455 30389 27461
rect 30331 27421 30343 27455
rect 30377 27452 30389 27455
rect 30484 27452 30512 27492
rect 30650 27480 30656 27532
rect 30708 27520 30714 27532
rect 31113 27523 31171 27529
rect 31113 27520 31125 27523
rect 30708 27492 31125 27520
rect 30708 27480 30714 27492
rect 31113 27489 31125 27492
rect 31159 27489 31171 27523
rect 31113 27483 31171 27489
rect 32677 27523 32735 27529
rect 32677 27489 32689 27523
rect 32723 27520 32735 27523
rect 33410 27520 33416 27532
rect 32723 27492 33416 27520
rect 32723 27489 32735 27492
rect 32677 27483 32735 27489
rect 33410 27480 33416 27492
rect 33468 27480 33474 27532
rect 33594 27480 33600 27532
rect 33652 27520 33658 27532
rect 37185 27523 37243 27529
rect 33652 27492 37044 27520
rect 33652 27480 33658 27492
rect 31021 27455 31079 27461
rect 31021 27452 31033 27455
rect 30377 27424 31033 27452
rect 30377 27421 30389 27424
rect 30331 27415 30389 27421
rect 31021 27421 31033 27424
rect 31067 27421 31079 27455
rect 31021 27415 31079 27421
rect 31297 27455 31355 27461
rect 31297 27421 31309 27455
rect 31343 27421 31355 27455
rect 31297 27415 31355 27421
rect 26844 27356 27844 27384
rect 30193 27387 30251 27393
rect 26844 27344 26850 27356
rect 30193 27353 30205 27387
rect 30239 27353 30251 27387
rect 30193 27347 30251 27353
rect 27246 27316 27252 27328
rect 26292 27288 27252 27316
rect 26292 27276 26298 27288
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 27798 27276 27804 27328
rect 27856 27316 27862 27328
rect 28077 27319 28135 27325
rect 28077 27316 28089 27319
rect 27856 27288 28089 27316
rect 27856 27276 27862 27288
rect 28077 27285 28089 27288
rect 28123 27285 28135 27319
rect 30208 27316 30236 27347
rect 30926 27344 30932 27396
rect 30984 27384 30990 27396
rect 31312 27384 31340 27415
rect 32950 27412 32956 27464
rect 33008 27412 33014 27464
rect 33686 27412 33692 27464
rect 33744 27412 33750 27464
rect 33962 27412 33968 27464
rect 34020 27452 34026 27464
rect 34057 27455 34115 27461
rect 34057 27452 34069 27455
rect 34020 27424 34069 27452
rect 34020 27412 34026 27424
rect 34057 27421 34069 27424
rect 34103 27421 34115 27455
rect 34057 27415 34115 27421
rect 34514 27412 34520 27464
rect 34572 27452 34578 27464
rect 34885 27455 34943 27461
rect 34885 27452 34897 27455
rect 34572 27424 34897 27452
rect 34572 27412 34578 27424
rect 34885 27421 34897 27424
rect 34931 27421 34943 27455
rect 34885 27415 34943 27421
rect 34974 27412 34980 27464
rect 35032 27412 35038 27464
rect 35161 27455 35219 27461
rect 35161 27421 35173 27455
rect 35207 27452 35219 27455
rect 35526 27452 35532 27464
rect 35207 27424 35532 27452
rect 35207 27421 35219 27424
rect 35161 27415 35219 27421
rect 35526 27412 35532 27424
rect 35584 27412 35590 27464
rect 36909 27455 36967 27461
rect 36909 27421 36921 27455
rect 36955 27421 36967 27455
rect 37016 27452 37044 27492
rect 37185 27489 37197 27523
rect 37231 27520 37243 27523
rect 38930 27520 38936 27532
rect 37231 27492 38936 27520
rect 37231 27489 37243 27492
rect 37185 27483 37243 27489
rect 38930 27480 38936 27492
rect 38988 27480 38994 27532
rect 37829 27455 37887 27461
rect 37829 27452 37841 27455
rect 37016 27424 37841 27452
rect 36909 27415 36967 27421
rect 37829 27421 37841 27424
rect 37875 27421 37887 27455
rect 37829 27415 37887 27421
rect 30984 27356 31340 27384
rect 33781 27387 33839 27393
rect 30984 27344 30990 27356
rect 33781 27353 33793 27387
rect 33827 27353 33839 27387
rect 33781 27347 33839 27353
rect 30282 27316 30288 27328
rect 30208 27288 30288 27316
rect 28077 27279 28135 27285
rect 30282 27276 30288 27288
rect 30340 27276 30346 27328
rect 32030 27276 32036 27328
rect 32088 27316 32094 27328
rect 33796 27316 33824 27347
rect 33870 27344 33876 27396
rect 33928 27344 33934 27396
rect 35345 27387 35403 27393
rect 35345 27353 35357 27387
rect 35391 27384 35403 27387
rect 36924 27384 36952 27415
rect 37918 27384 37924 27396
rect 35391 27356 37924 27384
rect 35391 27353 35403 27356
rect 35345 27347 35403 27353
rect 37918 27344 37924 27356
rect 37976 27344 37982 27396
rect 38105 27387 38163 27393
rect 38105 27353 38117 27387
rect 38151 27384 38163 27387
rect 39022 27384 39028 27396
rect 38151 27356 39028 27384
rect 38151 27353 38163 27356
rect 38105 27347 38163 27353
rect 39022 27344 39028 27356
rect 39080 27344 39086 27396
rect 32088 27288 33824 27316
rect 32088 27276 32094 27288
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 4157 27115 4215 27121
rect 4157 27081 4169 27115
rect 4203 27112 4215 27115
rect 4430 27112 4436 27124
rect 4203 27084 4436 27112
rect 4203 27081 4215 27084
rect 4157 27075 4215 27081
rect 4430 27072 4436 27084
rect 4488 27112 4494 27124
rect 6733 27115 6791 27121
rect 4488 27084 6684 27112
rect 4488 27072 4494 27084
rect 3044 27047 3102 27053
rect 3044 27013 3056 27047
rect 3090 27044 3102 27047
rect 3970 27044 3976 27056
rect 3090 27016 3976 27044
rect 3090 27013 3102 27016
rect 3044 27007 3102 27013
rect 3970 27004 3976 27016
rect 4028 27004 4034 27056
rect 5534 27004 5540 27056
rect 5592 27004 5598 27056
rect 6656 27044 6684 27084
rect 6733 27081 6745 27115
rect 6779 27112 6791 27115
rect 7285 27115 7343 27121
rect 7285 27112 7297 27115
rect 6779 27084 7297 27112
rect 6779 27081 6791 27084
rect 6733 27075 6791 27081
rect 7285 27081 7297 27084
rect 7331 27081 7343 27115
rect 7285 27075 7343 27081
rect 7374 27072 7380 27124
rect 7432 27112 7438 27124
rect 8202 27112 8208 27124
rect 7432 27084 8208 27112
rect 7432 27072 7438 27084
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 12802 27072 12808 27124
rect 12860 27072 12866 27124
rect 13096 27084 15056 27112
rect 13096 27044 13124 27084
rect 6656 27016 13124 27044
rect 13170 27004 13176 27056
rect 13228 27004 13234 27056
rect 13998 27044 14004 27056
rect 13280 27016 14004 27044
rect 2774 26936 2780 26988
rect 2832 26936 2838 26988
rect 4798 26936 4804 26988
rect 4856 26976 4862 26988
rect 5077 26979 5135 26985
rect 5077 26976 5089 26979
rect 4856 26948 5089 26976
rect 4856 26936 4862 26948
rect 5077 26945 5089 26948
rect 5123 26945 5135 26979
rect 5077 26939 5135 26945
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26976 5319 26979
rect 5350 26976 5356 26988
rect 5307 26948 5356 26976
rect 5307 26945 5319 26948
rect 5261 26939 5319 26945
rect 5350 26936 5356 26948
rect 5408 26976 5414 26988
rect 5902 26976 5908 26988
rect 5408 26948 5908 26976
rect 5408 26936 5414 26948
rect 5902 26936 5908 26948
rect 5960 26936 5966 26988
rect 6086 26936 6092 26988
rect 6144 26976 6150 26988
rect 6549 26979 6607 26985
rect 6549 26976 6561 26979
rect 6144 26948 6561 26976
rect 6144 26936 6150 26948
rect 6549 26945 6561 26948
rect 6595 26976 6607 26979
rect 6638 26976 6644 26988
rect 6595 26948 6644 26976
rect 6595 26945 6607 26948
rect 6549 26939 6607 26945
rect 6638 26936 6644 26948
rect 6696 26936 6702 26988
rect 6825 26979 6883 26985
rect 6825 26945 6837 26979
rect 6871 26945 6883 26979
rect 6825 26939 6883 26945
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 6840 26908 6868 26939
rect 7282 26936 7288 26988
rect 7340 26936 7346 26988
rect 7466 26936 7472 26988
rect 7524 26936 7530 26988
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26976 8079 26979
rect 8110 26976 8116 26988
rect 8067 26948 8116 26976
rect 8067 26945 8079 26948
rect 8021 26939 8079 26945
rect 6236 26880 6868 26908
rect 6236 26868 6242 26880
rect 6914 26868 6920 26920
rect 6972 26908 6978 26920
rect 8036 26908 8064 26939
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 8202 26936 8208 26988
rect 8260 26976 8266 26988
rect 8297 26979 8355 26985
rect 8297 26976 8309 26979
rect 8260 26948 8309 26976
rect 8260 26936 8266 26948
rect 8297 26945 8309 26948
rect 8343 26945 8355 26979
rect 8895 26979 8953 26985
rect 8895 26976 8907 26979
rect 8297 26939 8355 26945
rect 8680 26948 8907 26976
rect 6972 26880 8064 26908
rect 6972 26868 6978 26880
rect 8018 26800 8024 26852
rect 8076 26840 8082 26852
rect 8680 26840 8708 26948
rect 8895 26945 8907 26948
rect 8941 26945 8953 26979
rect 8895 26939 8953 26945
rect 9030 26936 9036 26988
rect 9088 26936 9094 26988
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26945 9183 26979
rect 9125 26939 9183 26945
rect 8754 26868 8760 26920
rect 8812 26868 8818 26920
rect 9140 26908 9168 26939
rect 9214 26936 9220 26988
rect 9272 26936 9278 26988
rect 10226 26936 10232 26988
rect 10284 26936 10290 26988
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26976 10471 26979
rect 10502 26976 10508 26988
rect 10459 26948 10508 26976
rect 10459 26945 10471 26948
rect 10413 26939 10471 26945
rect 10502 26936 10508 26948
rect 10560 26936 10566 26988
rect 12986 26936 12992 26988
rect 13044 26936 13050 26988
rect 13081 26979 13139 26985
rect 13081 26945 13093 26979
rect 13127 26976 13139 26979
rect 13280 26976 13308 27016
rect 13998 27004 14004 27016
rect 14056 27004 14062 27056
rect 15028 27044 15056 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 15933 27115 15991 27121
rect 15933 27112 15945 27115
rect 15160 27084 15945 27112
rect 15160 27072 15166 27084
rect 15933 27081 15945 27084
rect 15979 27112 15991 27115
rect 17126 27112 17132 27124
rect 15979 27084 17132 27112
rect 15979 27081 15991 27084
rect 15933 27075 15991 27081
rect 17126 27072 17132 27084
rect 17184 27072 17190 27124
rect 20165 27115 20223 27121
rect 20165 27081 20177 27115
rect 20211 27112 20223 27115
rect 20254 27112 20260 27124
rect 20211 27084 20260 27112
rect 20211 27081 20223 27084
rect 20165 27075 20223 27081
rect 20254 27072 20260 27084
rect 20312 27072 20318 27124
rect 22465 27115 22523 27121
rect 20364 27084 22416 27112
rect 16942 27044 16948 27056
rect 15028 27016 16948 27044
rect 16942 27004 16948 27016
rect 17000 27004 17006 27056
rect 17144 27016 19012 27044
rect 13127 26948 13308 26976
rect 13127 26945 13139 26948
rect 13081 26939 13139 26945
rect 13354 26936 13360 26988
rect 13412 26936 13418 26988
rect 14826 26985 14832 26988
rect 14820 26939 14832 26985
rect 14826 26936 14832 26939
rect 14884 26936 14890 26988
rect 9048 26880 9168 26908
rect 8076 26812 8708 26840
rect 8076 26800 8082 26812
rect 4706 26732 4712 26784
rect 4764 26772 4770 26784
rect 4893 26775 4951 26781
rect 4893 26772 4905 26775
rect 4764 26744 4905 26772
rect 4764 26732 4770 26744
rect 4893 26741 4905 26744
rect 4939 26741 4951 26775
rect 4893 26735 4951 26741
rect 5445 26775 5503 26781
rect 5445 26741 5457 26775
rect 5491 26772 5503 26775
rect 6549 26775 6607 26781
rect 6549 26772 6561 26775
rect 5491 26744 6561 26772
rect 5491 26741 5503 26744
rect 5445 26735 5503 26741
rect 6549 26741 6561 26744
rect 6595 26741 6607 26775
rect 6549 26735 6607 26741
rect 8202 26732 8208 26784
rect 8260 26772 8266 26784
rect 9048 26772 9076 26880
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 13372 26908 13400 26936
rect 12492 26880 13400 26908
rect 12492 26868 12498 26880
rect 14458 26868 14464 26920
rect 14516 26908 14522 26920
rect 14553 26911 14611 26917
rect 14553 26908 14565 26911
rect 14516 26880 14565 26908
rect 14516 26868 14522 26880
rect 14553 26877 14565 26880
rect 14599 26877 14611 26911
rect 14553 26871 14611 26877
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 17144 26917 17172 27016
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26976 18107 26979
rect 18230 26976 18236 26988
rect 18095 26948 18236 26976
rect 18095 26945 18107 26948
rect 18049 26939 18107 26945
rect 18230 26936 18236 26948
rect 18288 26936 18294 26988
rect 18984 26985 19012 27016
rect 19058 27004 19064 27056
rect 19116 27044 19122 27056
rect 19116 27016 20116 27044
rect 19116 27004 19122 27016
rect 18969 26979 19027 26985
rect 18969 26945 18981 26979
rect 19015 26945 19027 26979
rect 18969 26939 19027 26945
rect 19245 26979 19303 26985
rect 19245 26945 19257 26979
rect 19291 26976 19303 26979
rect 19794 26976 19800 26988
rect 19291 26948 19800 26976
rect 19291 26945 19303 26948
rect 19245 26939 19303 26945
rect 19794 26936 19800 26948
rect 19852 26936 19858 26988
rect 20088 26985 20116 27016
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26945 20131 26979
rect 20073 26939 20131 26945
rect 17129 26911 17187 26917
rect 17129 26908 17141 26911
rect 16816 26880 17141 26908
rect 16816 26868 16822 26880
rect 17129 26877 17141 26880
rect 17175 26877 17187 26911
rect 17129 26871 17187 26877
rect 18138 26868 18144 26920
rect 18196 26868 18202 26920
rect 20088 26908 20116 26939
rect 20254 26936 20260 26988
rect 20312 26976 20318 26988
rect 20364 26976 20392 27084
rect 20530 27004 20536 27056
rect 20588 27044 20594 27056
rect 22005 27047 22063 27053
rect 22005 27044 22017 27047
rect 20588 27016 22017 27044
rect 20588 27004 20594 27016
rect 22005 27013 22017 27016
rect 22051 27013 22063 27047
rect 22388 27044 22416 27084
rect 22465 27081 22477 27115
rect 22511 27112 22523 27115
rect 22511 27084 23888 27112
rect 22511 27081 22523 27084
rect 22465 27075 22523 27081
rect 22388 27016 23520 27044
rect 22005 27007 22063 27013
rect 20312 26948 20392 26976
rect 20809 26979 20867 26985
rect 20312 26936 20318 26948
rect 20809 26945 20821 26979
rect 20855 26976 20867 26979
rect 20990 26976 20996 26988
rect 20855 26948 20996 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 22281 26979 22339 26985
rect 22281 26945 22293 26979
rect 22327 26976 22339 26979
rect 22646 26976 22652 26988
rect 22327 26948 22652 26976
rect 22327 26945 22339 26948
rect 22281 26939 22339 26945
rect 22646 26936 22652 26948
rect 22704 26936 22710 26988
rect 22922 26936 22928 26988
rect 22980 26936 22986 26988
rect 23198 26936 23204 26988
rect 23256 26936 23262 26988
rect 20088 26880 20852 26908
rect 9401 26843 9459 26849
rect 9401 26809 9413 26843
rect 9447 26840 9459 26843
rect 14366 26840 14372 26852
rect 9447 26812 14372 26840
rect 9447 26809 9459 26812
rect 9401 26803 9459 26809
rect 14366 26800 14372 26812
rect 14424 26800 14430 26852
rect 17034 26800 17040 26852
rect 17092 26800 17098 26852
rect 17218 26800 17224 26852
rect 17276 26840 17282 26852
rect 18322 26840 18328 26852
rect 17276 26812 18328 26840
rect 17276 26800 17282 26812
rect 18322 26800 18328 26812
rect 18380 26800 18386 26852
rect 18969 26843 19027 26849
rect 18969 26809 18981 26843
rect 19015 26809 19027 26843
rect 20824 26840 20852 26880
rect 20898 26868 20904 26920
rect 20956 26868 20962 26920
rect 21726 26908 21732 26920
rect 20999 26880 21732 26908
rect 20999 26840 21027 26880
rect 21726 26868 21732 26880
rect 21784 26868 21790 26920
rect 22097 26911 22155 26917
rect 22097 26877 22109 26911
rect 22143 26877 22155 26911
rect 23017 26911 23075 26917
rect 23017 26908 23029 26911
rect 22097 26871 22155 26877
rect 22204 26880 23029 26908
rect 20824 26812 21027 26840
rect 21177 26843 21235 26849
rect 18969 26803 19027 26809
rect 21177 26809 21189 26843
rect 21223 26840 21235 26843
rect 22112 26840 22140 26871
rect 21223 26812 22140 26840
rect 21223 26809 21235 26812
rect 21177 26803 21235 26809
rect 8260 26744 9076 26772
rect 8260 26732 8266 26744
rect 10226 26732 10232 26784
rect 10284 26732 10290 26784
rect 10410 26732 10416 26784
rect 10468 26772 10474 26784
rect 16390 26772 16396 26784
rect 10468 26744 16396 26772
rect 10468 26732 10474 26744
rect 16390 26732 16396 26744
rect 16448 26732 16454 26784
rect 16482 26732 16488 26784
rect 16540 26772 16546 26784
rect 18984 26772 19012 26803
rect 20714 26772 20720 26784
rect 16540 26744 20720 26772
rect 16540 26732 16546 26744
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 20993 26775 21051 26781
rect 20993 26741 21005 26775
rect 21039 26772 21051 26775
rect 21082 26772 21088 26784
rect 21039 26744 21088 26772
rect 21039 26741 21051 26744
rect 20993 26735 21051 26741
rect 21082 26732 21088 26744
rect 21140 26772 21146 26784
rect 21542 26772 21548 26784
rect 21140 26744 21548 26772
rect 21140 26732 21146 26744
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 22094 26732 22100 26784
rect 22152 26772 22158 26784
rect 22204 26772 22232 26880
rect 23017 26877 23029 26880
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 23385 26843 23443 26849
rect 23385 26840 23397 26843
rect 22296 26812 23397 26840
rect 22296 26781 22324 26812
rect 23385 26809 23397 26812
rect 23431 26809 23443 26843
rect 23385 26803 23443 26809
rect 22152 26744 22232 26772
rect 22281 26775 22339 26781
rect 22152 26732 22158 26744
rect 22281 26741 22293 26775
rect 22327 26741 22339 26775
rect 22281 26735 22339 26741
rect 23014 26732 23020 26784
rect 23072 26732 23078 26784
rect 23492 26772 23520 27016
rect 23860 26908 23888 27084
rect 24578 27072 24584 27124
rect 24636 27072 24642 27124
rect 24946 27072 24952 27124
rect 25004 27112 25010 27124
rect 26329 27115 26387 27121
rect 25004 27084 26280 27112
rect 25004 27072 25010 27084
rect 24029 27047 24087 27053
rect 24029 27013 24041 27047
rect 24075 27044 24087 27047
rect 25498 27044 25504 27056
rect 24075 27016 25504 27044
rect 24075 27013 24087 27016
rect 24029 27007 24087 27013
rect 23934 26936 23940 26988
rect 23992 26936 23998 26988
rect 24118 26936 24124 26988
rect 24176 26936 24182 26988
rect 24762 26936 24768 26988
rect 24820 26936 24826 26988
rect 24854 26936 24860 26988
rect 24912 26936 24918 26988
rect 25056 26985 25084 27016
rect 25498 27004 25504 27016
rect 25556 27004 25562 27056
rect 26142 27004 26148 27056
rect 26200 27004 26206 27056
rect 26252 27044 26280 27084
rect 26329 27081 26341 27115
rect 26375 27112 26387 27115
rect 27154 27112 27160 27124
rect 26375 27084 27160 27112
rect 26375 27081 26387 27084
rect 26329 27075 26387 27081
rect 27154 27072 27160 27084
rect 27212 27072 27218 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 31110 27112 31116 27124
rect 27672 27084 31116 27112
rect 27672 27072 27678 27084
rect 31110 27072 31116 27084
rect 31168 27072 31174 27124
rect 32950 27072 32956 27124
rect 33008 27112 33014 27124
rect 37550 27112 37556 27124
rect 33008 27084 37556 27112
rect 33008 27072 33014 27084
rect 37550 27072 37556 27084
rect 37608 27072 37614 27124
rect 37918 27072 37924 27124
rect 37976 27072 37982 27124
rect 30377 27047 30435 27053
rect 26252 27016 28120 27044
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 25130 26936 25136 26988
rect 25188 26976 25194 26988
rect 25225 26979 25283 26985
rect 25225 26976 25237 26979
rect 25188 26948 25237 26976
rect 25188 26936 25194 26948
rect 25225 26945 25237 26948
rect 25271 26945 25283 26979
rect 25225 26939 25283 26945
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 27396 26948 27568 26976
rect 27396 26936 27402 26948
rect 27430 26908 27436 26920
rect 23860 26880 27436 26908
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 27540 26908 27568 26948
rect 27614 26936 27620 26988
rect 27672 26936 27678 26988
rect 28092 26985 28120 27016
rect 30377 27013 30389 27047
rect 30423 27044 30435 27047
rect 31389 27047 31447 27053
rect 31389 27044 31401 27047
rect 30423 27016 31401 27044
rect 30423 27013 30435 27016
rect 30377 27007 30435 27013
rect 31389 27013 31401 27016
rect 31435 27044 31447 27047
rect 32214 27044 32220 27056
rect 31435 27016 32220 27044
rect 31435 27013 31447 27016
rect 31389 27007 31447 27013
rect 32214 27004 32220 27016
rect 32272 27004 32278 27056
rect 34790 27044 34796 27056
rect 32600 27016 34796 27044
rect 32600 26988 32628 27016
rect 34790 27004 34796 27016
rect 34848 27004 34854 27056
rect 35621 27047 35679 27053
rect 35621 27013 35633 27047
rect 35667 27044 35679 27047
rect 36354 27044 36360 27056
rect 35667 27016 36360 27044
rect 35667 27013 35679 27016
rect 35621 27007 35679 27013
rect 36354 27004 36360 27016
rect 36412 27004 36418 27056
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26976 28135 26979
rect 28994 26976 29000 26988
rect 28123 26948 29000 26976
rect 28123 26945 28135 26948
rect 28077 26939 28135 26945
rect 28994 26936 29000 26948
rect 29052 26976 29058 26988
rect 29089 26979 29147 26985
rect 29089 26976 29101 26979
rect 29052 26948 29101 26976
rect 29052 26936 29058 26948
rect 29089 26945 29101 26948
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 29730 26936 29736 26988
rect 29788 26936 29794 26988
rect 30098 26936 30104 26988
rect 30156 26976 30162 26988
rect 30837 26979 30895 26985
rect 30837 26976 30849 26979
rect 30156 26948 30849 26976
rect 30156 26936 30162 26948
rect 30837 26945 30849 26948
rect 30883 26945 30895 26979
rect 30837 26939 30895 26945
rect 31205 26979 31263 26985
rect 31205 26945 31217 26979
rect 31251 26976 31263 26979
rect 31478 26976 31484 26988
rect 31251 26948 31484 26976
rect 31251 26945 31263 26948
rect 31205 26939 31263 26945
rect 31478 26936 31484 26948
rect 31536 26936 31542 26988
rect 32582 26936 32588 26988
rect 32640 26936 32646 26988
rect 33042 26936 33048 26988
rect 33100 26976 33106 26988
rect 34146 26976 34152 26988
rect 33100 26948 34152 26976
rect 33100 26936 33106 26948
rect 34146 26936 34152 26948
rect 34204 26936 34210 26988
rect 34333 26979 34391 26985
rect 34333 26945 34345 26979
rect 34379 26976 34391 26979
rect 34698 26976 34704 26988
rect 34379 26948 34704 26976
rect 34379 26945 34391 26948
rect 34333 26939 34391 26945
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 37826 26936 37832 26988
rect 37884 26936 37890 26988
rect 28353 26911 28411 26917
rect 28353 26908 28365 26911
rect 27540 26880 28365 26908
rect 28353 26877 28365 26880
rect 28399 26908 28411 26911
rect 31386 26908 31392 26920
rect 28399 26880 31392 26908
rect 28399 26877 28411 26880
rect 28353 26871 28411 26877
rect 31386 26868 31392 26880
rect 31444 26868 31450 26920
rect 32674 26868 32680 26920
rect 32732 26908 32738 26920
rect 33318 26908 33324 26920
rect 32732 26880 33324 26908
rect 32732 26868 32738 26880
rect 33318 26868 33324 26880
rect 33376 26868 33382 26920
rect 33410 26868 33416 26920
rect 33468 26908 33474 26920
rect 38013 26911 38071 26917
rect 38013 26908 38025 26911
rect 33468 26880 38025 26908
rect 33468 26868 33474 26880
rect 38013 26877 38025 26880
rect 38059 26908 38071 26911
rect 38102 26908 38108 26920
rect 38059 26880 38108 26908
rect 38059 26877 38071 26880
rect 38013 26871 38071 26877
rect 38102 26868 38108 26880
rect 38160 26868 38166 26920
rect 23566 26800 23572 26852
rect 23624 26840 23630 26852
rect 24854 26840 24860 26852
rect 23624 26812 24860 26840
rect 23624 26800 23630 26812
rect 24854 26800 24860 26812
rect 24912 26800 24918 26852
rect 24946 26800 24952 26852
rect 25004 26800 25010 26852
rect 26513 26843 26571 26849
rect 26513 26809 26525 26843
rect 26559 26840 26571 26843
rect 32950 26840 32956 26852
rect 26559 26812 32956 26840
rect 26559 26809 26571 26812
rect 26513 26803 26571 26809
rect 32950 26800 32956 26812
rect 33008 26800 33014 26852
rect 34974 26800 34980 26852
rect 35032 26840 35038 26852
rect 35802 26840 35808 26852
rect 35032 26812 35808 26840
rect 35032 26800 35038 26812
rect 35802 26800 35808 26812
rect 35860 26800 35866 26852
rect 25038 26772 25044 26784
rect 23492 26744 25044 26772
rect 25038 26732 25044 26744
rect 25096 26732 25102 26784
rect 26326 26732 26332 26784
rect 26384 26732 26390 26784
rect 34333 26775 34391 26781
rect 34333 26741 34345 26775
rect 34379 26772 34391 26775
rect 36262 26772 36268 26784
rect 34379 26744 36268 26772
rect 34379 26741 34391 26744
rect 34333 26735 34391 26741
rect 36262 26732 36268 26744
rect 36320 26732 36326 26784
rect 36814 26732 36820 26784
rect 36872 26772 36878 26784
rect 37461 26775 37519 26781
rect 37461 26772 37473 26775
rect 36872 26744 37473 26772
rect 36872 26732 36878 26744
rect 37461 26741 37473 26744
rect 37507 26741 37519 26775
rect 37461 26735 37519 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 8110 26528 8116 26580
rect 8168 26568 8174 26580
rect 9309 26571 9367 26577
rect 9309 26568 9321 26571
rect 8168 26540 9321 26568
rect 8168 26528 8174 26540
rect 9309 26537 9321 26540
rect 9355 26568 9367 26571
rect 10318 26568 10324 26580
rect 9355 26540 10324 26568
rect 9355 26537 9367 26540
rect 9309 26531 9367 26537
rect 10318 26528 10324 26540
rect 10376 26568 10382 26580
rect 12250 26568 12256 26580
rect 10376 26540 12256 26568
rect 10376 26528 10382 26540
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 14737 26571 14795 26577
rect 14737 26537 14749 26571
rect 14783 26568 14795 26571
rect 14826 26568 14832 26580
rect 14783 26540 14832 26568
rect 14783 26537 14795 26540
rect 14737 26531 14795 26537
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 16390 26528 16396 26580
rect 16448 26568 16454 26580
rect 19426 26568 19432 26580
rect 16448 26540 19432 26568
rect 16448 26528 16454 26540
rect 19426 26528 19432 26540
rect 19484 26528 19490 26580
rect 22833 26571 22891 26577
rect 22833 26537 22845 26571
rect 22879 26568 22891 26571
rect 23014 26568 23020 26580
rect 22879 26540 23020 26568
rect 22879 26537 22891 26540
rect 22833 26531 22891 26537
rect 23014 26528 23020 26540
rect 23072 26568 23078 26580
rect 23477 26571 23535 26577
rect 23477 26568 23489 26571
rect 23072 26540 23489 26568
rect 23072 26528 23078 26540
rect 23477 26537 23489 26540
rect 23523 26537 23535 26571
rect 23477 26531 23535 26537
rect 23658 26528 23664 26580
rect 23716 26568 23722 26580
rect 25866 26568 25872 26580
rect 23716 26540 25872 26568
rect 23716 26528 23722 26540
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 26510 26528 26516 26580
rect 26568 26568 26574 26580
rect 26568 26540 28994 26568
rect 26568 26528 26574 26540
rect 6362 26460 6368 26512
rect 6420 26500 6426 26512
rect 10410 26500 10416 26512
rect 6420 26472 10416 26500
rect 6420 26460 6426 26472
rect 10410 26460 10416 26472
rect 10468 26460 10474 26512
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 20438 26500 20444 26512
rect 14148 26472 15332 26500
rect 14148 26460 14154 26472
rect 5077 26435 5135 26441
rect 5077 26401 5089 26435
rect 5123 26432 5135 26435
rect 5442 26432 5448 26444
rect 5123 26404 5448 26432
rect 5123 26401 5135 26404
rect 5077 26395 5135 26401
rect 5442 26392 5448 26404
rect 5500 26432 5506 26444
rect 5997 26435 6055 26441
rect 5997 26432 6009 26435
rect 5500 26404 6009 26432
rect 5500 26392 5506 26404
rect 5997 26401 6009 26404
rect 6043 26401 6055 26435
rect 5997 26395 6055 26401
rect 8386 26392 8392 26444
rect 8444 26432 8450 26444
rect 11057 26435 11115 26441
rect 11057 26432 11069 26435
rect 8444 26404 11069 26432
rect 8444 26392 8450 26404
rect 11057 26401 11069 26404
rect 11103 26401 11115 26435
rect 11057 26395 11115 26401
rect 14366 26392 14372 26444
rect 14424 26432 14430 26444
rect 15304 26441 15332 26472
rect 20272 26472 20444 26500
rect 15197 26435 15255 26441
rect 15197 26432 15209 26435
rect 14424 26404 15209 26432
rect 14424 26392 14430 26404
rect 15197 26401 15209 26404
rect 15243 26401 15255 26435
rect 15197 26395 15255 26401
rect 15289 26435 15347 26441
rect 15289 26401 15301 26435
rect 15335 26401 15347 26435
rect 15289 26395 15347 26401
rect 16025 26435 16083 26441
rect 16025 26401 16037 26435
rect 16071 26432 16083 26435
rect 17218 26432 17224 26444
rect 16071 26404 17224 26432
rect 16071 26401 16083 26404
rect 16025 26395 16083 26401
rect 17218 26392 17224 26404
rect 17276 26392 17282 26444
rect 17954 26432 17960 26444
rect 17604 26404 17960 26432
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 5169 26367 5227 26373
rect 5169 26364 5181 26367
rect 4948 26336 5181 26364
rect 4948 26324 4954 26336
rect 5169 26333 5181 26336
rect 5215 26333 5227 26367
rect 5169 26327 5227 26333
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26364 5411 26367
rect 5626 26364 5632 26376
rect 5399 26336 5632 26364
rect 5399 26333 5411 26336
rect 5353 26327 5411 26333
rect 5276 26296 5304 26327
rect 5626 26324 5632 26336
rect 5684 26324 5690 26376
rect 5902 26324 5908 26376
rect 5960 26324 5966 26376
rect 6086 26324 6092 26376
rect 6144 26324 6150 26376
rect 8294 26324 8300 26376
rect 8352 26324 8358 26376
rect 8573 26367 8631 26373
rect 8573 26333 8585 26367
rect 8619 26364 8631 26367
rect 8754 26364 8760 26376
rect 8619 26336 8760 26364
rect 8619 26333 8631 26336
rect 8573 26327 8631 26333
rect 8754 26324 8760 26336
rect 8812 26364 8818 26376
rect 10597 26367 10655 26373
rect 8812 26336 9168 26364
rect 8812 26324 8818 26336
rect 5718 26296 5724 26308
rect 5276 26268 5724 26296
rect 5718 26256 5724 26268
rect 5776 26256 5782 26308
rect 6178 26256 6184 26308
rect 6236 26296 6242 26308
rect 8205 26299 8263 26305
rect 8205 26296 8217 26299
rect 6236 26268 8217 26296
rect 6236 26256 6242 26268
rect 8205 26265 8217 26268
rect 8251 26265 8263 26299
rect 8205 26259 8263 26265
rect 4614 26188 4620 26240
rect 4672 26228 4678 26240
rect 9140 26237 9168 26336
rect 10597 26333 10609 26367
rect 10643 26364 10655 26367
rect 10643 26336 12434 26364
rect 10643 26333 10655 26336
rect 10597 26327 10655 26333
rect 9490 26256 9496 26308
rect 9548 26256 9554 26308
rect 11146 26256 11152 26308
rect 11204 26296 11210 26308
rect 11302 26299 11360 26305
rect 11302 26296 11314 26299
rect 11204 26268 11314 26296
rect 11204 26256 11210 26268
rect 11302 26265 11314 26268
rect 11348 26265 11360 26299
rect 12406 26296 12434 26336
rect 15102 26324 15108 26376
rect 15160 26324 15166 26376
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26364 16267 26367
rect 17034 26364 17040 26376
rect 16255 26336 17040 26364
rect 16255 26333 16267 26336
rect 16209 26327 16267 26333
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 17604 26373 17632 26404
rect 17954 26392 17960 26404
rect 18012 26392 18018 26444
rect 20272 26432 20300 26472
rect 20438 26460 20444 26472
rect 20496 26500 20502 26512
rect 21266 26500 21272 26512
rect 20496 26472 21272 26500
rect 20496 26460 20502 26472
rect 21266 26460 21272 26472
rect 21324 26460 21330 26512
rect 21450 26460 21456 26512
rect 21508 26500 21514 26512
rect 21545 26503 21603 26509
rect 21545 26500 21557 26503
rect 21508 26472 21557 26500
rect 21508 26460 21514 26472
rect 21545 26469 21557 26472
rect 21591 26469 21603 26503
rect 21545 26463 21603 26469
rect 21726 26460 21732 26512
rect 21784 26500 21790 26512
rect 21784 26472 23980 26500
rect 21784 26460 21790 26472
rect 18248 26404 20300 26432
rect 17589 26367 17647 26373
rect 17589 26364 17601 26367
rect 17144 26336 17601 26364
rect 13630 26296 13636 26308
rect 12406 26268 13636 26296
rect 11302 26259 11360 26265
rect 13630 26256 13636 26268
rect 13688 26256 13694 26308
rect 16393 26299 16451 26305
rect 16393 26265 16405 26299
rect 16439 26296 16451 26299
rect 17144 26296 17172 26336
rect 17589 26333 17601 26336
rect 17635 26333 17647 26367
rect 17589 26327 17647 26333
rect 17678 26324 17684 26376
rect 17736 26324 17742 26376
rect 18248 26373 18276 26404
rect 20346 26392 20352 26444
rect 20404 26432 20410 26444
rect 20625 26435 20683 26441
rect 20625 26432 20637 26435
rect 20404 26404 20637 26432
rect 20404 26392 20410 26404
rect 20625 26401 20637 26404
rect 20671 26401 20683 26435
rect 21634 26432 21640 26444
rect 20625 26395 20683 26401
rect 20916 26404 21640 26432
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 18380 26336 19564 26364
rect 18380 26324 18386 26336
rect 16439 26268 17172 26296
rect 16439 26265 16451 26268
rect 16393 26259 16451 26265
rect 17218 26256 17224 26308
rect 17276 26296 17282 26308
rect 19429 26299 19487 26305
rect 19429 26296 19441 26299
rect 17276 26268 19441 26296
rect 17276 26256 17282 26268
rect 19429 26265 19441 26268
rect 19475 26265 19487 26299
rect 19536 26296 19564 26336
rect 19610 26324 19616 26376
rect 19668 26324 19674 26376
rect 19702 26324 19708 26376
rect 19760 26324 19766 26376
rect 19794 26324 19800 26376
rect 19852 26364 19858 26376
rect 20530 26364 20536 26376
rect 19852 26336 20536 26364
rect 19852 26324 19858 26336
rect 20530 26324 20536 26336
rect 20588 26364 20594 26376
rect 20916 26373 20944 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 22649 26435 22707 26441
rect 22649 26432 22661 26435
rect 21836 26404 22661 26432
rect 20901 26367 20959 26373
rect 20901 26364 20913 26367
rect 20588 26336 20913 26364
rect 20588 26324 20594 26336
rect 20901 26333 20913 26336
rect 20947 26333 20959 26367
rect 20901 26327 20959 26333
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26364 21143 26367
rect 21174 26364 21180 26376
rect 21131 26336 21180 26364
rect 21131 26333 21143 26336
rect 21085 26327 21143 26333
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 21450 26324 21456 26376
rect 21508 26364 21514 26376
rect 21748 26367 21806 26373
rect 21748 26364 21760 26367
rect 21508 26336 21760 26364
rect 21508 26324 21514 26336
rect 21748 26333 21760 26336
rect 21794 26333 21806 26367
rect 21748 26327 21806 26333
rect 21836 26296 21864 26404
rect 22649 26401 22661 26404
rect 22695 26432 22707 26435
rect 23842 26432 23848 26444
rect 22695 26404 23848 26432
rect 22695 26401 22707 26404
rect 22649 26395 22707 26401
rect 23842 26392 23848 26404
rect 23900 26392 23906 26444
rect 23952 26432 23980 26472
rect 24026 26460 24032 26512
rect 24084 26500 24090 26512
rect 26326 26500 26332 26512
rect 24084 26472 26332 26500
rect 24084 26460 24090 26472
rect 23952 26404 24808 26432
rect 22002 26324 22008 26376
rect 22060 26324 22066 26376
rect 22830 26324 22836 26376
rect 22888 26364 22894 26376
rect 23382 26364 23388 26376
rect 22888 26336 23388 26364
rect 22888 26324 22894 26336
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 23566 26364 23572 26376
rect 23523 26336 23572 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 23658 26324 23664 26376
rect 23716 26324 23722 26376
rect 24780 26373 24808 26404
rect 24765 26367 24823 26373
rect 24765 26333 24777 26367
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 19536 26268 21864 26296
rect 22557 26299 22615 26305
rect 19429 26259 19487 26265
rect 22557 26265 22569 26299
rect 22603 26265 22615 26299
rect 22557 26259 22615 26265
rect 24581 26299 24639 26305
rect 24581 26265 24593 26299
rect 24627 26296 24639 26299
rect 24670 26296 24676 26308
rect 24627 26268 24676 26296
rect 24627 26265 24639 26268
rect 24581 26259 24639 26265
rect 9306 26237 9312 26240
rect 4893 26231 4951 26237
rect 4893 26228 4905 26231
rect 4672 26200 4905 26228
rect 4672 26188 4678 26200
rect 4893 26197 4905 26200
rect 4939 26197 4951 26231
rect 4893 26191 4951 26197
rect 9125 26231 9183 26237
rect 9125 26197 9137 26231
rect 9171 26197 9183 26231
rect 9125 26191 9183 26197
rect 9293 26231 9312 26237
rect 9293 26197 9305 26231
rect 9293 26191 9312 26197
rect 9306 26188 9312 26191
rect 9364 26188 9370 26240
rect 9766 26188 9772 26240
rect 9824 26228 9830 26240
rect 10413 26231 10471 26237
rect 10413 26228 10425 26231
rect 9824 26200 10425 26228
rect 9824 26188 9830 26200
rect 10413 26197 10425 26200
rect 10459 26228 10471 26231
rect 10962 26228 10968 26240
rect 10459 26200 10968 26228
rect 10459 26197 10471 26200
rect 10413 26191 10471 26197
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 12437 26231 12495 26237
rect 12437 26197 12449 26231
rect 12483 26228 12495 26231
rect 12526 26228 12532 26240
rect 12483 26200 12532 26228
rect 12483 26197 12495 26200
rect 12437 26191 12495 26197
rect 12526 26188 12532 26200
rect 12584 26188 12590 26240
rect 18046 26188 18052 26240
rect 18104 26188 18110 26240
rect 18138 26188 18144 26240
rect 18196 26228 18202 26240
rect 19702 26228 19708 26240
rect 18196 26200 19708 26228
rect 18196 26188 18202 26200
rect 19702 26188 19708 26200
rect 19760 26228 19766 26240
rect 20070 26228 20076 26240
rect 19760 26200 20076 26228
rect 19760 26188 19766 26200
rect 20070 26188 20076 26200
rect 20128 26188 20134 26240
rect 21913 26231 21971 26237
rect 21913 26197 21925 26231
rect 21959 26228 21971 26231
rect 22002 26228 22008 26240
rect 21959 26200 22008 26228
rect 21959 26197 21971 26200
rect 21913 26191 21971 26197
rect 22002 26188 22008 26200
rect 22060 26188 22066 26240
rect 22370 26188 22376 26240
rect 22428 26228 22434 26240
rect 22572 26228 22600 26259
rect 24670 26256 24676 26268
rect 24728 26256 24734 26308
rect 24780 26296 24808 26327
rect 24946 26324 24952 26376
rect 25004 26324 25010 26376
rect 25038 26324 25044 26376
rect 25096 26324 25102 26376
rect 25130 26324 25136 26376
rect 25188 26324 25194 26376
rect 25317 26367 25375 26373
rect 25317 26333 25329 26367
rect 25363 26364 25375 26367
rect 25516 26364 25544 26472
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 27706 26460 27712 26512
rect 27764 26500 27770 26512
rect 27982 26500 27988 26512
rect 27764 26472 27988 26500
rect 27764 26460 27770 26472
rect 27982 26460 27988 26472
rect 28040 26500 28046 26512
rect 28040 26472 28120 26500
rect 28040 26460 28046 26472
rect 25363 26336 25544 26364
rect 27709 26367 27767 26373
rect 25363 26333 25375 26336
rect 25317 26327 25375 26333
rect 27709 26333 27721 26367
rect 27755 26333 27767 26367
rect 27709 26327 27767 26333
rect 26786 26296 26792 26308
rect 24780 26268 26792 26296
rect 26786 26256 26792 26268
rect 26844 26256 26850 26308
rect 27724 26296 27752 26327
rect 27890 26324 27896 26376
rect 27948 26324 27954 26376
rect 27982 26324 27988 26376
rect 28040 26324 28046 26376
rect 28092 26373 28120 26472
rect 28258 26460 28264 26512
rect 28316 26460 28322 26512
rect 28966 26500 28994 26540
rect 29546 26528 29552 26580
rect 29604 26568 29610 26580
rect 33870 26568 33876 26580
rect 29604 26540 33876 26568
rect 29604 26528 29610 26540
rect 33870 26528 33876 26540
rect 33928 26568 33934 26580
rect 33928 26540 35389 26568
rect 33928 26528 33934 26540
rect 29914 26500 29920 26512
rect 28966 26472 29920 26500
rect 29914 26460 29920 26472
rect 29972 26500 29978 26512
rect 30929 26503 30987 26509
rect 30929 26500 30941 26503
rect 29972 26472 30941 26500
rect 29972 26460 29978 26472
rect 30929 26469 30941 26472
rect 30975 26500 30987 26503
rect 32674 26500 32680 26512
rect 30975 26472 31340 26500
rect 30975 26469 30987 26472
rect 30929 26463 30987 26469
rect 30190 26392 30196 26444
rect 30248 26432 30254 26444
rect 30285 26435 30343 26441
rect 30285 26432 30297 26435
rect 30248 26404 30297 26432
rect 30248 26392 30254 26404
rect 30285 26401 30297 26404
rect 30331 26401 30343 26435
rect 30285 26395 30343 26401
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 28534 26324 28540 26376
rect 28592 26364 28598 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 28592 26336 29745 26364
rect 28592 26324 28598 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 31312 26364 31340 26472
rect 32324 26472 32680 26500
rect 32324 26441 32352 26472
rect 32674 26460 32680 26472
rect 32732 26460 32738 26512
rect 33594 26500 33600 26512
rect 33244 26472 33600 26500
rect 33244 26441 33272 26472
rect 33594 26460 33600 26472
rect 33652 26460 33658 26512
rect 34057 26503 34115 26509
rect 34057 26469 34069 26503
rect 34103 26500 34115 26503
rect 34146 26500 34152 26512
rect 34103 26472 34152 26500
rect 34103 26469 34115 26472
rect 34057 26463 34115 26469
rect 34146 26460 34152 26472
rect 34204 26460 34210 26512
rect 34238 26460 34244 26512
rect 34296 26460 34302 26512
rect 35361 26500 35389 26540
rect 35526 26528 35532 26580
rect 35584 26528 35590 26580
rect 37826 26568 37832 26580
rect 35636 26540 37832 26568
rect 35636 26500 35664 26540
rect 37826 26528 37832 26540
rect 37884 26568 37890 26580
rect 37921 26571 37979 26577
rect 37921 26568 37933 26571
rect 37884 26540 37933 26568
rect 37884 26528 37890 26540
rect 37921 26537 37933 26540
rect 37967 26537 37979 26571
rect 37921 26531 37979 26537
rect 35361 26472 35664 26500
rect 32309 26435 32367 26441
rect 32309 26401 32321 26435
rect 32355 26401 32367 26435
rect 32309 26395 32367 26401
rect 33229 26435 33287 26441
rect 33229 26401 33241 26435
rect 33275 26401 33287 26435
rect 33229 26395 33287 26401
rect 33410 26392 33416 26444
rect 33468 26392 33474 26444
rect 34256 26432 34284 26460
rect 34514 26432 34520 26444
rect 34256 26404 34520 26432
rect 34514 26392 34520 26404
rect 34572 26432 34578 26444
rect 34572 26404 35112 26432
rect 34572 26392 34578 26404
rect 33137 26367 33195 26373
rect 33137 26364 33149 26367
rect 31312 26358 32352 26364
rect 32472 26358 33149 26364
rect 31312 26336 33149 26358
rect 32324 26330 32500 26336
rect 33137 26333 33149 26336
rect 33183 26364 33195 26367
rect 33962 26364 33968 26376
rect 33183 26336 33968 26364
rect 33183 26333 33195 26336
rect 33137 26327 33195 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34054 26324 34060 26376
rect 34112 26324 34118 26376
rect 34238 26324 34244 26376
rect 34296 26324 34302 26376
rect 34974 26324 34980 26376
rect 35032 26324 35038 26376
rect 35084 26373 35112 26404
rect 36354 26392 36360 26444
rect 36412 26432 36418 26444
rect 36541 26435 36599 26441
rect 36541 26432 36553 26435
rect 36412 26404 36553 26432
rect 36412 26392 36418 26404
rect 36541 26401 36553 26404
rect 36587 26401 36599 26435
rect 36541 26395 36599 26401
rect 35069 26367 35127 26373
rect 35069 26333 35081 26367
rect 35115 26333 35127 26367
rect 35069 26327 35127 26333
rect 35250 26324 35256 26376
rect 35308 26324 35314 26376
rect 35342 26324 35348 26376
rect 35400 26324 35406 26376
rect 36814 26373 36820 26376
rect 36808 26364 36820 26373
rect 36775 26336 36820 26364
rect 36808 26327 36820 26336
rect 36814 26324 36820 26327
rect 36872 26324 36878 26376
rect 29546 26296 29552 26308
rect 27724 26268 29552 26296
rect 29546 26256 29552 26268
rect 29604 26256 29610 26308
rect 32064 26299 32122 26305
rect 32064 26265 32076 26299
rect 32110 26296 32122 26299
rect 32110 26268 32449 26296
rect 32110 26265 32122 26268
rect 32064 26259 32122 26265
rect 22428 26200 22600 26228
rect 22428 26188 22434 26200
rect 22922 26188 22928 26240
rect 22980 26228 22986 26240
rect 23017 26231 23075 26237
rect 23017 26228 23029 26231
rect 22980 26200 23029 26228
rect 22980 26188 22986 26200
rect 23017 26197 23029 26200
rect 23063 26197 23075 26231
rect 23017 26191 23075 26197
rect 30190 26188 30196 26240
rect 30248 26188 30254 26240
rect 32421 26228 32449 26268
rect 32769 26231 32827 26237
rect 32769 26228 32781 26231
rect 32421 26200 32781 26228
rect 32769 26197 32781 26200
rect 32815 26197 32827 26231
rect 32769 26191 32827 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 4890 25984 4896 26036
rect 4948 26024 4954 26036
rect 5629 26027 5687 26033
rect 5629 26024 5641 26027
rect 4948 25996 5641 26024
rect 4948 25984 4954 25996
rect 5629 25993 5641 25996
rect 5675 26024 5687 26027
rect 6914 26024 6920 26036
rect 5675 25996 6920 26024
rect 5675 25993 5687 25996
rect 5629 25987 5687 25993
rect 6914 25984 6920 25996
rect 6972 25984 6978 26036
rect 10594 25984 10600 26036
rect 10652 25984 10658 26036
rect 11146 25984 11152 26036
rect 11204 25984 11210 26036
rect 12805 26027 12863 26033
rect 12805 25993 12817 26027
rect 12851 26024 12863 26027
rect 14090 26024 14096 26036
rect 12851 25996 14096 26024
rect 12851 25993 12863 25996
rect 12805 25987 12863 25993
rect 5258 25916 5264 25968
rect 5316 25956 5322 25968
rect 6733 25959 6791 25965
rect 6733 25956 6745 25959
rect 5316 25928 6745 25956
rect 5316 25916 5322 25928
rect 6733 25925 6745 25928
rect 6779 25925 6791 25959
rect 6733 25919 6791 25925
rect 9677 25959 9735 25965
rect 9677 25925 9689 25959
rect 9723 25956 9735 25959
rect 10612 25956 10640 25984
rect 9723 25928 10640 25956
rect 9723 25925 9735 25928
rect 9677 25919 9735 25925
rect 12250 25916 12256 25968
rect 12308 25956 12314 25968
rect 12434 25956 12440 25968
rect 12308 25928 12440 25956
rect 12308 25916 12314 25928
rect 12434 25916 12440 25928
rect 12492 25916 12498 25968
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 5445 25891 5503 25897
rect 5445 25888 5457 25891
rect 4856 25860 5457 25888
rect 4856 25848 4862 25860
rect 5445 25857 5457 25860
rect 5491 25888 5503 25891
rect 5534 25888 5540 25900
rect 5491 25860 5540 25888
rect 5491 25857 5503 25860
rect 5445 25851 5503 25857
rect 5534 25848 5540 25860
rect 5592 25848 5598 25900
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 5810 25888 5816 25900
rect 5767 25860 5816 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 5810 25848 5816 25860
rect 5868 25848 5874 25900
rect 6638 25848 6644 25900
rect 6696 25848 6702 25900
rect 6822 25848 6828 25900
rect 6880 25888 6886 25900
rect 7282 25888 7288 25900
rect 6880 25860 7288 25888
rect 6880 25848 6886 25860
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 8110 25848 8116 25900
rect 8168 25848 8174 25900
rect 8570 25848 8576 25900
rect 8628 25888 8634 25900
rect 9490 25888 9496 25900
rect 8628 25860 9496 25888
rect 8628 25848 8634 25860
rect 9490 25848 9496 25860
rect 9548 25888 9554 25900
rect 9953 25891 10011 25897
rect 9953 25888 9965 25891
rect 9548 25860 9965 25888
rect 9548 25848 9554 25860
rect 9953 25857 9965 25860
rect 9999 25857 10011 25891
rect 9953 25851 10011 25857
rect 5166 25780 5172 25832
rect 5224 25820 5230 25832
rect 5261 25823 5319 25829
rect 5261 25820 5273 25823
rect 5224 25792 5273 25820
rect 5224 25780 5230 25792
rect 5261 25789 5273 25792
rect 5307 25789 5319 25823
rect 5261 25783 5319 25789
rect 5353 25823 5411 25829
rect 5353 25789 5365 25823
rect 5399 25820 5411 25823
rect 5902 25820 5908 25832
rect 5399 25792 5908 25820
rect 5399 25789 5411 25792
rect 5353 25783 5411 25789
rect 5902 25780 5908 25792
rect 5960 25820 5966 25832
rect 8205 25823 8263 25829
rect 8205 25820 8217 25823
rect 5960 25792 8217 25820
rect 5960 25780 5966 25792
rect 8205 25789 8217 25792
rect 8251 25820 8263 25823
rect 9398 25820 9404 25832
rect 8251 25792 9404 25820
rect 8251 25789 8263 25792
rect 8205 25783 8263 25789
rect 9398 25780 9404 25792
rect 9456 25780 9462 25832
rect 9766 25780 9772 25832
rect 9824 25780 9830 25832
rect 5810 25712 5816 25764
rect 5868 25752 5874 25764
rect 6638 25752 6644 25764
rect 5868 25724 6644 25752
rect 5868 25712 5874 25724
rect 6638 25712 6644 25724
rect 6696 25752 6702 25764
rect 8294 25752 8300 25764
rect 6696 25724 8300 25752
rect 6696 25712 6702 25724
rect 8294 25712 8300 25724
rect 8352 25712 8358 25764
rect 9968 25752 9996 25851
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10410 25888 10416 25900
rect 10284 25860 10416 25888
rect 10284 25848 10290 25860
rect 10410 25848 10416 25860
rect 10468 25888 10474 25900
rect 10597 25891 10655 25897
rect 10597 25888 10609 25891
rect 10468 25860 10609 25888
rect 10468 25848 10474 25860
rect 10597 25857 10609 25860
rect 10643 25857 10655 25891
rect 10597 25851 10655 25857
rect 10686 25848 10692 25900
rect 10744 25888 10750 25900
rect 10781 25891 10839 25897
rect 10781 25888 10793 25891
rect 10744 25860 10793 25888
rect 10744 25848 10750 25860
rect 10781 25857 10793 25860
rect 10827 25857 10839 25891
rect 10781 25851 10839 25857
rect 10873 25891 10931 25897
rect 10873 25857 10885 25891
rect 10919 25857 10931 25891
rect 10873 25851 10931 25857
rect 10888 25820 10916 25851
rect 10962 25848 10968 25900
rect 11020 25848 11026 25900
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 12526 25820 12532 25832
rect 10888 25792 12532 25820
rect 12526 25780 12532 25792
rect 12584 25780 12590 25832
rect 11974 25752 11980 25764
rect 9968 25724 11980 25752
rect 11974 25712 11980 25724
rect 12032 25712 12038 25764
rect 4890 25644 4896 25696
rect 4948 25684 4954 25696
rect 4985 25687 5043 25693
rect 4985 25684 4997 25687
rect 4948 25656 4997 25684
rect 4948 25644 4954 25656
rect 4985 25653 4997 25656
rect 5031 25653 5043 25687
rect 4985 25647 5043 25653
rect 9950 25644 9956 25696
rect 10008 25644 10014 25696
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25684 10195 25687
rect 10226 25684 10232 25696
rect 10183 25656 10232 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 10226 25644 10232 25656
rect 10284 25644 10290 25696
rect 10318 25644 10324 25696
rect 10376 25684 10382 25696
rect 12820 25684 12848 25987
rect 14090 25984 14096 25996
rect 14148 25984 14154 26036
rect 17313 26027 17371 26033
rect 17313 25993 17325 26027
rect 17359 26024 17371 26027
rect 18046 26024 18052 26036
rect 17359 25996 18052 26024
rect 17359 25993 17371 25996
rect 17313 25987 17371 25993
rect 18046 25984 18052 25996
rect 18104 25984 18110 26036
rect 19886 25984 19892 26036
rect 19944 26024 19950 26036
rect 20441 26027 20499 26033
rect 20441 26024 20453 26027
rect 19944 25996 20453 26024
rect 19944 25984 19950 25996
rect 20441 25993 20453 25996
rect 20487 25993 20499 26027
rect 20441 25987 20499 25993
rect 21358 25984 21364 26036
rect 21416 26024 21422 26036
rect 21416 25996 22600 26024
rect 21416 25984 21422 25996
rect 16942 25916 16948 25968
rect 17000 25956 17006 25968
rect 17037 25959 17095 25965
rect 17037 25956 17049 25959
rect 17000 25928 17049 25956
rect 17000 25916 17006 25928
rect 17037 25925 17049 25928
rect 17083 25925 17095 25959
rect 17037 25919 17095 25925
rect 17405 25959 17463 25965
rect 17405 25925 17417 25959
rect 17451 25956 17463 25959
rect 19334 25956 19340 25968
rect 17451 25928 19340 25956
rect 17451 25925 17463 25928
rect 17405 25919 17463 25925
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 20254 25916 20260 25968
rect 20312 25916 20318 25968
rect 20714 25916 20720 25968
rect 20772 25956 20778 25968
rect 21726 25956 21732 25968
rect 20772 25928 21732 25956
rect 20772 25916 20778 25928
rect 21726 25916 21732 25928
rect 21784 25956 21790 25968
rect 21784 25928 22232 25956
rect 21784 25916 21790 25928
rect 12986 25848 12992 25900
rect 13044 25848 13050 25900
rect 13630 25848 13636 25900
rect 13688 25888 13694 25900
rect 14093 25891 14151 25897
rect 14093 25888 14105 25891
rect 13688 25860 14105 25888
rect 13688 25848 13694 25860
rect 14093 25857 14105 25860
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 14369 25891 14427 25897
rect 14369 25857 14381 25891
rect 14415 25888 14427 25891
rect 15194 25888 15200 25900
rect 14415 25860 15200 25888
rect 14415 25857 14427 25860
rect 14369 25851 14427 25857
rect 15194 25848 15200 25860
rect 15252 25848 15258 25900
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25888 17279 25891
rect 17678 25888 17684 25900
rect 17267 25860 17684 25888
rect 17267 25857 17279 25860
rect 17221 25851 17279 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 18138 25848 18144 25900
rect 18196 25848 18202 25900
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 20272 25888 20300 25916
rect 18647 25860 20300 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 22002 25848 22008 25900
rect 22060 25888 22066 25900
rect 22094 25888 22100 25900
rect 22060 25860 22100 25888
rect 22060 25848 22066 25860
rect 22094 25848 22100 25860
rect 22152 25848 22158 25900
rect 22204 25897 22232 25928
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 17310 25780 17316 25832
rect 17368 25820 17374 25832
rect 17770 25820 17776 25832
rect 17368 25792 17776 25820
rect 17368 25780 17374 25792
rect 17770 25780 17776 25792
rect 17828 25820 17834 25832
rect 18509 25823 18567 25829
rect 18509 25820 18521 25823
rect 17828 25792 18521 25820
rect 17828 25780 17834 25792
rect 18509 25789 18521 25792
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 20070 25780 20076 25832
rect 20128 25780 20134 25832
rect 20165 25823 20223 25829
rect 20165 25789 20177 25823
rect 20211 25820 20223 25823
rect 20806 25820 20812 25832
rect 20211 25792 20812 25820
rect 20211 25789 20223 25792
rect 20165 25783 20223 25789
rect 17494 25712 17500 25764
rect 17552 25752 17558 25764
rect 17552 25724 17908 25752
rect 17552 25712 17558 25724
rect 10376 25656 12848 25684
rect 10376 25644 10382 25656
rect 13170 25644 13176 25696
rect 13228 25644 13234 25696
rect 17589 25687 17647 25693
rect 17589 25653 17601 25687
rect 17635 25684 17647 25687
rect 17770 25684 17776 25696
rect 17635 25656 17776 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 17770 25644 17776 25656
rect 17828 25644 17834 25696
rect 17880 25684 17908 25724
rect 18138 25712 18144 25764
rect 18196 25752 18202 25764
rect 20180 25752 20208 25783
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 22572 25829 22600 25996
rect 26234 25984 26240 26036
rect 26292 26024 26298 26036
rect 31205 26027 31263 26033
rect 26292 25996 28028 26024
rect 26292 25984 26298 25996
rect 22738 25916 22744 25968
rect 22796 25956 22802 25968
rect 27614 25956 27620 25968
rect 22796 25928 27620 25956
rect 22796 25916 22802 25928
rect 27614 25916 27620 25928
rect 27672 25916 27678 25968
rect 27890 25916 27896 25968
rect 27948 25916 27954 25968
rect 23290 25848 23296 25900
rect 23348 25848 23354 25900
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25888 23627 25891
rect 23750 25888 23756 25900
rect 23615 25860 23756 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 23750 25848 23756 25860
rect 23808 25888 23814 25900
rect 25130 25888 25136 25900
rect 23808 25860 25136 25888
rect 23808 25848 23814 25860
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 27706 25848 27712 25900
rect 27764 25848 27770 25900
rect 27801 25891 27859 25897
rect 27801 25857 27813 25891
rect 27847 25888 27859 25891
rect 27847 25860 27936 25888
rect 27847 25857 27859 25860
rect 27801 25851 27859 25857
rect 22557 25823 22615 25829
rect 22557 25789 22569 25823
rect 22603 25820 22615 25823
rect 24854 25820 24860 25832
rect 22603 25792 24860 25820
rect 22603 25789 22615 25792
rect 22557 25783 22615 25789
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 18196 25724 20208 25752
rect 18196 25712 18202 25724
rect 23290 25712 23296 25764
rect 23348 25712 23354 25764
rect 20898 25684 20904 25696
rect 17880 25656 20904 25684
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 27522 25644 27528 25696
rect 27580 25644 27586 25696
rect 27908 25684 27936 25860
rect 28000 25752 28028 25996
rect 31205 25993 31217 26027
rect 31251 26024 31263 26027
rect 32398 26024 32404 26036
rect 31251 25996 32404 26024
rect 31251 25993 31263 25996
rect 31205 25987 31263 25993
rect 32398 25984 32404 25996
rect 32456 25984 32462 26036
rect 33686 25984 33692 26036
rect 33744 26024 33750 26036
rect 34517 26027 34575 26033
rect 33744 25996 34376 26024
rect 33744 25984 33750 25996
rect 28994 25916 29000 25968
rect 29052 25916 29058 25968
rect 33134 25916 33140 25968
rect 33192 25956 33198 25968
rect 34241 25959 34299 25965
rect 34241 25956 34253 25959
rect 33192 25928 34253 25956
rect 33192 25916 33198 25928
rect 34241 25925 34253 25928
rect 34287 25925 34299 25959
rect 34241 25919 34299 25925
rect 28077 25891 28135 25897
rect 28077 25857 28089 25891
rect 28123 25888 28135 25891
rect 29454 25888 29460 25900
rect 28123 25860 29460 25888
rect 28123 25857 28135 25860
rect 28077 25851 28135 25857
rect 29454 25848 29460 25860
rect 29512 25848 29518 25900
rect 30190 25848 30196 25900
rect 30248 25848 30254 25900
rect 30650 25848 30656 25900
rect 30708 25848 30714 25900
rect 30742 25848 30748 25900
rect 30800 25848 30806 25900
rect 30929 25891 30987 25897
rect 30929 25857 30941 25891
rect 30975 25857 30987 25891
rect 30929 25851 30987 25857
rect 30282 25780 30288 25832
rect 30340 25820 30346 25832
rect 30944 25820 30972 25851
rect 31018 25848 31024 25900
rect 31076 25848 31082 25900
rect 33870 25848 33876 25900
rect 33928 25888 33934 25900
rect 34348 25897 34376 25996
rect 34517 25993 34529 26027
rect 34563 26024 34575 26027
rect 34974 26024 34980 26036
rect 34563 25996 34980 26024
rect 34563 25993 34575 25996
rect 34517 25987 34575 25993
rect 34974 25984 34980 25996
rect 35032 25984 35038 26036
rect 36262 25916 36268 25968
rect 36320 25956 36326 25968
rect 36366 25959 36424 25965
rect 36366 25956 36378 25959
rect 36320 25928 36378 25956
rect 36320 25916 36326 25928
rect 36366 25925 36378 25928
rect 36412 25925 36424 25959
rect 36366 25919 36424 25925
rect 33965 25891 34023 25897
rect 33965 25888 33977 25891
rect 33928 25860 33977 25888
rect 33928 25848 33934 25860
rect 33965 25857 33977 25860
rect 34011 25857 34023 25891
rect 33965 25851 34023 25857
rect 34149 25891 34207 25897
rect 34149 25857 34161 25891
rect 34195 25857 34207 25891
rect 34149 25851 34207 25857
rect 34333 25891 34391 25897
rect 34333 25857 34345 25891
rect 34379 25857 34391 25891
rect 34333 25851 34391 25857
rect 37829 25891 37887 25897
rect 37829 25857 37841 25891
rect 37875 25888 37887 25891
rect 37918 25888 37924 25900
rect 37875 25860 37924 25888
rect 37875 25857 37887 25860
rect 37829 25851 37887 25857
rect 31662 25820 31668 25832
rect 30340 25792 31668 25820
rect 30340 25780 30346 25792
rect 31662 25780 31668 25792
rect 31720 25780 31726 25832
rect 33778 25780 33784 25832
rect 33836 25820 33842 25832
rect 34164 25820 34192 25851
rect 37918 25848 37924 25860
rect 37976 25848 37982 25900
rect 33836 25792 34192 25820
rect 36633 25823 36691 25829
rect 33836 25780 33842 25792
rect 36633 25789 36645 25823
rect 36679 25820 36691 25823
rect 36722 25820 36728 25832
rect 36679 25792 36728 25820
rect 36679 25789 36691 25792
rect 36633 25783 36691 25789
rect 36722 25780 36728 25792
rect 36780 25780 36786 25832
rect 38105 25823 38163 25829
rect 38105 25789 38117 25823
rect 38151 25820 38163 25823
rect 39022 25820 39028 25832
rect 38151 25792 39028 25820
rect 38151 25789 38163 25792
rect 38105 25783 38163 25789
rect 39022 25780 39028 25792
rect 39080 25780 39086 25832
rect 32030 25752 32036 25764
rect 28000 25724 32036 25752
rect 32030 25712 32036 25724
rect 32088 25712 32094 25764
rect 30742 25684 30748 25696
rect 27908 25656 30748 25684
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 33410 25644 33416 25696
rect 33468 25684 33474 25696
rect 35253 25687 35311 25693
rect 35253 25684 35265 25687
rect 33468 25656 35265 25684
rect 33468 25644 33474 25656
rect 35253 25653 35265 25656
rect 35299 25653 35311 25687
rect 35253 25647 35311 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 5626 25440 5632 25492
rect 5684 25480 5690 25492
rect 6549 25483 6607 25489
rect 6549 25480 6561 25483
rect 5684 25452 6561 25480
rect 5684 25440 5690 25452
rect 6549 25449 6561 25452
rect 6595 25449 6607 25483
rect 6549 25443 6607 25449
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 9306 25480 9312 25492
rect 6972 25452 9312 25480
rect 6972 25440 6978 25452
rect 9306 25440 9312 25452
rect 9364 25480 9370 25492
rect 9493 25483 9551 25489
rect 9493 25480 9505 25483
rect 9364 25452 9505 25480
rect 9364 25440 9370 25452
rect 9493 25449 9505 25452
rect 9539 25449 9551 25483
rect 9493 25443 9551 25449
rect 12986 25440 12992 25492
rect 13044 25480 13050 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 13044 25452 14289 25480
rect 13044 25440 13050 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 17678 25440 17684 25492
rect 17736 25480 17742 25492
rect 24302 25480 24308 25492
rect 17736 25452 24308 25480
rect 17736 25440 17742 25452
rect 24302 25440 24308 25452
rect 24360 25440 24366 25492
rect 25225 25483 25283 25489
rect 25225 25449 25237 25483
rect 25271 25480 25283 25483
rect 25314 25480 25320 25492
rect 25271 25452 25320 25480
rect 25271 25449 25283 25452
rect 25225 25443 25283 25449
rect 25314 25440 25320 25452
rect 25372 25440 25378 25492
rect 28074 25440 28080 25492
rect 28132 25480 28138 25492
rect 28132 25452 29960 25480
rect 28132 25440 28138 25452
rect 4341 25415 4399 25421
rect 4341 25381 4353 25415
rect 4387 25412 4399 25415
rect 5074 25412 5080 25424
rect 4387 25384 5080 25412
rect 4387 25381 4399 25384
rect 4341 25375 4399 25381
rect 5074 25372 5080 25384
rect 5132 25412 5138 25424
rect 10318 25412 10324 25424
rect 5132 25384 10324 25412
rect 5132 25372 5138 25384
rect 10318 25372 10324 25384
rect 10376 25372 10382 25424
rect 18601 25415 18659 25421
rect 18601 25412 18613 25415
rect 13372 25384 18613 25412
rect 4614 25344 4620 25356
rect 4172 25316 4620 25344
rect 4172 25285 4200 25316
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 4890 25304 4896 25356
rect 4948 25304 4954 25356
rect 5258 25304 5264 25356
rect 5316 25304 5322 25356
rect 5350 25304 5356 25356
rect 5408 25304 5414 25356
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7561 25347 7619 25353
rect 7561 25344 7573 25347
rect 6871 25316 7573 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 7561 25313 7573 25316
rect 7607 25313 7619 25347
rect 7561 25307 7619 25313
rect 8202 25304 8208 25356
rect 8260 25344 8266 25356
rect 10134 25344 10140 25356
rect 8260 25316 10140 25344
rect 8260 25304 8266 25316
rect 10134 25304 10140 25316
rect 10192 25304 10198 25356
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 4433 25279 4491 25285
rect 4433 25245 4445 25279
rect 4479 25276 4491 25279
rect 4479 25248 4660 25276
rect 4479 25245 4491 25248
rect 4433 25239 4491 25245
rect 4632 25220 4660 25248
rect 4614 25168 4620 25220
rect 4672 25168 4678 25220
rect 5276 25208 5304 25304
rect 6730 25236 6736 25288
rect 6788 25236 6794 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 7009 25279 7067 25285
rect 7009 25245 7021 25279
rect 7055 25276 7067 25279
rect 9674 25276 9680 25288
rect 7055 25248 9680 25276
rect 7055 25245 7067 25248
rect 7009 25239 7067 25245
rect 6932 25208 6960 25239
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25276 9827 25279
rect 10594 25276 10600 25288
rect 9815 25248 10600 25276
rect 9815 25245 9827 25248
rect 9769 25239 9827 25245
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 12342 25236 12348 25288
rect 12400 25236 12406 25288
rect 12612 25279 12670 25285
rect 12612 25245 12624 25279
rect 12658 25276 12670 25279
rect 13170 25276 13176 25288
rect 12658 25248 13176 25276
rect 12658 25245 12670 25248
rect 12612 25239 12670 25245
rect 13170 25236 13176 25248
rect 13228 25236 13234 25288
rect 5276 25180 6960 25208
rect 7745 25211 7803 25217
rect 7745 25177 7757 25211
rect 7791 25208 7803 25211
rect 7834 25208 7840 25220
rect 7791 25180 7840 25208
rect 7791 25177 7803 25180
rect 7745 25171 7803 25177
rect 7834 25168 7840 25180
rect 7892 25168 7898 25220
rect 7929 25211 7987 25217
rect 7929 25177 7941 25211
rect 7975 25208 7987 25211
rect 8202 25208 8208 25220
rect 7975 25180 8208 25208
rect 7975 25177 7987 25180
rect 7929 25171 7987 25177
rect 8202 25168 8208 25180
rect 8260 25168 8266 25220
rect 8294 25168 8300 25220
rect 8352 25208 8358 25220
rect 9309 25211 9367 25217
rect 9309 25208 9321 25211
rect 8352 25180 9321 25208
rect 8352 25168 8358 25180
rect 9309 25177 9321 25180
rect 9355 25208 9367 25211
rect 9950 25208 9956 25220
rect 9355 25180 9956 25208
rect 9355 25177 9367 25180
rect 9309 25171 9367 25177
rect 9950 25168 9956 25180
rect 10008 25168 10014 25220
rect 12526 25168 12532 25220
rect 12584 25208 12590 25220
rect 13372 25208 13400 25384
rect 18601 25381 18613 25384
rect 18647 25381 18659 25415
rect 18601 25375 18659 25381
rect 19886 25372 19892 25424
rect 19944 25412 19950 25424
rect 20070 25412 20076 25424
rect 19944 25384 20076 25412
rect 19944 25372 19950 25384
rect 20070 25372 20076 25384
rect 20128 25372 20134 25424
rect 24854 25372 24860 25424
rect 24912 25412 24918 25424
rect 25498 25412 25504 25424
rect 24912 25384 25504 25412
rect 24912 25372 24918 25384
rect 25498 25372 25504 25384
rect 25556 25412 25562 25424
rect 27706 25412 27712 25424
rect 25556 25384 27712 25412
rect 25556 25372 25562 25384
rect 13630 25304 13636 25356
rect 13688 25344 13694 25356
rect 16669 25347 16727 25353
rect 13688 25316 14780 25344
rect 13688 25304 13694 25316
rect 13446 25236 13452 25288
rect 13504 25276 13510 25288
rect 14752 25285 14780 25316
rect 16669 25313 16681 25347
rect 16715 25344 16727 25347
rect 18046 25344 18052 25356
rect 16715 25316 18052 25344
rect 16715 25313 16727 25316
rect 16669 25307 16727 25313
rect 18046 25304 18052 25316
rect 18104 25304 18110 25356
rect 18322 25304 18328 25356
rect 18380 25344 18386 25356
rect 19058 25344 19064 25356
rect 18380 25316 19064 25344
rect 18380 25304 18386 25316
rect 19058 25304 19064 25316
rect 19116 25344 19122 25356
rect 19429 25347 19487 25353
rect 19429 25344 19441 25347
rect 19116 25316 19441 25344
rect 19116 25304 19122 25316
rect 19429 25313 19441 25316
rect 19475 25313 19487 25347
rect 20254 25344 20260 25356
rect 19429 25307 19487 25313
rect 19628 25316 20260 25344
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 13504 25248 14473 25276
rect 13504 25236 13510 25248
rect 14461 25245 14473 25248
rect 14507 25245 14519 25279
rect 14461 25239 14519 25245
rect 14737 25279 14795 25285
rect 14737 25245 14749 25279
rect 14783 25276 14795 25279
rect 15746 25276 15752 25288
rect 14783 25248 15752 25276
rect 14783 25245 14795 25248
rect 14737 25239 14795 25245
rect 15746 25236 15752 25248
rect 15804 25236 15810 25288
rect 16114 25236 16120 25288
rect 16172 25236 16178 25288
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 14645 25211 14703 25217
rect 14645 25208 14657 25211
rect 12584 25180 13400 25208
rect 13740 25180 14657 25208
rect 12584 25168 12590 25180
rect 3970 25100 3976 25152
rect 4028 25100 4034 25152
rect 5534 25100 5540 25152
rect 5592 25100 5598 25152
rect 7098 25100 7104 25152
rect 7156 25140 7162 25152
rect 8478 25140 8484 25152
rect 7156 25112 8484 25140
rect 7156 25100 7162 25112
rect 8478 25100 8484 25112
rect 8536 25140 8542 25152
rect 13740 25149 13768 25180
rect 14645 25177 14657 25180
rect 14691 25208 14703 25211
rect 16224 25208 16252 25239
rect 16574 25236 16580 25288
rect 16632 25236 16638 25288
rect 18138 25236 18144 25288
rect 18196 25276 18202 25288
rect 18233 25279 18291 25285
rect 18233 25276 18245 25279
rect 18196 25248 18245 25276
rect 18196 25236 18202 25248
rect 18233 25245 18245 25248
rect 18279 25245 18291 25279
rect 18417 25279 18475 25285
rect 18417 25276 18429 25279
rect 18233 25239 18291 25245
rect 18340 25248 18429 25276
rect 14691 25180 16252 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 16758 25168 16764 25220
rect 16816 25208 16822 25220
rect 17221 25211 17279 25217
rect 17221 25208 17233 25211
rect 16816 25180 17233 25208
rect 16816 25168 16822 25180
rect 17221 25177 17233 25180
rect 17267 25177 17279 25211
rect 17221 25171 17279 25177
rect 9493 25143 9551 25149
rect 9493 25140 9505 25143
rect 8536 25112 9505 25140
rect 8536 25100 8542 25112
rect 9493 25109 9505 25112
rect 9539 25109 9551 25143
rect 9493 25103 9551 25109
rect 13725 25143 13783 25149
rect 13725 25109 13737 25143
rect 13771 25109 13783 25143
rect 13725 25103 13783 25109
rect 13998 25100 14004 25152
rect 14056 25140 14062 25152
rect 18340 25140 18368 25248
rect 18417 25245 18429 25248
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18506 25236 18512 25288
rect 18564 25236 18570 25288
rect 18690 25236 18696 25288
rect 18748 25236 18754 25288
rect 19628 25285 19656 25316
rect 20254 25304 20260 25316
rect 20312 25304 20318 25356
rect 24486 25344 24492 25356
rect 20364 25316 24492 25344
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20364 25276 20392 25316
rect 24486 25304 24492 25316
rect 24544 25304 24550 25356
rect 26206 25344 26234 25384
rect 27706 25372 27712 25384
rect 27764 25372 27770 25424
rect 28534 25372 28540 25424
rect 28592 25412 28598 25424
rect 28721 25415 28779 25421
rect 28721 25412 28733 25415
rect 28592 25384 28733 25412
rect 28592 25372 28598 25384
rect 28721 25381 28733 25384
rect 28767 25381 28779 25415
rect 28721 25375 28779 25381
rect 29932 25353 29960 25452
rect 32585 25415 32643 25421
rect 32585 25381 32597 25415
rect 32631 25412 32643 25415
rect 32631 25384 33088 25412
rect 32631 25381 32643 25384
rect 32585 25375 32643 25381
rect 26160 25316 26234 25344
rect 27433 25347 27491 25353
rect 20036 25248 20392 25276
rect 20036 25236 20042 25248
rect 20530 25236 20536 25288
rect 20588 25236 20594 25288
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25276 21051 25279
rect 21174 25276 21180 25288
rect 21039 25248 21180 25276
rect 21039 25245 21051 25248
rect 20993 25239 21051 25245
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 23106 25236 23112 25288
rect 23164 25236 23170 25288
rect 23566 25236 23572 25288
rect 23624 25236 23630 25288
rect 25130 25236 25136 25288
rect 25188 25236 25194 25288
rect 26160 25285 26188 25316
rect 27433 25313 27445 25347
rect 27479 25344 27491 25347
rect 28629 25347 28687 25353
rect 28629 25344 28641 25347
rect 27479 25316 28641 25344
rect 27479 25313 27491 25316
rect 27433 25307 27491 25313
rect 28629 25313 28641 25316
rect 28675 25344 28687 25347
rect 29917 25347 29975 25353
rect 28675 25316 28948 25344
rect 28675 25313 28687 25316
rect 28629 25307 28687 25313
rect 26145 25279 26203 25285
rect 26145 25245 26157 25279
rect 26191 25245 26203 25279
rect 26145 25239 26203 25245
rect 26234 25236 26240 25288
rect 26292 25236 26298 25288
rect 26510 25236 26516 25288
rect 26568 25236 26574 25288
rect 26878 25236 26884 25288
rect 26936 25276 26942 25288
rect 27065 25279 27123 25285
rect 27065 25276 27077 25279
rect 26936 25248 27077 25276
rect 26936 25236 26942 25248
rect 27065 25245 27077 25248
rect 27111 25245 27123 25279
rect 27065 25239 27123 25245
rect 27246 25236 27252 25288
rect 27304 25236 27310 25288
rect 28074 25236 28080 25288
rect 28132 25276 28138 25288
rect 28537 25279 28595 25285
rect 28537 25276 28549 25279
rect 28132 25248 28549 25276
rect 28132 25236 28138 25248
rect 28537 25245 28549 25248
rect 28583 25245 28595 25279
rect 28537 25239 28595 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25245 28871 25279
rect 28920 25276 28948 25316
rect 29917 25313 29929 25347
rect 29963 25313 29975 25347
rect 29917 25307 29975 25313
rect 30377 25347 30435 25353
rect 30377 25313 30389 25347
rect 30423 25344 30435 25347
rect 30558 25344 30564 25356
rect 30423 25316 30564 25344
rect 30423 25313 30435 25316
rect 30377 25307 30435 25313
rect 30558 25304 30564 25316
rect 30616 25344 30622 25356
rect 31018 25344 31024 25356
rect 30616 25316 31024 25344
rect 30616 25304 30622 25316
rect 31018 25304 31024 25316
rect 31076 25344 31082 25356
rect 31076 25316 32260 25344
rect 31076 25304 31082 25316
rect 30009 25279 30067 25285
rect 30009 25276 30021 25279
rect 28920 25248 30021 25276
rect 28813 25239 28871 25245
rect 30009 25245 30021 25248
rect 30055 25245 30067 25279
rect 30009 25239 30067 25245
rect 19889 25211 19947 25217
rect 19889 25177 19901 25211
rect 19935 25208 19947 25211
rect 20898 25208 20904 25220
rect 19935 25180 20904 25208
rect 19935 25177 19947 25180
rect 19889 25171 19947 25177
rect 20898 25168 20904 25180
rect 20956 25168 20962 25220
rect 24946 25168 24952 25220
rect 25004 25168 25010 25220
rect 26329 25211 26387 25217
rect 26329 25208 26341 25211
rect 25792 25180 26341 25208
rect 14056 25112 18368 25140
rect 18877 25143 18935 25149
rect 14056 25100 14062 25112
rect 18877 25109 18889 25143
rect 18923 25140 18935 25143
rect 19426 25140 19432 25152
rect 18923 25112 19432 25140
rect 18923 25109 18935 25112
rect 18877 25103 18935 25109
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 20622 25100 20628 25152
rect 20680 25140 20686 25152
rect 20717 25143 20775 25149
rect 20717 25140 20729 25143
rect 20680 25112 20729 25140
rect 20680 25100 20686 25112
rect 20717 25109 20729 25112
rect 20763 25109 20775 25143
rect 20717 25103 20775 25109
rect 22094 25100 22100 25152
rect 22152 25140 22158 25152
rect 22649 25143 22707 25149
rect 22649 25140 22661 25143
rect 22152 25112 22661 25140
rect 22152 25100 22158 25112
rect 22649 25109 22661 25112
rect 22695 25109 22707 25143
rect 22649 25103 22707 25109
rect 24118 25100 24124 25152
rect 24176 25140 24182 25152
rect 25792 25140 25820 25180
rect 26329 25177 26341 25180
rect 26375 25208 26387 25211
rect 28626 25208 28632 25220
rect 26375 25180 28632 25208
rect 26375 25177 26387 25180
rect 26329 25171 26387 25177
rect 28626 25168 28632 25180
rect 28684 25168 28690 25220
rect 28828 25208 28856 25239
rect 31846 25236 31852 25288
rect 31904 25276 31910 25288
rect 31941 25279 31999 25285
rect 31941 25276 31953 25279
rect 31904 25248 31953 25276
rect 31904 25236 31910 25248
rect 31941 25245 31953 25248
rect 31987 25245 31999 25279
rect 31941 25239 31999 25245
rect 32030 25236 32036 25288
rect 32088 25276 32094 25288
rect 32232 25276 32260 25316
rect 32306 25304 32312 25356
rect 32364 25344 32370 25356
rect 33060 25353 33088 25384
rect 33045 25347 33103 25353
rect 32364 25316 32536 25344
rect 32364 25304 32370 25316
rect 32406 25279 32464 25285
rect 32406 25276 32418 25279
rect 32088 25248 32133 25276
rect 32232 25248 32418 25276
rect 32088 25236 32094 25248
rect 32406 25245 32418 25248
rect 32452 25245 32464 25279
rect 32508 25276 32536 25316
rect 33045 25313 33057 25347
rect 33091 25313 33103 25347
rect 33045 25307 33103 25313
rect 33410 25276 33416 25288
rect 32508 25248 33416 25276
rect 32406 25239 32464 25245
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 33594 25236 33600 25288
rect 33652 25236 33658 25288
rect 34790 25236 34796 25288
rect 34848 25276 34854 25288
rect 34977 25279 35035 25285
rect 34977 25276 34989 25279
rect 34848 25248 34989 25276
rect 34848 25236 34854 25248
rect 34977 25245 34989 25248
rect 35023 25245 35035 25279
rect 34977 25239 35035 25245
rect 35805 25279 35863 25285
rect 35805 25245 35817 25279
rect 35851 25276 35863 25279
rect 36633 25279 36691 25285
rect 36633 25276 36645 25279
rect 35851 25248 36645 25276
rect 35851 25245 35863 25248
rect 35805 25239 35863 25245
rect 36633 25245 36645 25248
rect 36679 25276 36691 25279
rect 36722 25276 36728 25288
rect 36679 25248 36728 25276
rect 36679 25245 36691 25248
rect 36633 25239 36691 25245
rect 36722 25236 36728 25248
rect 36780 25236 36786 25288
rect 30098 25208 30104 25220
rect 28828 25180 30104 25208
rect 30098 25168 30104 25180
rect 30156 25168 30162 25220
rect 30282 25168 30288 25220
rect 30340 25168 30346 25220
rect 32214 25168 32220 25220
rect 32272 25168 32278 25220
rect 32309 25211 32367 25217
rect 32309 25177 32321 25211
rect 32355 25208 32367 25211
rect 32490 25208 32496 25220
rect 32355 25180 32496 25208
rect 32355 25177 32367 25180
rect 32309 25171 32367 25177
rect 32490 25168 32496 25180
rect 32548 25168 32554 25220
rect 36900 25211 36958 25217
rect 36900 25177 36912 25211
rect 36946 25208 36958 25211
rect 37458 25208 37464 25220
rect 36946 25180 37464 25208
rect 36946 25177 36958 25180
rect 36900 25171 36958 25177
rect 37458 25168 37464 25180
rect 37516 25168 37522 25220
rect 24176 25112 25820 25140
rect 24176 25100 24182 25112
rect 25958 25100 25964 25152
rect 26016 25100 26022 25152
rect 28994 25100 29000 25152
rect 29052 25100 29058 25152
rect 29733 25143 29791 25149
rect 29733 25109 29745 25143
rect 29779 25140 29791 25143
rect 31938 25140 31944 25152
rect 29779 25112 31944 25140
rect 29779 25109 29791 25112
rect 29733 25103 29791 25109
rect 31938 25100 31944 25112
rect 31996 25100 32002 25152
rect 33413 25143 33471 25149
rect 33413 25109 33425 25143
rect 33459 25140 33471 25143
rect 34054 25140 34060 25152
rect 33459 25112 34060 25140
rect 33459 25109 33471 25112
rect 33413 25103 33471 25109
rect 34054 25100 34060 25112
rect 34112 25100 34118 25152
rect 38010 25100 38016 25152
rect 38068 25100 38074 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7650 24896 7656 24948
rect 7708 24936 7714 24948
rect 7708 24908 8432 24936
rect 7708 24896 7714 24908
rect 3044 24871 3102 24877
rect 3044 24837 3056 24871
rect 3090 24868 3102 24871
rect 3970 24868 3976 24880
rect 3090 24840 3976 24868
rect 3090 24837 3102 24840
rect 3044 24831 3102 24837
rect 3970 24828 3976 24840
rect 4028 24828 4034 24880
rect 5534 24828 5540 24880
rect 5592 24828 5598 24880
rect 7009 24871 7067 24877
rect 7009 24837 7021 24871
rect 7055 24868 7067 24871
rect 7834 24868 7840 24880
rect 7055 24840 7840 24868
rect 7055 24837 7067 24840
rect 7009 24831 7067 24837
rect 7834 24828 7840 24840
rect 7892 24828 7898 24880
rect 8404 24877 8432 24908
rect 19242 24896 19248 24948
rect 19300 24896 19306 24948
rect 24302 24896 24308 24948
rect 24360 24896 24366 24948
rect 37458 24896 37464 24948
rect 37516 24896 37522 24948
rect 8389 24871 8447 24877
rect 8389 24837 8401 24871
rect 8435 24837 8447 24871
rect 8389 24831 8447 24837
rect 8478 24828 8484 24880
rect 8536 24868 8542 24880
rect 8589 24871 8647 24877
rect 8589 24868 8601 24871
rect 8536 24840 8601 24868
rect 8536 24828 8542 24840
rect 8589 24837 8601 24840
rect 8635 24837 8647 24871
rect 9766 24868 9772 24880
rect 8589 24831 8647 24837
rect 9416 24840 9772 24868
rect 2774 24760 2780 24812
rect 2832 24760 2838 24812
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24800 5135 24803
rect 5552 24800 5580 24828
rect 5123 24772 5580 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 5626 24760 5632 24812
rect 5684 24800 5690 24812
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 5684 24772 6837 24800
rect 5684 24760 5690 24772
rect 6825 24769 6837 24772
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 9416 24809 9444 24840
rect 9766 24828 9772 24840
rect 9824 24868 9830 24880
rect 9824 24840 10364 24868
rect 9824 24828 9830 24840
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 6972 24772 7113 24800
rect 6972 24760 6978 24772
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 9674 24760 9680 24812
rect 9732 24800 9738 24812
rect 10229 24803 10287 24809
rect 10229 24800 10241 24803
rect 9732 24772 10241 24800
rect 9732 24760 9738 24772
rect 10229 24769 10241 24772
rect 10275 24769 10287 24803
rect 10336 24800 10364 24840
rect 10410 24828 10416 24880
rect 10468 24828 10474 24880
rect 13446 24828 13452 24880
rect 13504 24828 13510 24880
rect 19334 24868 19340 24880
rect 18524 24840 19340 24868
rect 10336 24772 10456 24800
rect 10229 24763 10287 24769
rect 10428 24744 10456 24772
rect 10502 24760 10508 24812
rect 10560 24760 10566 24812
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 5166 24692 5172 24744
rect 5224 24692 5230 24744
rect 5261 24735 5319 24741
rect 5261 24701 5273 24735
rect 5307 24701 5319 24735
rect 5261 24695 5319 24701
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24732 5411 24735
rect 5442 24732 5448 24744
rect 5399 24704 5448 24732
rect 5399 24701 5411 24704
rect 5353 24695 5411 24701
rect 4982 24624 4988 24676
rect 5040 24664 5046 24676
rect 5276 24664 5304 24695
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 9217 24735 9275 24741
rect 5583 24704 8984 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 5040 24636 5304 24664
rect 5040 24624 5046 24636
rect 4157 24599 4215 24605
rect 4157 24565 4169 24599
rect 4203 24596 4215 24599
rect 4614 24596 4620 24608
rect 4203 24568 4620 24596
rect 4203 24565 4215 24568
rect 4157 24559 4215 24565
rect 4614 24556 4620 24568
rect 4672 24556 4678 24608
rect 5276 24596 5304 24636
rect 6730 24624 6736 24676
rect 6788 24664 6794 24676
rect 6825 24667 6883 24673
rect 6825 24664 6837 24667
rect 6788 24636 6837 24664
rect 6788 24624 6794 24636
rect 6825 24633 6837 24636
rect 6871 24633 6883 24667
rect 8956 24664 8984 24704
rect 9217 24701 9229 24735
rect 9263 24732 9275 24735
rect 9766 24732 9772 24744
rect 9263 24704 9772 24732
rect 9263 24701 9275 24704
rect 9217 24695 9275 24701
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 10410 24692 10416 24744
rect 10468 24732 10474 24744
rect 10612 24732 10640 24763
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 13265 24803 13323 24809
rect 13265 24800 13277 24803
rect 12492 24772 13277 24800
rect 12492 24760 12498 24772
rect 13265 24769 13277 24772
rect 13311 24769 13323 24803
rect 13265 24763 13323 24769
rect 13541 24803 13599 24809
rect 13541 24769 13553 24803
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 10468 24704 10640 24732
rect 10468 24692 10474 24704
rect 12710 24664 12716 24676
rect 8956 24636 12716 24664
rect 6825 24627 6883 24633
rect 12710 24624 12716 24636
rect 12768 24624 12774 24676
rect 8573 24599 8631 24605
rect 8573 24596 8585 24599
rect 5276 24568 8585 24596
rect 8573 24565 8585 24568
rect 8619 24565 8631 24599
rect 8573 24559 8631 24565
rect 8757 24599 8815 24605
rect 8757 24565 8769 24599
rect 8803 24596 8815 24599
rect 9490 24596 9496 24608
rect 8803 24568 9496 24596
rect 8803 24565 8815 24568
rect 8757 24559 8815 24565
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 9582 24556 9588 24608
rect 9640 24556 9646 24608
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 10870 24596 10876 24608
rect 10827 24568 10876 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 13556 24596 13584 24763
rect 13630 24760 13636 24812
rect 13688 24760 13694 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 13832 24772 14565 24800
rect 13832 24673 13860 24772
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 16850 24760 16856 24812
rect 16908 24760 16914 24812
rect 17678 24760 17684 24812
rect 17736 24760 17742 24812
rect 18046 24760 18052 24812
rect 18104 24760 18110 24812
rect 18524 24809 18552 24840
rect 19334 24828 19340 24840
rect 19392 24828 19398 24880
rect 20530 24868 20536 24880
rect 20180 24840 20536 24868
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 20180 24800 20208 24840
rect 20530 24828 20536 24840
rect 20588 24828 20594 24880
rect 21266 24828 21272 24880
rect 21324 24868 21330 24880
rect 22738 24868 22744 24880
rect 21324 24840 22744 24868
rect 21324 24828 21330 24840
rect 22738 24828 22744 24840
rect 22796 24828 22802 24880
rect 25041 24871 25099 24877
rect 25041 24868 25053 24871
rect 24228 24840 25053 24868
rect 19291 24772 20208 24800
rect 20257 24803 20315 24809
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 20257 24769 20269 24803
rect 20303 24800 20315 24803
rect 20438 24800 20444 24812
rect 20303 24772 20444 24800
rect 20303 24769 20315 24772
rect 20257 24763 20315 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 21910 24760 21916 24812
rect 21968 24800 21974 24812
rect 21968 24772 22094 24800
rect 21968 24760 21974 24772
rect 13906 24692 13912 24744
rect 13964 24732 13970 24744
rect 14277 24735 14335 24741
rect 14277 24732 14289 24735
rect 13964 24704 14289 24732
rect 13964 24692 13970 24704
rect 14277 24701 14289 24704
rect 14323 24732 14335 24735
rect 14458 24732 14464 24744
rect 14323 24704 14464 24732
rect 14323 24701 14335 24704
rect 14277 24695 14335 24701
rect 14458 24692 14464 24704
rect 14516 24732 14522 24744
rect 16574 24732 16580 24744
rect 14516 24704 16580 24732
rect 14516 24692 14522 24704
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 22066 24732 22094 24772
rect 23106 24760 23112 24812
rect 23164 24760 23170 24812
rect 23290 24760 23296 24812
rect 23348 24760 23354 24812
rect 23382 24760 23388 24812
rect 23440 24800 23446 24812
rect 23477 24803 23535 24809
rect 23477 24800 23489 24803
rect 23440 24772 23489 24800
rect 23440 24760 23446 24772
rect 23477 24769 23489 24772
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24800 23811 24803
rect 24228 24800 24256 24840
rect 25041 24837 25053 24840
rect 25087 24868 25099 24871
rect 25682 24868 25688 24880
rect 25087 24840 25688 24868
rect 25087 24837 25099 24840
rect 25041 24831 25099 24837
rect 25682 24828 25688 24840
rect 25740 24868 25746 24880
rect 30926 24868 30932 24880
rect 25740 24840 26234 24868
rect 25740 24828 25746 24840
rect 23799 24772 24256 24800
rect 23799 24769 23811 24772
rect 23753 24763 23811 24769
rect 24302 24760 24308 24812
rect 24360 24760 24366 24812
rect 24578 24760 24584 24812
rect 24636 24760 24642 24812
rect 24946 24760 24952 24812
rect 25004 24800 25010 24812
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 25004 24772 25237 24800
rect 25004 24760 25010 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 26206 24800 26234 24840
rect 30300 24840 30932 24868
rect 27617 24803 27675 24809
rect 27617 24800 27629 24803
rect 26206 24772 27629 24800
rect 25777 24763 25835 24769
rect 27617 24769 27629 24772
rect 27663 24800 27675 24803
rect 27706 24800 27712 24812
rect 27663 24772 27712 24800
rect 27663 24769 27675 24772
rect 27617 24763 27675 24769
rect 22925 24735 22983 24741
rect 22925 24732 22937 24735
rect 22066 24704 22937 24732
rect 22925 24701 22937 24704
rect 22971 24732 22983 24735
rect 24762 24732 24768 24744
rect 22971 24704 24768 24732
rect 22971 24701 22983 24704
rect 22925 24695 22983 24701
rect 24762 24692 24768 24704
rect 24820 24692 24826 24744
rect 25130 24692 25136 24744
rect 25188 24732 25194 24744
rect 25792 24732 25820 24763
rect 27706 24760 27712 24772
rect 27764 24760 27770 24812
rect 27890 24760 27896 24812
rect 27948 24760 27954 24812
rect 28994 24760 29000 24812
rect 29052 24760 29058 24812
rect 29454 24760 29460 24812
rect 29512 24760 29518 24812
rect 29549 24803 29607 24809
rect 29549 24769 29561 24803
rect 29595 24800 29607 24803
rect 29914 24800 29920 24812
rect 29595 24772 29920 24800
rect 29595 24769 29607 24772
rect 29549 24763 29607 24769
rect 29914 24760 29920 24772
rect 29972 24760 29978 24812
rect 30101 24803 30159 24809
rect 30101 24769 30113 24803
rect 30147 24800 30159 24803
rect 30300 24800 30328 24840
rect 30926 24828 30932 24840
rect 30984 24828 30990 24880
rect 32030 24828 32036 24880
rect 32088 24868 32094 24880
rect 37829 24871 37887 24877
rect 37829 24868 37841 24871
rect 32088 24840 37841 24868
rect 32088 24828 32094 24840
rect 37829 24837 37841 24840
rect 37875 24868 37887 24871
rect 38010 24868 38016 24880
rect 37875 24840 38016 24868
rect 37875 24837 37887 24840
rect 37829 24831 37887 24837
rect 38010 24828 38016 24840
rect 38068 24828 38074 24880
rect 30147 24772 30328 24800
rect 30147 24769 30159 24772
rect 30101 24763 30159 24769
rect 30374 24760 30380 24812
rect 30432 24760 30438 24812
rect 33686 24760 33692 24812
rect 33744 24800 33750 24812
rect 33781 24803 33839 24809
rect 33781 24800 33793 24803
rect 33744 24772 33793 24800
rect 33744 24760 33750 24772
rect 33781 24769 33793 24772
rect 33827 24769 33839 24803
rect 34957 24803 35015 24809
rect 34957 24800 34969 24803
rect 33781 24763 33839 24769
rect 34164 24772 34969 24800
rect 26142 24732 26148 24744
rect 25188 24704 26148 24732
rect 25188 24692 25194 24704
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 28077 24735 28135 24741
rect 28077 24701 28089 24735
rect 28123 24732 28135 24735
rect 28534 24732 28540 24744
rect 28123 24704 28540 24732
rect 28123 24701 28135 24704
rect 28077 24695 28135 24701
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 28810 24692 28816 24744
rect 28868 24692 28874 24744
rect 30837 24735 30895 24741
rect 30837 24701 30849 24735
rect 30883 24732 30895 24735
rect 31294 24732 31300 24744
rect 30883 24704 31300 24732
rect 30883 24701 30895 24704
rect 30837 24695 30895 24701
rect 31294 24692 31300 24704
rect 31352 24692 31358 24744
rect 33870 24692 33876 24744
rect 33928 24692 33934 24744
rect 34164 24741 34192 24772
rect 34957 24769 34969 24772
rect 35003 24769 35015 24803
rect 34957 24763 35015 24769
rect 34149 24735 34207 24741
rect 34149 24701 34161 24735
rect 34195 24701 34207 24735
rect 34149 24695 34207 24701
rect 34701 24735 34759 24741
rect 34701 24701 34713 24735
rect 34747 24701 34759 24735
rect 34701 24695 34759 24701
rect 13817 24667 13875 24673
rect 13817 24633 13829 24667
rect 13863 24633 13875 24667
rect 13817 24627 13875 24633
rect 15841 24667 15899 24673
rect 15841 24633 15853 24667
rect 15887 24664 15899 24667
rect 26234 24664 26240 24676
rect 15887 24636 26240 24664
rect 15887 24633 15899 24636
rect 15841 24627 15899 24633
rect 15856 24596 15884 24627
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 26476 24636 28396 24664
rect 26476 24624 26482 24636
rect 13556 24568 15884 24596
rect 18414 24556 18420 24608
rect 18472 24556 18478 24608
rect 27614 24556 27620 24608
rect 27672 24596 27678 24608
rect 27709 24599 27767 24605
rect 27709 24596 27721 24599
rect 27672 24568 27721 24596
rect 27672 24556 27678 24568
rect 27709 24565 27721 24568
rect 27755 24565 27767 24599
rect 28368 24596 28396 24636
rect 28626 24624 28632 24676
rect 28684 24664 28690 24676
rect 29546 24664 29552 24676
rect 28684 24636 29552 24664
rect 28684 24624 28690 24636
rect 29546 24624 29552 24636
rect 29604 24624 29610 24676
rect 29914 24624 29920 24676
rect 29972 24664 29978 24676
rect 30193 24667 30251 24673
rect 30193 24664 30205 24667
rect 29972 24636 30205 24664
rect 29972 24624 29978 24636
rect 30193 24633 30205 24636
rect 30239 24633 30251 24667
rect 30193 24627 30251 24633
rect 32674 24624 32680 24676
rect 32732 24664 32738 24676
rect 34716 24664 34744 24695
rect 37918 24692 37924 24744
rect 37976 24692 37982 24744
rect 38102 24692 38108 24744
rect 38160 24692 38166 24744
rect 32732 24636 34744 24664
rect 32732 24624 32738 24636
rect 30006 24596 30012 24608
rect 28368 24568 30012 24596
rect 27709 24559 27767 24565
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 35986 24556 35992 24608
rect 36044 24596 36050 24608
rect 36081 24599 36139 24605
rect 36081 24596 36093 24599
rect 36044 24568 36093 24596
rect 36044 24556 36050 24568
rect 36081 24565 36093 24568
rect 36127 24565 36139 24599
rect 36081 24559 36139 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 5166 24352 5172 24404
rect 5224 24392 5230 24404
rect 5994 24392 6000 24404
rect 5224 24364 6000 24392
rect 5224 24352 5230 24364
rect 5994 24352 6000 24364
rect 6052 24352 6058 24404
rect 10502 24352 10508 24404
rect 10560 24392 10566 24404
rect 11977 24395 12035 24401
rect 11977 24392 11989 24395
rect 10560 24364 11989 24392
rect 10560 24352 10566 24364
rect 11977 24361 11989 24364
rect 12023 24361 12035 24395
rect 11977 24355 12035 24361
rect 5718 24284 5724 24336
rect 5776 24324 5782 24336
rect 11992 24324 12020 24355
rect 12066 24352 12072 24404
rect 12124 24392 12130 24404
rect 16850 24392 16856 24404
rect 12124 24364 16856 24392
rect 12124 24352 12130 24364
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 23198 24352 23204 24404
rect 23256 24352 23262 24404
rect 24118 24392 24124 24404
rect 23308 24364 24124 24392
rect 18690 24324 18696 24336
rect 5776 24296 7144 24324
rect 11992 24296 18696 24324
rect 5776 24284 5782 24296
rect 5350 24216 5356 24268
rect 5408 24256 5414 24268
rect 5626 24256 5632 24268
rect 5408 24228 5632 24256
rect 5408 24216 5414 24228
rect 5626 24216 5632 24228
rect 5684 24256 5690 24268
rect 7116 24256 7144 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 8018 24256 8024 24268
rect 5684 24228 6040 24256
rect 5684 24216 5690 24228
rect 5718 24148 5724 24200
rect 5776 24148 5782 24200
rect 5810 24148 5816 24200
rect 5868 24148 5874 24200
rect 6012 24197 6040 24228
rect 7116 24228 8024 24256
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 6546 24148 6552 24200
rect 6604 24188 6610 24200
rect 7116 24197 7144 24228
rect 8018 24216 8024 24228
rect 8076 24256 8082 24268
rect 9309 24259 9367 24265
rect 9309 24256 9321 24259
rect 8076 24228 9321 24256
rect 8076 24216 8082 24228
rect 9309 24225 9321 24228
rect 9355 24225 9367 24259
rect 9309 24219 9367 24225
rect 9398 24216 9404 24268
rect 9456 24216 9462 24268
rect 9582 24216 9588 24268
rect 9640 24216 9646 24268
rect 16850 24216 16856 24268
rect 16908 24256 16914 24268
rect 16908 24228 19748 24256
rect 16908 24216 16914 24228
rect 6825 24191 6883 24197
rect 6825 24188 6837 24191
rect 6604 24160 6837 24188
rect 6604 24148 6610 24160
rect 6825 24157 6837 24160
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 7101 24191 7159 24197
rect 7101 24157 7113 24191
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 8110 24188 8116 24200
rect 7699 24160 8116 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 10318 24188 10324 24200
rect 9539 24160 10324 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 12342 24188 12348 24200
rect 10643 24160 12348 24188
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24188 17279 24191
rect 17310 24188 17316 24200
rect 17267 24160 17316 24188
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17402 24148 17408 24200
rect 17460 24148 17466 24200
rect 17770 24148 17776 24200
rect 17828 24148 17834 24200
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18230 24148 18236 24200
rect 18288 24148 18294 24200
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 18840 24160 19625 24188
rect 18840 24148 18846 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19720 24188 19748 24228
rect 20806 24216 20812 24268
rect 20864 24256 20870 24268
rect 20864 24228 22048 24256
rect 20864 24216 20870 24228
rect 21450 24188 21456 24200
rect 19720 24160 21456 24188
rect 19613 24151 19671 24157
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22020 24197 22048 24228
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 22704 24228 23152 24256
rect 22704 24216 22710 24228
rect 21821 24191 21879 24197
rect 21821 24188 21833 24191
rect 21784 24160 21833 24188
rect 21784 24148 21790 24160
rect 21821 24157 21833 24160
rect 21867 24157 21879 24191
rect 21821 24151 21879 24157
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 10870 24129 10876 24132
rect 10864 24120 10876 24129
rect 4672 24092 9260 24120
rect 10831 24092 10876 24120
rect 4672 24080 4678 24092
rect 6178 24012 6184 24064
rect 6236 24012 6242 24064
rect 6638 24012 6644 24064
rect 6696 24012 6702 24064
rect 7006 24012 7012 24064
rect 7064 24052 7070 24064
rect 7650 24052 7656 24064
rect 7064 24024 7656 24052
rect 7064 24012 7070 24024
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24052 7803 24055
rect 7834 24052 7840 24064
rect 7791 24024 7840 24052
rect 7791 24021 7803 24024
rect 7745 24015 7803 24021
rect 7834 24012 7840 24024
rect 7892 24012 7898 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 9232 24052 9260 24092
rect 10864 24083 10876 24092
rect 10870 24080 10876 24083
rect 10928 24080 10934 24132
rect 15286 24080 15292 24132
rect 15344 24120 15350 24132
rect 18248 24120 18276 24148
rect 15344 24092 18276 24120
rect 18693 24123 18751 24129
rect 15344 24080 15350 24092
rect 18693 24089 18705 24123
rect 18739 24120 18751 24123
rect 19334 24120 19340 24132
rect 18739 24092 19340 24120
rect 18739 24089 18751 24092
rect 18693 24083 18751 24089
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 19705 24123 19763 24129
rect 19705 24089 19717 24123
rect 19751 24120 19763 24123
rect 20717 24123 20775 24129
rect 20717 24120 20729 24123
rect 19751 24092 20729 24120
rect 19751 24089 19763 24092
rect 19705 24083 19763 24089
rect 20717 24089 20729 24092
rect 20763 24089 20775 24123
rect 22020 24120 22048 24151
rect 23014 24148 23020 24200
rect 23072 24148 23078 24200
rect 23124 24188 23152 24228
rect 23198 24216 23204 24268
rect 23256 24256 23262 24268
rect 23308 24265 23336 24364
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 24302 24352 24308 24404
rect 24360 24392 24366 24404
rect 24360 24364 27108 24392
rect 24360 24352 24366 24364
rect 25222 24324 25228 24336
rect 24044 24296 25228 24324
rect 23293 24259 23351 24265
rect 23293 24256 23305 24259
rect 23256 24228 23305 24256
rect 23256 24216 23262 24228
rect 23293 24225 23305 24228
rect 23339 24225 23351 24259
rect 23293 24219 23351 24225
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 24044 24256 24072 24296
rect 25222 24284 25228 24296
rect 25280 24284 25286 24336
rect 26142 24284 26148 24336
rect 26200 24324 26206 24336
rect 27080 24333 27108 24364
rect 27614 24352 27620 24404
rect 27672 24392 27678 24404
rect 30374 24392 30380 24404
rect 27672 24364 30380 24392
rect 27672 24352 27678 24364
rect 27065 24327 27123 24333
rect 26200 24296 27016 24324
rect 26200 24284 26206 24296
rect 23440 24228 24072 24256
rect 23440 24216 23446 24228
rect 23124 24160 23428 24188
rect 23400 24132 23428 24160
rect 23842 24148 23848 24200
rect 23900 24148 23906 24200
rect 24044 24197 24072 24228
rect 24394 24216 24400 24268
rect 24452 24256 24458 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24452 24228 24593 24256
rect 24452 24216 24458 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 25774 24216 25780 24268
rect 25832 24256 25838 24268
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 25832 24228 26341 24256
rect 25832 24216 25838 24228
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26329 24219 26387 24225
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24157 24087 24191
rect 24029 24151 24087 24157
rect 24670 24148 24676 24200
rect 24728 24188 24734 24200
rect 24857 24191 24915 24197
rect 24857 24188 24869 24191
rect 24728 24160 24869 24188
rect 24728 24148 24734 24160
rect 24857 24157 24869 24160
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24188 26847 24191
rect 26878 24188 26884 24200
rect 26835 24160 26884 24188
rect 26835 24157 26847 24160
rect 26789 24151 26847 24157
rect 26878 24148 26884 24160
rect 26936 24148 26942 24200
rect 26988 24188 27016 24296
rect 27065 24293 27077 24327
rect 27111 24324 27123 24327
rect 29362 24324 29368 24336
rect 27111 24296 29368 24324
rect 27111 24293 27123 24296
rect 27065 24287 27123 24293
rect 29362 24284 29368 24296
rect 29420 24284 29426 24336
rect 28718 24256 28724 24268
rect 28431 24228 28724 24256
rect 27249 24191 27307 24197
rect 27249 24188 27261 24191
rect 26988 24160 27261 24188
rect 27249 24157 27261 24160
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 27890 24148 27896 24200
rect 27948 24188 27954 24200
rect 28431 24197 28459 24228
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 28031 24191 28089 24197
rect 28031 24188 28043 24191
rect 27948 24160 28043 24188
rect 27948 24148 27954 24160
rect 28031 24157 28043 24160
rect 28077 24157 28089 24191
rect 28431 24191 28502 24197
rect 28431 24160 28456 24191
rect 28031 24151 28089 24157
rect 28444 24157 28456 24160
rect 28490 24157 28502 24191
rect 28444 24151 28502 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24188 28595 24191
rect 28626 24188 28632 24200
rect 28583 24160 28632 24188
rect 28583 24157 28595 24160
rect 28537 24151 28595 24157
rect 28626 24148 28632 24160
rect 28684 24148 28690 24200
rect 29546 24148 29552 24200
rect 29604 24188 29610 24200
rect 29825 24191 29883 24197
rect 29825 24188 29837 24191
rect 29604 24160 29837 24188
rect 29604 24148 29610 24160
rect 29825 24157 29837 24160
rect 29871 24157 29883 24191
rect 29825 24151 29883 24157
rect 29914 24148 29920 24200
rect 29972 24148 29978 24200
rect 30116 24197 30144 24364
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 33778 24392 33784 24404
rect 31726 24364 33784 24392
rect 31726 24324 31754 24364
rect 33778 24352 33784 24364
rect 33836 24352 33842 24404
rect 34149 24395 34207 24401
rect 34149 24361 34161 24395
rect 34195 24392 34207 24395
rect 34238 24392 34244 24404
rect 34195 24364 34244 24392
rect 34195 24361 34207 24364
rect 34149 24355 34207 24361
rect 34238 24352 34244 24364
rect 34296 24352 34302 24404
rect 34698 24352 34704 24404
rect 34756 24392 34762 24404
rect 34885 24395 34943 24401
rect 34885 24392 34897 24395
rect 34756 24364 34897 24392
rect 34756 24352 34762 24364
rect 34885 24361 34897 24364
rect 34931 24361 34943 24395
rect 34885 24355 34943 24361
rect 30576 24296 31754 24324
rect 30576 24265 30604 24296
rect 31846 24284 31852 24336
rect 31904 24324 31910 24336
rect 31904 24296 32536 24324
rect 31904 24284 31910 24296
rect 30561 24259 30619 24265
rect 30561 24225 30573 24259
rect 30607 24225 30619 24259
rect 31478 24256 31484 24268
rect 30561 24219 30619 24225
rect 31368 24228 31484 24256
rect 30101 24191 30159 24197
rect 30101 24157 30113 24191
rect 30147 24157 30159 24191
rect 30101 24151 30159 24157
rect 31202 24148 31208 24200
rect 31260 24148 31266 24200
rect 31368 24197 31396 24228
rect 31478 24216 31484 24228
rect 31536 24216 31542 24268
rect 32030 24256 32036 24268
rect 31588 24228 32036 24256
rect 31588 24197 31616 24228
rect 32030 24216 32036 24228
rect 32088 24216 32094 24268
rect 32398 24216 32404 24268
rect 32456 24216 32462 24268
rect 31353 24191 31411 24197
rect 31353 24157 31365 24191
rect 31399 24157 31411 24191
rect 31353 24151 31411 24157
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24157 31631 24191
rect 31573 24151 31631 24157
rect 31670 24191 31728 24197
rect 31670 24157 31682 24191
rect 31716 24157 31728 24191
rect 31670 24151 31728 24157
rect 22020 24092 23336 24120
rect 20717 24083 20775 24089
rect 23308 24064 23336 24092
rect 23382 24080 23388 24132
rect 23440 24080 23446 24132
rect 24949 24123 25007 24129
rect 24949 24120 24961 24123
rect 24688 24092 24961 24120
rect 12066 24052 12072 24064
rect 9232 24024 12072 24052
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 20254 24012 20260 24064
rect 20312 24012 20318 24064
rect 20625 24055 20683 24061
rect 20625 24021 20637 24055
rect 20671 24052 20683 24055
rect 21082 24052 21088 24064
rect 20671 24024 21088 24052
rect 20671 24021 20683 24024
rect 20625 24015 20683 24021
rect 21082 24012 21088 24024
rect 21140 24012 21146 24064
rect 22830 24012 22836 24064
rect 22888 24012 22894 24064
rect 23290 24012 23296 24064
rect 23348 24012 23354 24064
rect 23937 24055 23995 24061
rect 23937 24021 23949 24055
rect 23983 24052 23995 24055
rect 24688 24052 24716 24092
rect 24949 24089 24961 24092
rect 24995 24089 25007 24123
rect 24949 24083 25007 24089
rect 25317 24123 25375 24129
rect 25317 24089 25329 24123
rect 25363 24120 25375 24123
rect 27154 24120 27160 24132
rect 25363 24092 27160 24120
rect 25363 24089 25375 24092
rect 25317 24083 25375 24089
rect 27154 24080 27160 24092
rect 27212 24080 27218 24132
rect 27706 24080 27712 24132
rect 27764 24120 27770 24132
rect 27764 24092 28120 24120
rect 27764 24080 27770 24092
rect 23983 24024 24716 24052
rect 23983 24021 23995 24024
rect 23937 24015 23995 24021
rect 24762 24012 24768 24064
rect 24820 24012 24826 24064
rect 27893 24055 27951 24061
rect 27893 24021 27905 24055
rect 27939 24052 27951 24055
rect 27982 24052 27988 24064
rect 27939 24024 27988 24052
rect 27939 24021 27951 24024
rect 27893 24015 27951 24021
rect 27982 24012 27988 24024
rect 28040 24012 28046 24064
rect 28092 24052 28120 24092
rect 28166 24080 28172 24132
rect 28224 24080 28230 24132
rect 28261 24123 28319 24129
rect 28261 24089 28273 24123
rect 28307 24120 28319 24123
rect 28810 24120 28816 24132
rect 28307 24092 28816 24120
rect 28307 24089 28319 24092
rect 28261 24083 28319 24089
rect 28810 24080 28816 24092
rect 28868 24080 28874 24132
rect 29730 24120 29736 24132
rect 29196 24092 29736 24120
rect 29196 24052 29224 24092
rect 29730 24080 29736 24092
rect 29788 24080 29794 24132
rect 30006 24080 30012 24132
rect 30064 24120 30070 24132
rect 31481 24123 31539 24129
rect 31481 24120 31493 24123
rect 30064 24092 31493 24120
rect 30064 24080 30070 24092
rect 31481 24089 31493 24092
rect 31527 24089 31539 24123
rect 31481 24083 31539 24089
rect 28092 24024 29224 24052
rect 29270 24012 29276 24064
rect 29328 24052 29334 24064
rect 30834 24052 30840 24064
rect 29328 24024 30840 24052
rect 29328 24012 29334 24024
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 31294 24012 31300 24064
rect 31352 24052 31358 24064
rect 31685 24052 31713 24151
rect 32306 24148 32312 24200
rect 32364 24148 32370 24200
rect 32508 24188 32536 24296
rect 33686 24216 33692 24268
rect 33744 24256 33750 24268
rect 34256 24256 34284 24352
rect 35253 24259 35311 24265
rect 35253 24256 35265 24259
rect 33744 24228 34008 24256
rect 34256 24228 35265 24256
rect 33744 24216 33750 24228
rect 32585 24191 32643 24197
rect 32585 24188 32597 24191
rect 32508 24160 32597 24188
rect 32585 24157 32597 24160
rect 32631 24157 32643 24191
rect 32585 24151 32643 24157
rect 32677 24191 32735 24197
rect 32677 24157 32689 24191
rect 32723 24157 32735 24191
rect 32677 24151 32735 24157
rect 33781 24191 33839 24197
rect 33781 24157 33793 24191
rect 33827 24188 33839 24191
rect 33870 24188 33876 24200
rect 33827 24160 33876 24188
rect 33827 24157 33839 24160
rect 33781 24151 33839 24157
rect 32692 24120 32720 24151
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 33980 24197 34008 24228
rect 35253 24225 35265 24228
rect 35299 24225 35311 24259
rect 35253 24219 35311 24225
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 34054 24148 34060 24200
rect 34112 24188 34118 24200
rect 35069 24191 35127 24197
rect 35069 24188 35081 24191
rect 34112 24160 35081 24188
rect 34112 24148 34118 24160
rect 35069 24157 35081 24160
rect 35115 24157 35127 24191
rect 35069 24151 35127 24157
rect 37826 24148 37832 24200
rect 37884 24148 37890 24200
rect 31864 24092 32720 24120
rect 38105 24123 38163 24129
rect 31864 24061 31892 24092
rect 38105 24089 38117 24123
rect 38151 24120 38163 24123
rect 39022 24120 39028 24132
rect 38151 24092 39028 24120
rect 38151 24089 38163 24092
rect 38105 24083 38163 24089
rect 39022 24080 39028 24092
rect 39080 24080 39086 24132
rect 31352 24024 31713 24052
rect 31849 24055 31907 24061
rect 31352 24012 31358 24024
rect 31849 24021 31861 24055
rect 31895 24021 31907 24055
rect 31849 24015 31907 24021
rect 32030 24012 32036 24064
rect 32088 24052 32094 24064
rect 32490 24052 32496 24064
rect 32088 24024 32496 24052
rect 32088 24012 32094 24024
rect 32490 24012 32496 24024
rect 32548 24012 32554 24064
rect 32861 24055 32919 24061
rect 32861 24021 32873 24055
rect 32907 24052 32919 24055
rect 37918 24052 37924 24064
rect 32907 24024 37924 24052
rect 32907 24021 32919 24024
rect 32861 24015 32919 24021
rect 37918 24012 37924 24024
rect 37976 24012 37982 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 4157 23851 4215 23857
rect 4157 23817 4169 23851
rect 4203 23848 4215 23851
rect 4890 23848 4896 23860
rect 4203 23820 4896 23848
rect 4203 23817 4215 23820
rect 4157 23811 4215 23817
rect 4890 23808 4896 23820
rect 4948 23848 4954 23860
rect 17954 23848 17960 23860
rect 4948 23820 17960 23848
rect 4948 23808 4954 23820
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 21450 23808 21456 23860
rect 21508 23848 21514 23860
rect 29914 23848 29920 23860
rect 21508 23820 29920 23848
rect 21508 23808 21514 23820
rect 29914 23808 29920 23820
rect 29972 23808 29978 23860
rect 32858 23808 32864 23860
rect 32916 23808 32922 23860
rect 33321 23851 33379 23857
rect 33321 23817 33333 23851
rect 33367 23848 33379 23851
rect 33367 23820 33824 23848
rect 33367 23817 33379 23820
rect 33321 23811 33379 23817
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 5534 23780 5540 23792
rect 4120 23752 4936 23780
rect 4120 23740 4126 23752
rect 2774 23672 2780 23724
rect 2832 23672 2838 23724
rect 3044 23715 3102 23721
rect 3044 23681 3056 23715
rect 3090 23712 3102 23715
rect 3970 23712 3976 23724
rect 3090 23684 3976 23712
rect 3090 23681 3102 23684
rect 3044 23675 3102 23681
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 4908 23721 4936 23752
rect 5092 23752 5540 23780
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23712 4951 23715
rect 4982 23712 4988 23724
rect 4939 23684 4988 23712
rect 4939 23681 4951 23684
rect 4893 23675 4951 23681
rect 4982 23672 4988 23684
rect 5040 23672 5046 23724
rect 5092 23721 5120 23752
rect 5534 23740 5540 23752
rect 5592 23740 5598 23792
rect 5902 23780 5908 23792
rect 5644 23752 5908 23780
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23681 5135 23715
rect 5077 23675 5135 23681
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5644 23721 5672 23752
rect 5902 23740 5908 23752
rect 5960 23740 5966 23792
rect 5994 23740 6000 23792
rect 6052 23780 6058 23792
rect 7006 23780 7012 23792
rect 6052 23752 7012 23780
rect 6052 23740 6058 23752
rect 7006 23740 7012 23752
rect 7064 23740 7070 23792
rect 7834 23740 7840 23792
rect 7892 23780 7898 23792
rect 8656 23783 8714 23789
rect 7892 23752 8524 23780
rect 7892 23740 7898 23752
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 6012 23712 6040 23740
rect 5859 23684 6040 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6730 23672 6736 23724
rect 6788 23672 6794 23724
rect 8386 23672 8392 23724
rect 8444 23672 8450 23724
rect 8496 23712 8524 23752
rect 8656 23749 8668 23783
rect 8702 23780 8714 23783
rect 9122 23780 9128 23792
rect 8702 23752 9128 23780
rect 8702 23749 8714 23752
rect 8656 23743 8714 23749
rect 9122 23740 9128 23752
rect 9180 23740 9186 23792
rect 12342 23740 12348 23792
rect 12400 23780 12406 23792
rect 13906 23780 13912 23792
rect 12400 23752 13912 23780
rect 12400 23740 12406 23752
rect 12728 23721 12756 23752
rect 13906 23740 13912 23752
rect 13964 23740 13970 23792
rect 18230 23740 18236 23792
rect 18288 23780 18294 23792
rect 21266 23780 21272 23792
rect 18288 23752 21272 23780
rect 18288 23740 18294 23752
rect 12713 23715 12771 23721
rect 8496 23684 12434 23712
rect 4816 23644 4844 23672
rect 5721 23647 5779 23653
rect 5721 23644 5733 23647
rect 4816 23616 5733 23644
rect 5721 23613 5733 23616
rect 5767 23613 5779 23647
rect 12406 23644 12434 23684
rect 12713 23681 12725 23715
rect 12759 23681 12771 23715
rect 12969 23715 13027 23721
rect 12969 23712 12981 23715
rect 12713 23675 12771 23681
rect 12820 23684 12981 23712
rect 12820 23644 12848 23684
rect 12969 23681 12981 23684
rect 13015 23681 13027 23715
rect 12969 23675 13027 23681
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 17218 23712 17224 23724
rect 17083 23684 17224 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 20456 23721 20484 23752
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 22186 23740 22192 23792
rect 22244 23780 22250 23792
rect 22244 23752 25636 23780
rect 22244 23740 22250 23752
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 19484 23684 20269 23712
rect 19484 23672 19490 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20257 23675 20315 23681
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23681 20499 23715
rect 20441 23675 20499 23681
rect 20533 23715 20591 23721
rect 20533 23681 20545 23715
rect 20579 23712 20591 23715
rect 20806 23712 20812 23724
rect 20579 23684 20812 23712
rect 20579 23681 20591 23684
rect 20533 23675 20591 23681
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 23106 23672 23112 23724
rect 23164 23712 23170 23724
rect 23201 23715 23259 23721
rect 23201 23712 23213 23715
rect 23164 23684 23213 23712
rect 23164 23672 23170 23684
rect 23201 23681 23213 23684
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 23382 23672 23388 23724
rect 23440 23672 23446 23724
rect 24213 23715 24271 23721
rect 24213 23681 24225 23715
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 12406 23616 12848 23644
rect 5721 23607 5779 23613
rect 17126 23604 17132 23656
rect 17184 23644 17190 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 17184 23616 17417 23644
rect 17184 23604 17190 23616
rect 17405 23613 17417 23616
rect 17451 23644 17463 23647
rect 21634 23644 21640 23656
rect 17451 23616 21640 23644
rect 17451 23613 17463 23616
rect 17405 23607 17463 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 24228 23644 24256 23675
rect 24762 23672 24768 23724
rect 24820 23672 24826 23724
rect 25608 23721 25636 23752
rect 26234 23740 26240 23792
rect 26292 23780 26298 23792
rect 27801 23783 27859 23789
rect 27801 23780 27813 23783
rect 26292 23752 27813 23780
rect 26292 23740 26298 23752
rect 27801 23749 27813 23752
rect 27847 23749 27859 23783
rect 27801 23743 27859 23749
rect 27982 23740 27988 23792
rect 28040 23740 28046 23792
rect 30193 23783 30251 23789
rect 29472 23752 30144 23780
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23681 25651 23715
rect 25593 23675 25651 23681
rect 27706 23672 27712 23724
rect 27764 23672 27770 23724
rect 28626 23672 28632 23724
rect 28684 23672 28690 23724
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23681 28871 23715
rect 28813 23675 28871 23681
rect 28997 23715 29055 23721
rect 28997 23681 29009 23715
rect 29043 23712 29055 23715
rect 29270 23712 29276 23724
rect 29043 23684 29276 23712
rect 29043 23681 29055 23684
rect 28997 23675 29055 23681
rect 24578 23644 24584 23656
rect 24228 23616 24584 23644
rect 24578 23604 24584 23616
rect 24636 23644 24642 23656
rect 25777 23647 25835 23653
rect 24636 23616 25084 23644
rect 24636 23604 24642 23616
rect 16298 23576 16304 23588
rect 14016 23548 16304 23576
rect 4614 23468 4620 23520
rect 4672 23468 4678 23520
rect 6825 23511 6883 23517
rect 6825 23477 6837 23511
rect 6871 23508 6883 23511
rect 8570 23508 8576 23520
rect 6871 23480 8576 23508
rect 6871 23477 6883 23480
rect 6825 23471 6883 23477
rect 8570 23468 8576 23480
rect 8628 23468 8634 23520
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 14016 23508 14044 23548
rect 16298 23536 16304 23548
rect 16356 23536 16362 23588
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 20622 23576 20628 23588
rect 20404 23548 20628 23576
rect 20404 23536 20410 23548
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 23474 23536 23480 23588
rect 23532 23536 23538 23588
rect 9824 23480 14044 23508
rect 14093 23511 14151 23517
rect 9824 23468 9830 23480
rect 14093 23477 14105 23511
rect 14139 23508 14151 23511
rect 16942 23508 16948 23520
rect 14139 23480 16948 23508
rect 14139 23477 14151 23480
rect 14093 23471 14151 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 20714 23468 20720 23520
rect 20772 23468 20778 23520
rect 25056 23517 25084 23616
rect 25777 23613 25789 23647
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 26053 23647 26111 23653
rect 26053 23613 26065 23647
rect 26099 23613 26111 23647
rect 26053 23607 26111 23613
rect 25130 23536 25136 23588
rect 25188 23576 25194 23588
rect 25792 23576 25820 23607
rect 25188 23548 25820 23576
rect 26068 23576 26096 23607
rect 26142 23604 26148 23656
rect 26200 23604 26206 23656
rect 27338 23604 27344 23656
rect 27396 23644 27402 23656
rect 28736 23644 28764 23675
rect 27396 23616 28764 23644
rect 28828 23644 28856 23675
rect 29270 23672 29276 23684
rect 29328 23672 29334 23724
rect 29362 23672 29368 23724
rect 29420 23712 29426 23724
rect 29472 23721 29500 23752
rect 29457 23715 29515 23721
rect 29457 23712 29469 23715
rect 29420 23684 29469 23712
rect 29420 23672 29426 23684
rect 29457 23681 29469 23684
rect 29503 23681 29515 23715
rect 29457 23675 29515 23681
rect 29730 23672 29736 23724
rect 29788 23672 29794 23724
rect 30116 23712 30144 23752
rect 30193 23749 30205 23783
rect 30239 23780 30251 23783
rect 30650 23780 30656 23792
rect 30239 23752 30656 23780
rect 30239 23749 30251 23752
rect 30193 23743 30251 23749
rect 30650 23740 30656 23752
rect 30708 23740 30714 23792
rect 32214 23740 32220 23792
rect 32272 23780 32278 23792
rect 32876 23780 32904 23808
rect 33796 23789 33824 23820
rect 33870 23808 33876 23860
rect 33928 23857 33934 23860
rect 33928 23848 33937 23857
rect 35529 23851 35587 23857
rect 33928 23820 33973 23848
rect 34164 23820 35480 23848
rect 33928 23811 33937 23820
rect 33928 23808 33934 23811
rect 34164 23792 34192 23820
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 32272 23752 32965 23780
rect 32272 23740 32278 23752
rect 32953 23749 32965 23752
rect 32999 23749 33011 23783
rect 32953 23743 33011 23749
rect 33781 23783 33839 23789
rect 33781 23749 33793 23783
rect 33827 23749 33839 23783
rect 33781 23743 33839 23749
rect 33965 23783 34023 23789
rect 33965 23749 33977 23783
rect 34011 23780 34023 23783
rect 34146 23780 34152 23792
rect 34011 23752 34152 23780
rect 34011 23749 34023 23752
rect 33965 23743 34023 23749
rect 34146 23740 34152 23752
rect 34204 23740 34210 23792
rect 34606 23740 34612 23792
rect 34664 23780 34670 23792
rect 35161 23783 35219 23789
rect 35161 23780 35173 23783
rect 34664 23752 35173 23780
rect 34664 23740 34670 23752
rect 35161 23749 35173 23752
rect 35207 23749 35219 23783
rect 35161 23743 35219 23749
rect 30558 23712 30564 23724
rect 30116 23684 30564 23712
rect 30558 23672 30564 23684
rect 30616 23672 30622 23724
rect 31018 23672 31024 23724
rect 31076 23672 31082 23724
rect 31570 23672 31576 23724
rect 31628 23672 31634 23724
rect 31754 23672 31760 23724
rect 31812 23712 31818 23724
rect 32677 23715 32735 23721
rect 32677 23712 32689 23715
rect 31812 23684 32689 23712
rect 31812 23672 31818 23684
rect 32677 23681 32689 23684
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32825 23715 32883 23721
rect 32825 23681 32837 23715
rect 32871 23681 32883 23715
rect 32825 23675 32883 23681
rect 28902 23644 28908 23656
rect 28828 23616 28908 23644
rect 27396 23604 27402 23616
rect 27890 23576 27896 23588
rect 26068 23548 27896 23576
rect 25188 23536 25194 23548
rect 27890 23536 27896 23548
rect 27948 23536 27954 23588
rect 27985 23579 28043 23585
rect 27985 23545 27997 23579
rect 28031 23576 28043 23579
rect 28074 23576 28080 23588
rect 28031 23548 28080 23576
rect 28031 23545 28043 23548
rect 27985 23539 28043 23545
rect 28074 23536 28080 23548
rect 28132 23536 28138 23588
rect 28736 23576 28764 23616
rect 28902 23604 28908 23616
rect 28960 23644 28966 23656
rect 29546 23644 29552 23656
rect 28960 23616 29552 23644
rect 28960 23604 28966 23616
rect 29546 23604 29552 23616
rect 29604 23604 29610 23656
rect 30837 23647 30895 23653
rect 30837 23613 30849 23647
rect 30883 23644 30895 23647
rect 31110 23644 31116 23656
rect 30883 23616 31116 23644
rect 30883 23613 30895 23616
rect 30837 23607 30895 23613
rect 31110 23604 31116 23616
rect 31168 23604 31174 23656
rect 32306 23644 32312 23656
rect 31496 23616 32312 23644
rect 31496 23576 31524 23616
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 28736 23548 31524 23576
rect 31573 23579 31631 23585
rect 31573 23545 31585 23579
rect 31619 23576 31631 23579
rect 32840 23576 32868 23675
rect 33042 23672 33048 23724
rect 33100 23672 33106 23724
rect 33183 23715 33241 23721
rect 33183 23681 33195 23715
rect 33229 23712 33241 23715
rect 33502 23712 33508 23724
rect 33229 23684 33508 23712
rect 33229 23681 33241 23684
rect 33183 23675 33241 23681
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 33594 23672 33600 23724
rect 33652 23712 33658 23724
rect 34057 23715 34115 23721
rect 34057 23712 34069 23715
rect 33652 23684 34069 23712
rect 33652 23672 33658 23684
rect 34057 23681 34069 23684
rect 34103 23681 34115 23715
rect 34057 23675 34115 23681
rect 34514 23672 34520 23724
rect 34572 23712 34578 23724
rect 34790 23712 34796 23724
rect 34572 23684 34796 23712
rect 34572 23672 34578 23684
rect 34790 23672 34796 23684
rect 34848 23712 34854 23724
rect 34885 23715 34943 23721
rect 34885 23712 34897 23715
rect 34848 23684 34897 23712
rect 34848 23672 34854 23684
rect 34885 23681 34897 23684
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 34978 23715 35036 23721
rect 34978 23681 34990 23715
rect 35024 23681 35036 23715
rect 34978 23675 35036 23681
rect 35253 23715 35311 23721
rect 35253 23681 35265 23715
rect 35299 23681 35311 23715
rect 35253 23675 35311 23681
rect 34698 23604 34704 23656
rect 34756 23644 34762 23656
rect 34992 23644 35020 23675
rect 34756 23616 35020 23644
rect 35268 23644 35296 23675
rect 35342 23672 35348 23724
rect 35400 23721 35406 23724
rect 35400 23675 35408 23721
rect 35452 23712 35480 23820
rect 35529 23817 35541 23851
rect 35575 23817 35587 23851
rect 35529 23811 35587 23817
rect 35544 23780 35572 23811
rect 37826 23808 37832 23860
rect 37884 23808 37890 23860
rect 36541 23783 36599 23789
rect 35544 23752 36400 23780
rect 35986 23712 35992 23724
rect 35452 23684 35992 23712
rect 35400 23672 35406 23675
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 36372 23721 36400 23752
rect 36541 23749 36553 23783
rect 36587 23780 36599 23783
rect 37844 23780 37872 23808
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 36587 23752 37933 23780
rect 36587 23749 36599 23752
rect 36541 23743 36599 23749
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 36357 23715 36415 23721
rect 36357 23681 36369 23715
rect 36403 23681 36415 23715
rect 37829 23715 37887 23721
rect 37829 23712 37841 23715
rect 36357 23675 36415 23681
rect 36464 23684 37841 23712
rect 36464 23644 36492 23684
rect 37829 23681 37841 23684
rect 37875 23712 37887 23715
rect 38194 23712 38200 23724
rect 37875 23684 38200 23712
rect 37875 23681 37887 23684
rect 37829 23675 37887 23681
rect 38194 23672 38200 23684
rect 38252 23672 38258 23724
rect 35268 23616 36492 23644
rect 34756 23604 34762 23616
rect 35268 23576 35296 23616
rect 38102 23604 38108 23656
rect 38160 23604 38166 23656
rect 31619 23548 31754 23576
rect 32840 23548 35296 23576
rect 31619 23545 31631 23548
rect 31573 23539 31631 23545
rect 25041 23511 25099 23517
rect 25041 23477 25053 23511
rect 25087 23508 25099 23511
rect 25498 23508 25504 23520
rect 25087 23480 25504 23508
rect 25087 23477 25099 23480
rect 25041 23471 25099 23477
rect 25498 23468 25504 23480
rect 25556 23468 25562 23520
rect 28442 23468 28448 23520
rect 28500 23468 28506 23520
rect 28534 23468 28540 23520
rect 28592 23508 28598 23520
rect 28902 23508 28908 23520
rect 28592 23480 28908 23508
rect 28592 23468 28598 23480
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 29362 23468 29368 23520
rect 29420 23508 29426 23520
rect 31478 23508 31484 23520
rect 29420 23480 31484 23508
rect 29420 23468 29426 23480
rect 31478 23468 31484 23480
rect 31536 23468 31542 23520
rect 31726 23508 31754 23548
rect 35802 23536 35808 23588
rect 35860 23576 35866 23588
rect 36081 23579 36139 23585
rect 36081 23576 36093 23579
rect 35860 23548 36093 23576
rect 35860 23536 35866 23548
rect 36081 23545 36093 23548
rect 36127 23545 36139 23579
rect 36081 23539 36139 23545
rect 32766 23508 32772 23520
rect 31726 23480 32772 23508
rect 32766 23468 32772 23480
rect 32824 23508 32830 23520
rect 33594 23508 33600 23520
rect 32824 23480 33600 23508
rect 32824 23468 32830 23480
rect 33594 23468 33600 23480
rect 33652 23468 33658 23520
rect 35618 23468 35624 23520
rect 35676 23508 35682 23520
rect 35894 23508 35900 23520
rect 35676 23480 35900 23508
rect 35676 23468 35682 23480
rect 35894 23468 35900 23480
rect 35952 23468 35958 23520
rect 37090 23468 37096 23520
rect 37148 23508 37154 23520
rect 37461 23511 37519 23517
rect 37461 23508 37473 23511
rect 37148 23480 37473 23508
rect 37148 23468 37154 23480
rect 37461 23477 37473 23480
rect 37507 23477 37519 23511
rect 37461 23471 37519 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 3970 23264 3976 23316
rect 4028 23264 4034 23316
rect 5166 23264 5172 23316
rect 5224 23264 5230 23316
rect 5537 23307 5595 23313
rect 5537 23273 5549 23307
rect 5583 23304 5595 23307
rect 5626 23304 5632 23316
rect 5583 23276 5632 23304
rect 5583 23273 5595 23276
rect 5537 23267 5595 23273
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 10428 23276 12434 23304
rect 3878 23196 3884 23248
rect 3936 23236 3942 23248
rect 6457 23239 6515 23245
rect 3936 23208 5304 23236
rect 3936 23196 3942 23208
rect 4525 23171 4583 23177
rect 4525 23137 4537 23171
rect 4571 23168 4583 23171
rect 5074 23168 5080 23180
rect 4571 23140 5080 23168
rect 4571 23137 4583 23140
rect 4525 23131 4583 23137
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23100 4491 23103
rect 4614 23100 4620 23112
rect 4479 23072 4620 23100
rect 4479 23069 4491 23072
rect 4433 23063 4491 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 5276 23100 5304 23208
rect 6457 23205 6469 23239
rect 6503 23236 6515 23239
rect 6638 23236 6644 23248
rect 6503 23208 6644 23236
rect 6503 23205 6515 23208
rect 6457 23199 6515 23205
rect 6638 23196 6644 23208
rect 6696 23196 6702 23248
rect 5629 23171 5687 23177
rect 5629 23137 5641 23171
rect 5675 23168 5687 23171
rect 5675 23140 6500 23168
rect 5675 23137 5687 23140
rect 5629 23131 5687 23137
rect 6472 23112 6500 23140
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 5276 23072 5365 23100
rect 5353 23069 5365 23072
rect 5399 23100 5411 23103
rect 5718 23100 5724 23112
rect 5399 23072 5724 23100
rect 5399 23069 5411 23072
rect 5353 23063 5411 23069
rect 5718 23060 5724 23072
rect 5776 23100 5782 23112
rect 6365 23103 6423 23109
rect 6365 23100 6377 23103
rect 5776 23072 6377 23100
rect 5776 23060 5782 23072
rect 6365 23069 6377 23072
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 6454 23060 6460 23112
rect 6512 23100 6518 23112
rect 6549 23103 6607 23109
rect 6549 23100 6561 23103
rect 6512 23072 6561 23100
rect 6512 23060 6518 23072
rect 6549 23069 6561 23072
rect 6595 23069 6607 23103
rect 6549 23063 6607 23069
rect 6638 23060 6644 23112
rect 6696 23060 6702 23112
rect 9950 23060 9956 23112
rect 10008 23100 10014 23112
rect 10137 23103 10195 23109
rect 10137 23100 10149 23103
rect 10008 23072 10149 23100
rect 10008 23060 10014 23072
rect 10137 23069 10149 23072
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 4341 23035 4399 23041
rect 4341 23001 4353 23035
rect 4387 23032 4399 23035
rect 4890 23032 4896 23044
rect 4387 23004 4896 23032
rect 4387 23001 4399 23004
rect 4341 22995 4399 23001
rect 4890 22992 4896 23004
rect 4948 22992 4954 23044
rect 6270 22992 6276 23044
rect 6328 23032 6334 23044
rect 6656 23032 6684 23060
rect 6328 23004 6684 23032
rect 6328 22992 6334 23004
rect 6825 22967 6883 22973
rect 6825 22933 6837 22967
rect 6871 22964 6883 22967
rect 7466 22964 7472 22976
rect 6871 22936 7472 22964
rect 6871 22933 6883 22936
rect 6825 22927 6883 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 10152 22964 10180 23063
rect 10318 22992 10324 23044
rect 10376 22992 10382 23044
rect 10428 23041 10456 23276
rect 10689 23239 10747 23245
rect 10689 23205 10701 23239
rect 10735 23205 10747 23239
rect 12406 23236 12434 23276
rect 22278 23264 22284 23316
rect 22336 23304 22342 23316
rect 22741 23307 22799 23313
rect 22741 23304 22753 23307
rect 22336 23276 22753 23304
rect 22336 23264 22342 23276
rect 22741 23273 22753 23276
rect 22787 23273 22799 23307
rect 22741 23267 22799 23273
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22888 23276 22937 23304
rect 22888 23264 22894 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 22925 23267 22983 23273
rect 26234 23264 26240 23316
rect 26292 23264 26298 23316
rect 35897 23307 35955 23313
rect 35897 23273 35909 23307
rect 35943 23304 35955 23307
rect 36262 23304 36268 23316
rect 35943 23276 36268 23304
rect 35943 23273 35955 23276
rect 35897 23267 35955 23273
rect 36262 23264 36268 23276
rect 36320 23264 36326 23316
rect 38194 23264 38200 23316
rect 38252 23264 38258 23316
rect 12529 23239 12587 23245
rect 12529 23236 12541 23239
rect 12406 23208 12541 23236
rect 10689 23199 10747 23205
rect 12529 23205 12541 23208
rect 12575 23236 12587 23239
rect 12575 23208 14320 23236
rect 12575 23205 12587 23208
rect 12529 23199 12587 23205
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10413 23035 10471 23041
rect 10413 23001 10425 23035
rect 10459 23001 10471 23035
rect 10704 23032 10732 23199
rect 11149 23103 11207 23109
rect 11149 23069 11161 23103
rect 11195 23100 11207 23103
rect 12342 23100 12348 23112
rect 11195 23072 12348 23100
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 14292 23109 14320 23208
rect 14642 23196 14648 23248
rect 14700 23236 14706 23248
rect 14921 23239 14979 23245
rect 14921 23236 14933 23239
rect 14700 23208 14933 23236
rect 14700 23196 14706 23208
rect 14921 23205 14933 23208
rect 14967 23205 14979 23239
rect 14921 23199 14979 23205
rect 24670 23196 24676 23248
rect 24728 23236 24734 23248
rect 26878 23236 26884 23248
rect 24728 23208 26884 23236
rect 24728 23196 24734 23208
rect 26878 23196 26884 23208
rect 26936 23196 26942 23248
rect 27341 23239 27399 23245
rect 27341 23205 27353 23239
rect 27387 23236 27399 23239
rect 30098 23236 30104 23248
rect 27387 23208 30104 23236
rect 27387 23205 27399 23208
rect 27341 23199 27399 23205
rect 30098 23196 30104 23208
rect 30156 23196 30162 23248
rect 16574 23128 16580 23180
rect 16632 23128 16638 23180
rect 19978 23128 19984 23180
rect 20036 23128 20042 23180
rect 20254 23128 20260 23180
rect 20312 23168 20318 23180
rect 20349 23171 20407 23177
rect 20349 23168 20361 23171
rect 20312 23140 20361 23168
rect 20312 23128 20318 23140
rect 20349 23137 20361 23140
rect 20395 23137 20407 23171
rect 20349 23131 20407 23137
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 20622 23168 20628 23180
rect 20496 23140 20628 23168
rect 20496 23128 20502 23140
rect 20622 23128 20628 23140
rect 20680 23128 20686 23180
rect 23017 23171 23075 23177
rect 23017 23168 23029 23171
rect 22066 23140 23029 23168
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14550 23100 14556 23112
rect 14323 23072 14556 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 14660 23072 15056 23100
rect 11394 23035 11452 23041
rect 11394 23032 11406 23035
rect 10704 23004 11406 23032
rect 10413 22995 10471 23001
rect 11394 23001 11406 23004
rect 11440 23001 11452 23035
rect 14660 23032 14688 23072
rect 11394 22995 11452 23001
rect 12406 23004 14688 23032
rect 12406 22964 12434 23004
rect 14826 22992 14832 23044
rect 14884 23032 14890 23044
rect 14921 23035 14979 23041
rect 14921 23032 14933 23035
rect 14884 23004 14933 23032
rect 14884 22992 14890 23004
rect 14921 23001 14933 23004
rect 14967 23001 14979 23035
rect 15028 23032 15056 23072
rect 15194 23060 15200 23112
rect 15252 23060 15258 23112
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23100 15899 23103
rect 15930 23100 15936 23112
rect 15887 23072 15936 23100
rect 15887 23069 15899 23072
rect 15841 23063 15899 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 16822 23035 16880 23041
rect 16822 23032 16834 23035
rect 15028 23004 16834 23032
rect 14921 22995 14979 23001
rect 16822 23001 16834 23004
rect 16868 23001 16880 23035
rect 19996 23032 20024 23128
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 22066 23100 22094 23140
rect 23017 23137 23029 23140
rect 23063 23137 23075 23171
rect 23017 23131 23075 23137
rect 25501 23171 25559 23177
rect 25501 23137 25513 23171
rect 25547 23168 25559 23171
rect 28994 23168 29000 23180
rect 25547 23140 29000 23168
rect 25547 23137 25559 23140
rect 25501 23131 25559 23137
rect 28994 23128 29000 23140
rect 29052 23168 29058 23180
rect 29178 23168 29184 23180
rect 29052 23140 29184 23168
rect 29052 23128 29058 23140
rect 29178 23128 29184 23140
rect 29236 23128 29242 23180
rect 29546 23168 29552 23180
rect 29288 23140 29552 23168
rect 20956 23072 22094 23100
rect 22925 23103 22983 23109
rect 20956 23060 20962 23072
rect 22925 23069 22937 23103
rect 22971 23100 22983 23103
rect 24302 23100 24308 23112
rect 22971 23072 24308 23100
rect 22971 23069 22983 23072
rect 22925 23063 22983 23069
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25317 23103 25375 23109
rect 25317 23100 25329 23103
rect 25004 23072 25329 23100
rect 25004 23060 25010 23072
rect 25317 23069 25329 23072
rect 25363 23069 25375 23103
rect 25317 23063 25375 23069
rect 25406 23060 25412 23112
rect 25464 23100 25470 23112
rect 26697 23103 26755 23109
rect 26697 23100 26709 23103
rect 25464 23072 26709 23100
rect 25464 23060 25470 23072
rect 26697 23069 26709 23072
rect 26743 23069 26755 23103
rect 26697 23063 26755 23069
rect 26970 23060 26976 23112
rect 27028 23100 27034 23112
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 27028 23072 27537 23100
rect 27028 23060 27034 23072
rect 27525 23069 27537 23072
rect 27571 23100 27583 23103
rect 27614 23100 27620 23112
rect 27571 23072 27620 23100
rect 27571 23069 27583 23072
rect 27525 23063 27583 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 28810 23060 28816 23112
rect 28868 23100 28874 23112
rect 29288 23100 29316 23140
rect 29546 23128 29552 23140
rect 29604 23168 29610 23180
rect 29604 23140 30236 23168
rect 29604 23128 29610 23140
rect 28868 23072 29316 23100
rect 28868 23060 28874 23072
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 30208 23109 30236 23140
rect 34698 23128 34704 23180
rect 34756 23168 34762 23180
rect 35713 23171 35771 23177
rect 35713 23168 35725 23171
rect 34756 23140 35725 23168
rect 34756 23128 34762 23140
rect 35713 23137 35725 23140
rect 35759 23137 35771 23171
rect 35713 23131 35771 23137
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23069 30251 23103
rect 30193 23063 30251 23069
rect 30558 23060 30564 23112
rect 30616 23060 30622 23112
rect 33042 23060 33048 23112
rect 33100 23100 33106 23112
rect 35345 23103 35403 23109
rect 35345 23100 35357 23103
rect 33100 23072 35357 23100
rect 33100 23060 33106 23072
rect 35345 23069 35357 23072
rect 35391 23069 35403 23103
rect 35345 23063 35403 23069
rect 35621 23103 35679 23109
rect 35621 23069 35633 23103
rect 35667 23069 35679 23103
rect 35621 23063 35679 23069
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 19996 23004 20269 23032
rect 16822 22995 16880 23001
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 10152 22936 12434 22964
rect 14369 22967 14427 22973
rect 14369 22933 14381 22967
rect 14415 22964 14427 22967
rect 15105 22967 15163 22973
rect 15105 22964 15117 22967
rect 14415 22936 15117 22964
rect 14415 22933 14427 22936
rect 14369 22927 14427 22933
rect 15105 22933 15117 22936
rect 15151 22933 15163 22967
rect 15105 22927 15163 22933
rect 15286 22924 15292 22976
rect 15344 22964 15350 22976
rect 15749 22967 15807 22973
rect 15749 22964 15761 22967
rect 15344 22936 15761 22964
rect 15344 22924 15350 22936
rect 15749 22933 15761 22936
rect 15795 22933 15807 22967
rect 15749 22927 15807 22933
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22964 18015 22967
rect 18506 22964 18512 22976
rect 18003 22936 18512 22964
rect 18003 22933 18015 22936
rect 17957 22927 18015 22933
rect 18506 22924 18512 22936
rect 18564 22924 18570 22976
rect 19889 22967 19947 22973
rect 19889 22933 19901 22967
rect 19935 22964 19947 22967
rect 20070 22964 20076 22976
rect 19935 22936 20076 22964
rect 19935 22933 19947 22936
rect 19889 22927 19947 22933
rect 20070 22924 20076 22936
rect 20128 22924 20134 22976
rect 20272 22964 20300 22995
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 21085 23035 21143 23041
rect 21085 23032 21097 23035
rect 20588 23004 21097 23032
rect 20588 22992 20594 23004
rect 21085 23001 21097 23004
rect 21131 23001 21143 23035
rect 21085 22995 21143 23001
rect 21269 23035 21327 23041
rect 21269 23001 21281 23035
rect 21315 23032 21327 23035
rect 21315 23004 22094 23032
rect 21315 23001 21327 23004
rect 21269 22995 21327 23001
rect 21358 22964 21364 22976
rect 20272 22936 21364 22964
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 21450 22924 21456 22976
rect 21508 22924 21514 22976
rect 22066 22964 22094 23004
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 23385 23035 23443 23041
rect 23385 23032 23397 23035
rect 22244 23004 23397 23032
rect 22244 22992 22250 23004
rect 23385 23001 23397 23004
rect 23431 23001 23443 23035
rect 23385 22995 23443 23001
rect 25133 23035 25191 23041
rect 25133 23001 25145 23035
rect 25179 23032 25191 23035
rect 25222 23032 25228 23044
rect 25179 23004 25228 23032
rect 25179 23001 25191 23004
rect 25133 22995 25191 23001
rect 25222 22992 25228 23004
rect 25280 22992 25286 23044
rect 28626 22992 28632 23044
rect 28684 23032 28690 23044
rect 30282 23032 30288 23044
rect 28684 23004 30288 23032
rect 28684 22992 28690 23004
rect 30282 22992 30288 23004
rect 30340 22992 30346 23044
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 35253 23035 35311 23041
rect 35253 23032 35265 23035
rect 34572 23004 35265 23032
rect 34572 22992 34578 23004
rect 35253 23001 35265 23004
rect 35299 23001 35311 23035
rect 35253 22995 35311 23001
rect 35636 22976 35664 23063
rect 36722 23060 36728 23112
rect 36780 23100 36786 23112
rect 37090 23109 37096 23112
rect 36817 23103 36875 23109
rect 36817 23100 36829 23103
rect 36780 23072 36829 23100
rect 36780 23060 36786 23072
rect 36817 23069 36829 23072
rect 36863 23069 36875 23103
rect 37084 23100 37096 23109
rect 37051 23072 37096 23100
rect 36817 23063 36875 23069
rect 37084 23063 37096 23072
rect 37090 23060 37096 23063
rect 37148 23060 37154 23112
rect 22646 22964 22652 22976
rect 22066 22936 22652 22964
rect 22646 22924 22652 22936
rect 22704 22924 22710 22976
rect 25314 22924 25320 22976
rect 25372 22964 25378 22976
rect 25590 22964 25596 22976
rect 25372 22936 25596 22964
rect 25372 22924 25378 22936
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 27890 22924 27896 22976
rect 27948 22964 27954 22976
rect 29086 22964 29092 22976
rect 27948 22936 29092 22964
rect 27948 22924 27954 22936
rect 29086 22924 29092 22936
rect 29144 22924 29150 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 30837 22967 30895 22973
rect 30837 22964 30849 22967
rect 30616 22936 30849 22964
rect 30616 22924 30622 22936
rect 30837 22933 30849 22936
rect 30883 22964 30895 22967
rect 35618 22964 35624 22976
rect 30883 22936 35624 22964
rect 30883 22933 30895 22936
rect 30837 22927 30895 22933
rect 35618 22924 35624 22936
rect 35676 22924 35682 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 5810 22720 5816 22772
rect 5868 22720 5874 22772
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8573 22763 8631 22769
rect 8573 22760 8585 22763
rect 8352 22732 8585 22760
rect 8352 22720 8358 22732
rect 8573 22729 8585 22732
rect 8619 22729 8631 22763
rect 8573 22723 8631 22729
rect 8849 22763 8907 22769
rect 8849 22729 8861 22763
rect 8895 22760 8907 22763
rect 10134 22760 10140 22772
rect 8895 22732 10140 22760
rect 8895 22729 8907 22732
rect 8849 22723 8907 22729
rect 10134 22720 10140 22732
rect 10192 22760 10198 22772
rect 10318 22760 10324 22772
rect 10192 22732 10324 22760
rect 10192 22720 10198 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 19978 22760 19984 22772
rect 11112 22732 19984 22760
rect 11112 22720 11118 22732
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20070 22720 20076 22772
rect 20128 22720 20134 22772
rect 20162 22720 20168 22772
rect 20220 22760 20226 22772
rect 20438 22760 20444 22772
rect 20220 22732 20444 22760
rect 20220 22720 20226 22732
rect 20438 22720 20444 22732
rect 20496 22720 20502 22772
rect 20530 22720 20536 22772
rect 20588 22720 20594 22772
rect 22278 22760 22284 22772
rect 22066 22732 22284 22760
rect 4982 22652 4988 22704
rect 5040 22692 5046 22704
rect 5040 22664 7696 22692
rect 5040 22652 5046 22664
rect 5626 22584 5632 22636
rect 5684 22624 5690 22636
rect 5905 22627 5963 22633
rect 5905 22624 5917 22627
rect 5684 22596 5917 22624
rect 5684 22584 5690 22596
rect 5905 22593 5917 22596
rect 5951 22624 5963 22627
rect 5994 22624 6000 22636
rect 5951 22596 6000 22624
rect 5951 22593 5963 22596
rect 5905 22587 5963 22593
rect 5994 22584 6000 22596
rect 6052 22584 6058 22636
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 7248 22596 7481 22624
rect 7248 22584 7254 22596
rect 7469 22593 7481 22596
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7558 22584 7564 22636
rect 7616 22584 7622 22636
rect 7668 22624 7696 22664
rect 7742 22652 7748 22704
rect 7800 22652 7806 22704
rect 8481 22695 8539 22701
rect 8481 22661 8493 22695
rect 8527 22692 8539 22695
rect 8754 22692 8760 22704
rect 8527 22664 8760 22692
rect 8527 22661 8539 22664
rect 8481 22655 8539 22661
rect 8754 22652 8760 22664
rect 8812 22652 8818 22704
rect 11974 22701 11980 22704
rect 11968 22692 11980 22701
rect 11935 22664 11980 22692
rect 11968 22655 11980 22664
rect 11974 22652 11980 22655
rect 12032 22652 12038 22704
rect 14826 22652 14832 22704
rect 14884 22692 14890 22704
rect 22066 22692 22094 22732
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 24762 22760 24768 22772
rect 24636 22732 24768 22760
rect 24636 22720 24642 22732
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 27338 22760 27344 22772
rect 25700 22732 27344 22760
rect 25700 22692 25728 22732
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 32582 22760 32588 22772
rect 27488 22732 32588 22760
rect 27488 22720 27494 22732
rect 32582 22720 32588 22732
rect 32640 22720 32646 22772
rect 26234 22692 26240 22704
rect 14884 22664 22094 22692
rect 22388 22664 25728 22692
rect 25792 22664 26240 22692
rect 14884 22652 14890 22664
rect 8202 22624 8208 22636
rect 7668 22596 8208 22624
rect 8202 22584 8208 22596
rect 8260 22624 8266 22636
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8260 22596 8677 22624
rect 8260 22584 8266 22596
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22624 11759 22627
rect 12342 22624 12348 22636
rect 11747 22596 12348 22624
rect 11747 22593 11759 22596
rect 11701 22587 11759 22593
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 14458 22584 14464 22636
rect 14516 22584 14522 22636
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 15194 22584 15200 22636
rect 15252 22584 15258 22636
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 14277 22559 14335 22565
rect 14277 22556 14289 22559
rect 14240 22528 14289 22556
rect 14240 22516 14246 22528
rect 14277 22525 14289 22528
rect 14323 22525 14335 22559
rect 14277 22519 14335 22525
rect 8294 22448 8300 22500
rect 8352 22448 8358 22500
rect 15396 22488 15424 22587
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15562 22584 15568 22636
rect 15620 22584 15626 22636
rect 15654 22584 15660 22636
rect 15712 22633 15718 22636
rect 15712 22627 15761 22633
rect 15712 22593 15715 22627
rect 15749 22624 15761 22627
rect 17218 22624 17224 22636
rect 15749 22596 17224 22624
rect 15749 22593 15761 22596
rect 15712 22587 15761 22593
rect 15712 22584 15718 22587
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 18506 22584 18512 22636
rect 18564 22584 18570 22636
rect 18874 22584 18880 22636
rect 18932 22584 18938 22636
rect 18984 22596 19472 22624
rect 15841 22559 15899 22565
rect 15841 22525 15853 22559
rect 15887 22556 15899 22559
rect 16666 22556 16672 22568
rect 15887 22528 16672 22556
rect 15887 22525 15899 22528
rect 15841 22519 15899 22525
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 18984 22556 19012 22596
rect 16960 22528 19012 22556
rect 19337 22559 19395 22565
rect 16850 22488 16856 22500
rect 15396 22460 16856 22488
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 7006 22380 7012 22432
rect 7064 22420 7070 22432
rect 7285 22423 7343 22429
rect 7285 22420 7297 22423
rect 7064 22392 7297 22420
rect 7064 22380 7070 22392
rect 7285 22389 7297 22392
rect 7331 22389 7343 22423
rect 7285 22383 7343 22389
rect 7466 22380 7472 22432
rect 7524 22380 7530 22432
rect 13081 22423 13139 22429
rect 13081 22389 13093 22423
rect 13127 22420 13139 22423
rect 15378 22420 15384 22432
rect 13127 22392 15384 22420
rect 13127 22389 13139 22392
rect 13081 22383 13139 22389
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 15930 22380 15936 22432
rect 15988 22420 15994 22432
rect 16960 22420 16988 22528
rect 19337 22525 19349 22559
rect 19383 22525 19395 22559
rect 19337 22519 19395 22525
rect 15988 22392 16988 22420
rect 19352 22420 19380 22519
rect 19444 22488 19472 22596
rect 20162 22584 20168 22636
rect 20220 22584 20226 22636
rect 22094 22584 22100 22636
rect 22152 22624 22158 22636
rect 22388 22633 22416 22664
rect 22229 22627 22287 22633
rect 22229 22624 22241 22627
rect 22152 22596 22241 22624
rect 22152 22584 22158 22596
rect 22229 22593 22241 22596
rect 22275 22593 22287 22627
rect 22229 22587 22287 22593
rect 22373 22627 22431 22633
rect 22373 22593 22385 22627
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22462 22584 22468 22636
rect 22520 22584 22526 22636
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 22738 22624 22744 22636
rect 22695 22596 22744 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 24486 22584 24492 22636
rect 24544 22584 24550 22636
rect 24670 22584 24676 22636
rect 24728 22584 24734 22636
rect 25682 22584 25688 22636
rect 25740 22584 25746 22636
rect 25792 22633 25820 22664
rect 26234 22652 26240 22664
rect 26292 22652 26298 22704
rect 27982 22652 27988 22704
rect 28040 22652 28046 22704
rect 30006 22692 30012 22704
rect 28276 22664 30012 22692
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22593 25835 22627
rect 25777 22587 25835 22593
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 26510 22624 26516 22636
rect 26200 22596 26516 22624
rect 26200 22584 26206 22596
rect 26510 22584 26516 22596
rect 26568 22624 26574 22636
rect 26568 22596 27568 22624
rect 26568 22584 26574 22596
rect 19981 22559 20039 22565
rect 19981 22525 19993 22559
rect 20027 22556 20039 22559
rect 20714 22556 20720 22568
rect 20027 22528 20720 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20714 22516 20720 22528
rect 20772 22516 20778 22568
rect 24504 22556 24532 22584
rect 24762 22556 24768 22568
rect 24504 22528 24768 22556
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 25700 22556 25728 22584
rect 26234 22556 26240 22568
rect 25700 22528 26240 22556
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 26329 22491 26387 22497
rect 19444 22460 22232 22488
rect 21818 22420 21824 22432
rect 19352 22392 21824 22420
rect 15988 22380 15994 22392
rect 21818 22380 21824 22392
rect 21876 22380 21882 22432
rect 22002 22380 22008 22432
rect 22060 22420 22066 22432
rect 22097 22423 22155 22429
rect 22097 22420 22109 22423
rect 22060 22392 22109 22420
rect 22060 22380 22066 22392
rect 22097 22389 22109 22392
rect 22143 22389 22155 22423
rect 22204 22420 22232 22460
rect 26329 22457 26341 22491
rect 26375 22488 26387 22491
rect 26418 22488 26424 22500
rect 26375 22460 26424 22488
rect 26375 22457 26387 22460
rect 26329 22451 26387 22457
rect 26418 22448 26424 22460
rect 26476 22448 26482 22500
rect 27540 22488 27568 22596
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 28276 22633 28304 22664
rect 30006 22652 30012 22664
rect 30064 22652 30070 22704
rect 31110 22692 31116 22704
rect 30944 22664 31116 22692
rect 27847 22627 27905 22633
rect 27847 22624 27859 22627
rect 27672 22596 27859 22624
rect 27672 22584 27678 22596
rect 27847 22593 27859 22596
rect 27893 22593 27905 22627
rect 27847 22587 27905 22593
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 28260 22627 28318 22633
rect 28260 22593 28272 22627
rect 28306 22593 28318 22627
rect 28260 22587 28318 22593
rect 27706 22516 27712 22568
rect 27764 22556 27770 22568
rect 28092 22556 28120 22587
rect 28350 22584 28356 22636
rect 28408 22584 28414 22636
rect 30944 22633 30972 22664
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 33229 22695 33287 22701
rect 33229 22661 33241 22695
rect 33275 22692 33287 22695
rect 33594 22692 33600 22704
rect 33275 22664 33600 22692
rect 33275 22661 33287 22664
rect 33229 22655 33287 22661
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 30561 22627 30619 22633
rect 30561 22593 30573 22627
rect 30607 22593 30619 22627
rect 30561 22587 30619 22593
rect 30929 22627 30987 22633
rect 30929 22593 30941 22627
rect 30975 22593 30987 22627
rect 30929 22587 30987 22593
rect 27764 22528 28120 22556
rect 27764 22516 27770 22528
rect 30576 22488 30604 22587
rect 31018 22584 31024 22636
rect 31076 22624 31082 22636
rect 31076 22596 31524 22624
rect 31076 22584 31082 22596
rect 31110 22516 31116 22568
rect 31168 22516 31174 22568
rect 31496 22556 31524 22596
rect 31570 22584 31576 22636
rect 31628 22584 31634 22636
rect 33413 22627 33471 22633
rect 33413 22593 33425 22627
rect 33459 22624 33471 22627
rect 33502 22624 33508 22636
rect 33459 22596 33508 22624
rect 33459 22593 33471 22596
rect 33413 22587 33471 22593
rect 33502 22584 33508 22596
rect 33560 22584 33566 22636
rect 37734 22584 37740 22636
rect 37792 22624 37798 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37792 22596 37841 22624
rect 37792 22584 37798 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 32490 22556 32496 22568
rect 31496 22528 32496 22556
rect 32490 22516 32496 22528
rect 32548 22516 32554 22568
rect 33597 22559 33655 22565
rect 33597 22525 33609 22559
rect 33643 22556 33655 22559
rect 33686 22556 33692 22568
rect 33643 22528 33692 22556
rect 33643 22525 33655 22528
rect 33597 22519 33655 22525
rect 33686 22516 33692 22528
rect 33744 22516 33750 22568
rect 38105 22559 38163 22565
rect 38105 22525 38117 22559
rect 38151 22556 38163 22559
rect 39022 22556 39028 22568
rect 38151 22528 39028 22556
rect 38151 22525 38163 22528
rect 38105 22519 38163 22525
rect 39022 22516 39028 22528
rect 39080 22516 39086 22568
rect 31754 22488 31760 22500
rect 27540 22460 31760 22488
rect 31754 22448 31760 22460
rect 31812 22488 31818 22500
rect 32306 22488 32312 22500
rect 31812 22460 32312 22488
rect 31812 22448 31818 22460
rect 32306 22448 32312 22460
rect 32364 22488 32370 22500
rect 33042 22488 33048 22500
rect 32364 22460 33048 22488
rect 32364 22448 32370 22460
rect 33042 22448 33048 22460
rect 33100 22448 33106 22500
rect 25038 22420 25044 22432
rect 22204 22392 25044 22420
rect 22097 22383 22155 22389
rect 25038 22380 25044 22392
rect 25096 22380 25102 22432
rect 25866 22380 25872 22432
rect 25924 22420 25930 22432
rect 27709 22423 27767 22429
rect 27709 22420 27721 22423
rect 25924 22392 27721 22420
rect 25924 22380 25930 22392
rect 27709 22389 27721 22392
rect 27755 22389 27767 22423
rect 27709 22383 27767 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 7190 22176 7196 22228
rect 7248 22176 7254 22228
rect 15470 22216 15476 22228
rect 7300 22188 15476 22216
rect 6822 22108 6828 22160
rect 6880 22148 6886 22160
rect 7300 22148 7328 22188
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 20622 22216 20628 22228
rect 20496 22188 20628 22216
rect 20496 22176 20502 22188
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 27706 22216 27712 22228
rect 25188 22188 27712 22216
rect 25188 22176 25194 22188
rect 27706 22176 27712 22188
rect 27764 22176 27770 22228
rect 27985 22219 28043 22225
rect 27985 22185 27997 22219
rect 28031 22216 28043 22219
rect 28350 22216 28356 22228
rect 28031 22188 28356 22216
rect 28031 22185 28043 22188
rect 27985 22179 28043 22185
rect 28350 22176 28356 22188
rect 28408 22176 28414 22228
rect 31665 22219 31723 22225
rect 31665 22185 31677 22219
rect 31711 22216 31723 22219
rect 31846 22216 31852 22228
rect 31711 22188 31852 22216
rect 31711 22185 31723 22188
rect 31665 22179 31723 22185
rect 31846 22176 31852 22188
rect 31904 22176 31910 22228
rect 32582 22176 32588 22228
rect 32640 22216 32646 22228
rect 35710 22216 35716 22228
rect 32640 22188 35716 22216
rect 32640 22176 32646 22188
rect 35710 22176 35716 22188
rect 35768 22176 35774 22228
rect 6880 22120 7328 22148
rect 6880 22108 6886 22120
rect 13998 22108 14004 22160
rect 14056 22148 14062 22160
rect 14550 22148 14556 22160
rect 14056 22120 14556 22148
rect 14056 22108 14062 22120
rect 14550 22108 14556 22120
rect 14608 22108 14614 22160
rect 15562 22108 15568 22160
rect 15620 22148 15626 22160
rect 15933 22151 15991 22157
rect 15933 22148 15945 22151
rect 15620 22120 15945 22148
rect 15620 22108 15626 22120
rect 15933 22117 15945 22120
rect 15979 22117 15991 22151
rect 15933 22111 15991 22117
rect 23477 22151 23535 22157
rect 23477 22117 23489 22151
rect 23523 22148 23535 22151
rect 23934 22148 23940 22160
rect 23523 22120 23940 22148
rect 23523 22117 23535 22120
rect 23477 22111 23535 22117
rect 23934 22108 23940 22120
rect 23992 22108 23998 22160
rect 27154 22108 27160 22160
rect 27212 22148 27218 22160
rect 27212 22120 27476 22148
rect 27212 22108 27218 22120
rect 4614 22040 4620 22092
rect 4672 22040 4678 22092
rect 6638 22080 6644 22092
rect 6288 22052 6644 22080
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4798 22012 4804 22024
rect 4479 21984 4804 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 6288 22021 6316 22052
rect 6638 22040 6644 22052
rect 6696 22040 6702 22092
rect 6730 22040 6736 22092
rect 6788 22080 6794 22092
rect 8294 22080 8300 22092
rect 6788 22052 8300 22080
rect 6788 22040 6794 22052
rect 6273 22015 6331 22021
rect 6273 21981 6285 22015
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 7561 22015 7619 22021
rect 7561 21981 7573 22015
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 6365 21947 6423 21953
rect 6365 21944 6377 21947
rect 5684 21916 6377 21944
rect 5684 21904 5690 21916
rect 6365 21913 6377 21916
rect 6411 21944 6423 21947
rect 7484 21944 7512 21975
rect 6411 21916 7512 21944
rect 7576 21944 7604 21975
rect 7650 21972 7656 22024
rect 7708 21972 7714 22024
rect 7852 22021 7880 22052
rect 8294 22040 8300 22052
rect 8352 22040 8358 22092
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 16850 22080 16856 22092
rect 14936 22052 16856 22080
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7883 21984 7917 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 14936 22021 14964 22052
rect 16850 22040 16856 22052
rect 16908 22080 16914 22092
rect 17126 22080 17132 22092
rect 16908 22052 17132 22080
rect 16908 22040 16914 22052
rect 17126 22040 17132 22052
rect 17184 22040 17190 22092
rect 23014 22040 23020 22092
rect 23072 22040 23078 22092
rect 25041 22083 25099 22089
rect 25041 22049 25053 22083
rect 25087 22080 25099 22083
rect 25314 22080 25320 22092
rect 25087 22052 25320 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 25314 22040 25320 22052
rect 25372 22080 25378 22092
rect 25372 22052 26188 22080
rect 25372 22040 25378 22052
rect 9585 22015 9643 22021
rect 9585 22012 9597 22015
rect 9180 21984 9597 22012
rect 9180 21972 9186 21984
rect 9585 21981 9597 21984
rect 9631 21981 9643 22015
rect 9585 21975 9643 21981
rect 14895 22015 14964 22021
rect 14895 21981 14907 22015
rect 14941 21984 14964 22015
rect 14941 21981 14953 21984
rect 14895 21975 14953 21981
rect 15010 21972 15016 22024
rect 15068 21972 15074 22024
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 22012 15255 22015
rect 15654 22012 15660 22024
rect 15243 21984 15660 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 16022 21972 16028 22024
rect 16080 21972 16086 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 20717 22015 20775 22021
rect 20717 22012 20729 22015
rect 19484 21984 20729 22012
rect 19484 21972 19490 21984
rect 20717 21981 20729 21984
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 20984 22015 21042 22021
rect 20984 21981 20996 22015
rect 21030 22012 21042 22015
rect 21450 22012 21456 22024
rect 21030 21984 21456 22012
rect 21030 21981 21042 21984
rect 20984 21975 21042 21981
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 22554 21972 22560 22024
rect 22612 22012 22618 22024
rect 23032 22012 23060 22040
rect 26160 22024 26188 22052
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 26844 22052 27384 22080
rect 26844 22040 26850 22052
rect 22612 21984 23060 22012
rect 23109 22015 23167 22021
rect 22612 21972 22618 21984
rect 23109 21981 23121 22015
rect 23155 22012 23167 22015
rect 23566 22012 23572 22024
rect 23155 21984 23572 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 25222 21972 25228 22024
rect 25280 21972 25286 22024
rect 25866 21972 25872 22024
rect 25924 21972 25930 22024
rect 26142 21972 26148 22024
rect 26200 22012 26206 22024
rect 26973 22015 27031 22021
rect 26973 22012 26985 22015
rect 26200 21984 26985 22012
rect 26200 21972 26206 21984
rect 26973 21981 26985 21984
rect 27019 21981 27031 22015
rect 26973 21975 27031 21981
rect 27062 21972 27068 22024
rect 27120 21972 27126 22024
rect 27356 22021 27384 22052
rect 27341 22015 27399 22021
rect 27341 21981 27353 22015
rect 27387 21981 27399 22015
rect 27448 22012 27476 22120
rect 28718 22108 28724 22160
rect 28776 22148 28782 22160
rect 29181 22151 29239 22157
rect 28776 22120 28994 22148
rect 28776 22108 28782 22120
rect 28966 22080 28994 22120
rect 29181 22117 29193 22151
rect 29227 22148 29239 22151
rect 29270 22148 29276 22160
rect 29227 22120 29276 22148
rect 29227 22117 29239 22120
rect 29181 22111 29239 22117
rect 29270 22108 29276 22120
rect 29328 22108 29334 22160
rect 29914 22108 29920 22160
rect 29972 22108 29978 22160
rect 29932 22080 29960 22108
rect 30466 22080 30472 22092
rect 28920 22052 29960 22080
rect 30024 22052 30472 22080
rect 27801 22015 27859 22021
rect 27801 22012 27813 22015
rect 27448 21984 27813 22012
rect 27341 21975 27399 21981
rect 27801 21981 27813 21984
rect 27847 21981 27859 22015
rect 27801 21975 27859 21981
rect 27982 21972 27988 22024
rect 28040 21972 28046 22024
rect 28534 21972 28540 22024
rect 28592 21972 28598 22024
rect 28630 22015 28688 22021
rect 28630 21981 28642 22015
rect 28676 21981 28688 22015
rect 28630 21975 28688 21981
rect 8110 21944 8116 21956
rect 7576 21916 8116 21944
rect 6411 21913 6423 21916
rect 6365 21907 6423 21913
rect 3970 21836 3976 21888
rect 4028 21836 4034 21888
rect 4338 21836 4344 21888
rect 4396 21836 4402 21888
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 6733 21879 6791 21885
rect 6733 21876 6745 21879
rect 6604 21848 6745 21876
rect 6604 21836 6610 21848
rect 6733 21845 6745 21848
rect 6779 21845 6791 21879
rect 7484 21876 7512 21916
rect 8110 21904 8116 21916
rect 8168 21904 8174 21956
rect 9852 21947 9910 21953
rect 9852 21913 9864 21947
rect 9898 21944 9910 21947
rect 9950 21944 9956 21956
rect 9898 21916 9956 21944
rect 9898 21913 9910 21916
rect 9852 21907 9910 21913
rect 9950 21904 9956 21916
rect 10008 21904 10014 21956
rect 15105 21947 15163 21953
rect 15105 21913 15117 21947
rect 15151 21944 15163 21947
rect 15562 21944 15568 21956
rect 15151 21916 15568 21944
rect 15151 21913 15163 21916
rect 15105 21907 15163 21913
rect 15562 21904 15568 21916
rect 15620 21904 15626 21956
rect 23290 21904 23296 21956
rect 23348 21944 23354 21956
rect 27157 21947 27215 21953
rect 27157 21944 27169 21947
rect 23348 21916 27169 21944
rect 23348 21904 23354 21916
rect 27157 21913 27169 21916
rect 27203 21944 27215 21947
rect 27614 21944 27620 21956
rect 27203 21916 27620 21944
rect 27203 21913 27215 21916
rect 27157 21907 27215 21913
rect 27614 21904 27620 21916
rect 27672 21944 27678 21956
rect 28074 21944 28080 21956
rect 27672 21916 28080 21944
rect 27672 21904 27678 21916
rect 28074 21904 28080 21916
rect 28132 21904 28138 21956
rect 28645 21944 28673 21975
rect 28718 21972 28724 22024
rect 28776 22012 28782 22024
rect 28920 22021 28948 22052
rect 29086 22021 29092 22024
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 28776 21984 28825 22012
rect 28776 21972 28782 21984
rect 28813 21981 28825 21984
rect 28859 21981 28871 22015
rect 28813 21975 28871 21981
rect 28902 22015 28960 22021
rect 28902 21981 28914 22015
rect 28948 21981 28960 22015
rect 28902 21975 28960 21981
rect 29043 22015 29092 22021
rect 29043 21981 29055 22015
rect 29089 21981 29092 22015
rect 29043 21975 29092 21981
rect 29086 21972 29092 21975
rect 29144 21972 29150 22024
rect 29178 21972 29184 22024
rect 29236 22012 29242 22024
rect 30024 22021 30052 22052
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 33226 22080 33232 22092
rect 30576 22052 33232 22080
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29236 21984 29929 22012
rect 29236 21972 29242 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 29917 21975 29975 21981
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 21981 30067 22015
rect 30009 21975 30067 21981
rect 30285 22015 30343 22021
rect 30285 21981 30297 22015
rect 30331 22012 30343 22015
rect 30374 22012 30380 22024
rect 30331 21984 30380 22012
rect 30331 21981 30343 21984
rect 30285 21975 30343 21981
rect 30374 21972 30380 21984
rect 30432 21972 30438 22024
rect 30101 21947 30159 21953
rect 28645 21916 30052 21944
rect 10870 21876 10876 21888
rect 7484 21848 10876 21876
rect 6733 21839 6791 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 10962 21836 10968 21888
rect 11020 21836 11026 21888
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 15381 21879 15439 21885
rect 15381 21876 15393 21879
rect 14700 21848 15393 21876
rect 14700 21836 14706 21848
rect 15381 21845 15393 21848
rect 15427 21845 15439 21879
rect 15381 21839 15439 21845
rect 15746 21836 15752 21888
rect 15804 21876 15810 21888
rect 16390 21876 16396 21888
rect 15804 21848 16396 21876
rect 15804 21836 15810 21848
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 22097 21879 22155 21885
rect 22097 21876 22109 21879
rect 20220 21848 22109 21876
rect 20220 21836 20226 21848
rect 22097 21845 22109 21848
rect 22143 21876 22155 21879
rect 25038 21876 25044 21888
rect 22143 21848 25044 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 25038 21836 25044 21848
rect 25096 21836 25102 21888
rect 25682 21836 25688 21888
rect 25740 21876 25746 21888
rect 25777 21879 25835 21885
rect 25777 21876 25789 21879
rect 25740 21848 25789 21876
rect 25740 21836 25746 21848
rect 25777 21845 25789 21848
rect 25823 21845 25835 21879
rect 25777 21839 25835 21845
rect 26786 21836 26792 21888
rect 26844 21836 26850 21888
rect 27062 21836 27068 21888
rect 27120 21876 27126 21888
rect 29362 21876 29368 21888
rect 27120 21848 29368 21876
rect 27120 21836 27126 21848
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 29638 21836 29644 21888
rect 29696 21876 29702 21888
rect 29733 21879 29791 21885
rect 29733 21876 29745 21879
rect 29696 21848 29745 21876
rect 29696 21836 29702 21848
rect 29733 21845 29745 21848
rect 29779 21845 29791 21879
rect 30024 21876 30052 21916
rect 30101 21913 30113 21947
rect 30147 21944 30159 21947
rect 30190 21944 30196 21956
rect 30147 21916 30196 21944
rect 30147 21913 30159 21916
rect 30101 21907 30159 21913
rect 30190 21904 30196 21916
rect 30248 21904 30254 21956
rect 30576 21876 30604 22052
rect 33226 22040 33232 22052
rect 33284 22040 33290 22092
rect 33594 22040 33600 22092
rect 33652 22040 33658 22092
rect 34054 22040 34060 22092
rect 34112 22040 34118 22092
rect 35621 22083 35679 22089
rect 35621 22049 35633 22083
rect 35667 22080 35679 22083
rect 35710 22080 35716 22092
rect 35667 22052 35716 22080
rect 35667 22049 35679 22052
rect 35621 22043 35679 22049
rect 35710 22040 35716 22052
rect 35768 22040 35774 22092
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 31113 22015 31171 22021
rect 31113 22012 31125 22015
rect 30984 21984 31125 22012
rect 30984 21972 30990 21984
rect 31113 21981 31125 21984
rect 31159 21981 31171 22015
rect 31113 21975 31171 21981
rect 31202 21972 31208 22024
rect 31260 22012 31266 22024
rect 31389 22015 31447 22021
rect 31389 22012 31401 22015
rect 31260 21984 31401 22012
rect 31260 21972 31266 21984
rect 31389 21981 31401 21984
rect 31435 21981 31447 22015
rect 31389 21975 31447 21981
rect 31478 21972 31484 22024
rect 31536 21972 31542 22024
rect 32490 21972 32496 22024
rect 32548 22021 32554 22024
rect 32548 22015 32597 22021
rect 32548 21981 32551 22015
rect 32585 21981 32597 22015
rect 32548 21975 32597 21981
rect 32769 22015 32827 22021
rect 32769 21981 32781 22015
rect 32815 22012 32827 22015
rect 32858 22012 32864 22024
rect 32815 21984 32864 22012
rect 32815 21981 32827 21984
rect 32769 21975 32827 21981
rect 32548 21972 32554 21975
rect 32858 21972 32864 21984
rect 32916 21972 32922 22024
rect 32952 22015 33010 22021
rect 32952 21981 32964 22015
rect 32998 21981 33010 22015
rect 32952 21975 33010 21981
rect 31021 21947 31079 21953
rect 31021 21913 31033 21947
rect 31067 21913 31079 21947
rect 31021 21907 31079 21913
rect 30024 21848 30604 21876
rect 31036 21876 31064 21907
rect 32674 21904 32680 21956
rect 32732 21904 32738 21956
rect 32968 21944 32996 21975
rect 33042 21972 33048 22024
rect 33100 21972 33106 22024
rect 33502 21972 33508 22024
rect 33560 22012 33566 22024
rect 33689 22015 33747 22021
rect 33689 22012 33701 22015
rect 33560 21984 33701 22012
rect 33560 21972 33566 21984
rect 33689 21981 33701 21984
rect 33735 21981 33747 22015
rect 33689 21975 33747 21981
rect 35526 21972 35532 22024
rect 35584 21972 35590 22024
rect 35802 21972 35808 22024
rect 35860 21972 35866 22024
rect 35897 22015 35955 22021
rect 35897 21981 35909 22015
rect 35943 22012 35955 22015
rect 36262 22012 36268 22024
rect 35943 21984 36268 22012
rect 35943 21981 35955 21984
rect 35897 21975 35955 21981
rect 36262 21972 36268 21984
rect 36320 21972 36326 22024
rect 36722 21972 36728 22024
rect 36780 22012 36786 22024
rect 36817 22015 36875 22021
rect 36817 22012 36829 22015
rect 36780 21984 36829 22012
rect 36780 21972 36786 21984
rect 36817 21981 36829 21984
rect 36863 21981 36875 22015
rect 36817 21975 36875 21981
rect 35986 21944 35992 21956
rect 32968 21916 35992 21944
rect 35986 21904 35992 21916
rect 36044 21904 36050 21956
rect 37084 21947 37142 21953
rect 37084 21913 37096 21947
rect 37130 21944 37142 21947
rect 37458 21944 37464 21956
rect 37130 21916 37464 21944
rect 37130 21913 37142 21916
rect 37084 21907 37142 21913
rect 37458 21904 37464 21916
rect 37516 21904 37522 21956
rect 31386 21876 31392 21888
rect 31036 21848 31392 21876
rect 29733 21839 29791 21845
rect 31386 21836 31392 21848
rect 31444 21836 31450 21888
rect 32398 21836 32404 21888
rect 32456 21836 32462 21888
rect 32692 21876 32720 21904
rect 35894 21876 35900 21888
rect 32692 21848 35900 21876
rect 35894 21836 35900 21848
rect 35952 21836 35958 21888
rect 36081 21879 36139 21885
rect 36081 21845 36093 21879
rect 36127 21876 36139 21879
rect 37734 21876 37740 21888
rect 36127 21848 37740 21876
rect 36127 21845 36139 21848
rect 36081 21839 36139 21845
rect 37734 21836 37740 21848
rect 37792 21876 37798 21888
rect 37918 21876 37924 21888
rect 37792 21848 37924 21876
rect 37792 21836 37798 21848
rect 37918 21836 37924 21848
rect 37976 21836 37982 21888
rect 38194 21836 38200 21888
rect 38252 21836 38258 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4338 21632 4344 21684
rect 4396 21672 4402 21684
rect 4433 21675 4491 21681
rect 4433 21672 4445 21675
rect 4396 21644 4445 21672
rect 4396 21632 4402 21644
rect 4433 21641 4445 21644
rect 4479 21672 4491 21675
rect 4479 21644 9628 21672
rect 4479 21641 4491 21644
rect 4433 21635 4491 21641
rect 3320 21607 3378 21613
rect 3320 21573 3332 21607
rect 3366 21604 3378 21607
rect 3970 21604 3976 21616
rect 3366 21576 3976 21604
rect 3366 21573 3378 21576
rect 3320 21567 3378 21573
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 7650 21604 7656 21616
rect 6696 21576 7656 21604
rect 6696 21564 6702 21576
rect 7650 21564 7656 21576
rect 7708 21564 7714 21616
rect 8294 21604 8300 21616
rect 8036 21576 8300 21604
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 5718 21536 5724 21548
rect 5675 21508 5724 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 6178 21496 6184 21548
rect 6236 21536 6242 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6236 21508 6561 21536
rect 6236 21496 6242 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 6822 21496 6828 21548
rect 6880 21496 6886 21548
rect 6914 21496 6920 21548
rect 6972 21496 6978 21548
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 8036 21545 8064 21576
rect 8294 21564 8300 21576
rect 8352 21604 8358 21616
rect 8352 21576 9076 21604
rect 8352 21564 8358 21576
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7064 21508 7941 21536
rect 7064 21496 7070 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 8021 21539 8079 21545
rect 8021 21505 8033 21539
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 8202 21496 8208 21548
rect 8260 21496 8266 21548
rect 9048 21545 9076 21576
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21536 9091 21539
rect 9490 21536 9496 21548
rect 9079 21508 9496 21536
rect 9079 21505 9091 21508
rect 9033 21499 9091 21505
rect 3050 21428 3056 21480
rect 3108 21428 3114 21480
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 4672 21440 5457 21468
rect 4672 21428 4678 21440
rect 5445 21437 5457 21440
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21468 5871 21471
rect 6748 21468 6776 21496
rect 5859 21440 6776 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 8110 21428 8116 21480
rect 8168 21468 8174 21480
rect 8956 21468 8984 21499
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 8168 21440 8984 21468
rect 9600 21468 9628 21644
rect 9950 21632 9956 21684
rect 10008 21632 10014 21684
rect 14458 21632 14464 21684
rect 14516 21632 14522 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 15436 21644 18000 21672
rect 15436 21632 15442 21644
rect 10321 21607 10379 21613
rect 10321 21573 10333 21607
rect 10367 21604 10379 21607
rect 10962 21604 10968 21616
rect 10367 21576 10968 21604
rect 10367 21573 10379 21576
rect 10321 21567 10379 21573
rect 10962 21564 10968 21576
rect 11020 21604 11026 21616
rect 16298 21604 16304 21616
rect 11020 21576 15424 21604
rect 11020 21564 11026 21576
rect 10134 21496 10140 21548
rect 10192 21496 10198 21548
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 10502 21536 10508 21548
rect 10459 21508 10508 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 10612 21508 11008 21536
rect 10612 21468 10640 21508
rect 9600 21440 10640 21468
rect 8168 21428 8174 21440
rect 8956 21400 8984 21440
rect 10870 21428 10876 21480
rect 10928 21428 10934 21480
rect 10980 21468 11008 21508
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11149 21539 11207 21545
rect 11149 21536 11161 21539
rect 11112 21508 11161 21536
rect 11112 21496 11118 21508
rect 11149 21505 11161 21508
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 14458 21496 14464 21548
rect 14516 21496 14522 21548
rect 14642 21496 14648 21548
rect 14700 21496 14706 21548
rect 15396 21468 15424 21576
rect 15856 21576 16304 21604
rect 15856 21545 15884 21576
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 17586 21564 17592 21616
rect 17644 21564 17650 21616
rect 17972 21613 18000 21644
rect 18874 21632 18880 21684
rect 18932 21632 18938 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 24854 21672 24860 21684
rect 22796 21644 24860 21672
rect 22796 21632 22802 21644
rect 17957 21607 18015 21613
rect 17957 21573 17969 21607
rect 18003 21573 18015 21607
rect 17957 21567 18015 21573
rect 18693 21607 18751 21613
rect 18693 21573 18705 21607
rect 18739 21604 18751 21607
rect 19978 21604 19984 21616
rect 18739 21576 19984 21604
rect 18739 21573 18751 21576
rect 18693 21567 18751 21573
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 23155 21613 23183 21644
rect 24854 21632 24860 21644
rect 24912 21632 24918 21684
rect 26418 21632 26424 21684
rect 26476 21672 26482 21684
rect 27246 21672 27252 21684
rect 26476 21644 27252 21672
rect 26476 21632 26482 21644
rect 27246 21632 27252 21644
rect 27304 21672 27310 21684
rect 28534 21672 28540 21684
rect 27304 21644 28540 21672
rect 27304 21632 27310 21644
rect 23140 21607 23198 21613
rect 23140 21573 23152 21607
rect 23186 21573 23198 21607
rect 27522 21604 27528 21616
rect 23140 21567 23198 21573
rect 23400 21576 27528 21604
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16390 21536 16396 21548
rect 15979 21508 16396 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21536 17923 21539
rect 18046 21536 18052 21548
rect 17911 21508 18052 21536
rect 17911 21505 17923 21508
rect 17865 21499 17923 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 18325 21539 18383 21545
rect 18325 21505 18337 21539
rect 18371 21536 18383 21539
rect 19150 21536 19156 21548
rect 18371 21508 19156 21536
rect 18371 21505 18383 21508
rect 18325 21499 18383 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 23400 21545 23428 21576
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 25590 21536 25596 21548
rect 24351 21508 25596 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 25590 21496 25596 21508
rect 25648 21496 25654 21548
rect 26602 21496 26608 21548
rect 26660 21536 26666 21548
rect 27154 21536 27160 21548
rect 26660 21508 27160 21536
rect 26660 21496 26666 21508
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27341 21539 27399 21545
rect 27341 21505 27353 21539
rect 27387 21505 27399 21539
rect 28368 21536 28396 21644
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 28810 21632 28816 21684
rect 28868 21672 28874 21684
rect 29638 21672 29644 21684
rect 28868 21644 29644 21672
rect 28868 21632 28874 21644
rect 29638 21632 29644 21644
rect 29696 21632 29702 21684
rect 29822 21632 29828 21684
rect 29880 21632 29886 21684
rect 29914 21632 29920 21684
rect 29972 21672 29978 21684
rect 32769 21675 32827 21681
rect 32769 21672 32781 21675
rect 29972 21644 32781 21672
rect 29972 21632 29978 21644
rect 32769 21641 32781 21644
rect 32815 21672 32827 21675
rect 35069 21675 35127 21681
rect 35069 21672 35081 21675
rect 32815 21644 35081 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 35069 21641 35081 21644
rect 35115 21672 35127 21675
rect 35526 21672 35532 21684
rect 35115 21644 35532 21672
rect 35115 21641 35127 21644
rect 35069 21635 35127 21641
rect 35526 21632 35532 21644
rect 35584 21632 35590 21684
rect 36262 21632 36268 21684
rect 36320 21632 36326 21684
rect 37458 21632 37464 21684
rect 37516 21632 37522 21684
rect 37918 21632 37924 21684
rect 37976 21632 37982 21684
rect 28442 21564 28448 21616
rect 28500 21604 28506 21616
rect 29840 21604 29868 21632
rect 30098 21604 30104 21616
rect 28500 21576 29040 21604
rect 28500 21564 28506 21576
rect 29012 21545 29040 21576
rect 29748 21576 30104 21604
rect 29748 21545 29776 21576
rect 30098 21564 30104 21576
rect 30156 21564 30162 21616
rect 30558 21564 30564 21616
rect 30616 21604 30622 21616
rect 31202 21604 31208 21616
rect 30616 21576 31208 21604
rect 30616 21564 30622 21576
rect 31202 21564 31208 21576
rect 31260 21564 31266 21616
rect 32398 21564 32404 21616
rect 32456 21604 32462 21616
rect 32585 21607 32643 21613
rect 32585 21604 32597 21607
rect 32456 21576 32597 21604
rect 32456 21564 32462 21576
rect 32585 21573 32597 21576
rect 32631 21573 32643 21607
rect 32585 21567 32643 21573
rect 33956 21607 34014 21613
rect 33956 21573 33968 21607
rect 34002 21604 34014 21607
rect 34054 21604 34060 21616
rect 34002 21576 34060 21604
rect 34002 21573 34014 21576
rect 33956 21567 34014 21573
rect 34054 21564 34060 21576
rect 34112 21564 34118 21616
rect 34606 21564 34612 21616
rect 34664 21604 34670 21616
rect 35897 21607 35955 21613
rect 35897 21604 35909 21607
rect 34664 21576 35909 21604
rect 34664 21564 34670 21576
rect 35897 21573 35909 21576
rect 35943 21573 35955 21607
rect 35897 21567 35955 21573
rect 35986 21564 35992 21616
rect 36044 21604 36050 21616
rect 37829 21607 37887 21613
rect 37829 21604 37841 21607
rect 36044 21576 37841 21604
rect 36044 21564 36050 21576
rect 37829 21573 37841 21576
rect 37875 21604 37887 21607
rect 38194 21604 38200 21616
rect 37875 21576 38200 21604
rect 37875 21573 37887 21576
rect 37829 21567 37887 21573
rect 38194 21564 38200 21576
rect 38252 21564 38258 21616
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 28368 21508 28733 21536
rect 27341 21499 27399 21505
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 28813 21539 28871 21545
rect 28813 21505 28825 21539
rect 28859 21505 28871 21539
rect 28813 21499 28871 21505
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29089 21539 29147 21545
rect 29089 21505 29101 21539
rect 29135 21536 29147 21539
rect 29733 21539 29791 21545
rect 29135 21508 29592 21536
rect 29135 21505 29147 21508
rect 29089 21499 29147 21505
rect 16022 21468 16028 21480
rect 10980 21440 12434 21468
rect 15396 21440 16028 21468
rect 11057 21403 11115 21409
rect 11057 21400 11069 21403
rect 8956 21372 11069 21400
rect 11057 21369 11069 21372
rect 11103 21369 11115 21403
rect 12406 21400 12434 21440
rect 16022 21428 16028 21440
rect 16080 21468 16086 21480
rect 16209 21471 16267 21477
rect 16209 21468 16221 21471
rect 16080 21440 16221 21468
rect 16080 21428 16086 21440
rect 16209 21437 16221 21440
rect 16255 21437 16267 21471
rect 16209 21431 16267 21437
rect 15930 21400 15936 21412
rect 12406 21372 15936 21400
rect 11057 21363 11115 21369
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 16224 21400 16252 21431
rect 16298 21428 16304 21480
rect 16356 21428 16362 21480
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17000 21440 17434 21468
rect 17000 21428 17006 21440
rect 24486 21428 24492 21480
rect 24544 21428 24550 21480
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 24673 21471 24731 21477
rect 24673 21437 24685 21471
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 24765 21471 24823 21477
rect 24765 21437 24777 21471
rect 24811 21468 24823 21471
rect 24854 21468 24860 21480
rect 24811 21440 24860 21468
rect 24811 21437 24823 21440
rect 24765 21431 24823 21437
rect 16574 21400 16580 21412
rect 16224 21372 16580 21400
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 7098 21292 7104 21344
rect 7156 21292 7162 21344
rect 8386 21292 8392 21344
rect 8444 21292 8450 21344
rect 8938 21292 8944 21344
rect 8996 21292 9002 21344
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 10965 21335 11023 21341
rect 10965 21332 10977 21335
rect 10376 21304 10977 21332
rect 10376 21292 10382 21304
rect 10965 21301 10977 21304
rect 11011 21301 11023 21335
rect 10965 21295 11023 21301
rect 15654 21292 15660 21344
rect 15712 21292 15718 21344
rect 22005 21335 22063 21341
rect 22005 21301 22017 21335
rect 22051 21332 22063 21335
rect 23566 21332 23572 21344
rect 22051 21304 23572 21332
rect 22051 21301 22063 21304
rect 22005 21295 22063 21301
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 24596 21332 24624 21431
rect 24688 21400 24716 21431
rect 24854 21428 24860 21440
rect 24912 21468 24918 21480
rect 27062 21468 27068 21480
rect 24912 21440 27068 21468
rect 24912 21428 24918 21440
rect 27062 21428 27068 21440
rect 27120 21428 27126 21480
rect 27356 21468 27384 21499
rect 27522 21468 27528 21480
rect 27356 21440 27528 21468
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 27890 21428 27896 21480
rect 27948 21468 27954 21480
rect 28828 21468 28856 21499
rect 27948 21440 28856 21468
rect 27948 21428 27954 21440
rect 24688 21372 24808 21400
rect 24780 21344 24808 21372
rect 25038 21360 25044 21412
rect 25096 21400 25102 21412
rect 25096 21372 25912 21400
rect 25096 21360 25102 21372
rect 24670 21332 24676 21344
rect 24596 21304 24676 21332
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 24762 21292 24768 21344
rect 24820 21292 24826 21344
rect 24949 21335 25007 21341
rect 24949 21301 24961 21335
rect 24995 21332 25007 21335
rect 25774 21332 25780 21344
rect 24995 21304 25780 21332
rect 24995 21301 25007 21304
rect 24949 21295 25007 21301
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 25884 21332 25912 21372
rect 27264 21372 27752 21400
rect 27264 21332 27292 21372
rect 25884 21304 27292 21332
rect 27341 21335 27399 21341
rect 27341 21301 27353 21335
rect 27387 21332 27399 21335
rect 27614 21332 27620 21344
rect 27387 21304 27620 21332
rect 27387 21301 27399 21304
rect 27341 21295 27399 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 27724 21332 27752 21372
rect 27982 21360 27988 21412
rect 28040 21400 28046 21412
rect 29362 21400 29368 21412
rect 28040 21372 29368 21400
rect 28040 21360 28046 21372
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 29564 21409 29592 21508
rect 29733 21505 29745 21539
rect 29779 21505 29791 21539
rect 29733 21499 29791 21505
rect 29822 21496 29828 21548
rect 29880 21536 29886 21548
rect 31478 21536 31484 21548
rect 29880 21508 31484 21536
rect 29880 21496 29886 21508
rect 31478 21496 31484 21508
rect 31536 21496 31542 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 32861 21539 32919 21545
rect 32861 21536 32873 21539
rect 32824 21508 32873 21536
rect 32824 21496 32830 21508
rect 32861 21505 32873 21508
rect 32907 21505 32919 21539
rect 32861 21499 32919 21505
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 35621 21539 35679 21545
rect 35621 21536 35633 21539
rect 34848 21508 35633 21536
rect 34848 21496 34854 21508
rect 35621 21505 35633 21508
rect 35667 21505 35679 21539
rect 35621 21499 35679 21505
rect 35714 21539 35772 21545
rect 35714 21505 35726 21539
rect 35760 21505 35772 21539
rect 36086 21539 36144 21545
rect 36086 21536 36098 21539
rect 35714 21499 35772 21505
rect 35820 21508 36098 21536
rect 30006 21428 30012 21480
rect 30064 21468 30070 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 30064 21440 30113 21468
rect 30064 21428 30070 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 29549 21403 29607 21409
rect 29549 21369 29561 21403
rect 29595 21369 29607 21403
rect 30116 21400 30144 21431
rect 30190 21428 30196 21480
rect 30248 21428 30254 21480
rect 32030 21468 32036 21480
rect 31726 21440 32036 21468
rect 30926 21400 30932 21412
rect 30116 21372 30932 21400
rect 29549 21363 29607 21369
rect 30926 21360 30932 21372
rect 30984 21400 30990 21412
rect 31726 21400 31754 21440
rect 32030 21428 32036 21440
rect 32088 21428 32094 21480
rect 33686 21428 33692 21480
rect 33744 21428 33750 21480
rect 35434 21468 35440 21480
rect 34716 21440 35440 21468
rect 30984 21372 31754 21400
rect 32585 21403 32643 21409
rect 30984 21360 30990 21372
rect 32585 21369 32597 21403
rect 32631 21400 32643 21403
rect 33594 21400 33600 21412
rect 32631 21372 33600 21400
rect 32631 21369 32643 21372
rect 32585 21363 32643 21369
rect 33594 21360 33600 21372
rect 33652 21360 33658 21412
rect 28442 21332 28448 21344
rect 27724 21304 28448 21332
rect 28442 21292 28448 21304
rect 28500 21292 28506 21344
rect 28534 21292 28540 21344
rect 28592 21292 28598 21344
rect 30742 21292 30748 21344
rect 30800 21332 30806 21344
rect 34716 21332 34744 21440
rect 35434 21428 35440 21440
rect 35492 21468 35498 21480
rect 35729 21468 35757 21499
rect 35492 21440 35757 21468
rect 35492 21428 35498 21440
rect 35342 21360 35348 21412
rect 35400 21400 35406 21412
rect 35820 21400 35848 21508
rect 36086 21505 36098 21508
rect 36132 21505 36144 21539
rect 36086 21499 36144 21505
rect 38010 21428 38016 21480
rect 38068 21428 38074 21480
rect 35400 21372 35848 21400
rect 35400 21360 35406 21372
rect 30800 21304 34744 21332
rect 30800 21292 30806 21304
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 5997 21131 6055 21137
rect 5997 21097 6009 21131
rect 6043 21128 6055 21131
rect 6822 21128 6828 21140
rect 6043 21100 6828 21128
rect 6043 21097 6055 21100
rect 5997 21091 6055 21097
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 7650 21088 7656 21140
rect 7708 21128 7714 21140
rect 9677 21131 9735 21137
rect 9677 21128 9689 21131
rect 7708 21100 9689 21128
rect 7708 21088 7714 21100
rect 9677 21097 9689 21100
rect 9723 21128 9735 21131
rect 9723 21100 10548 21128
rect 9723 21097 9735 21100
rect 9677 21091 9735 21097
rect 3050 20884 3056 20936
rect 3108 20924 3114 20936
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 3108 20896 4629 20924
rect 3108 20884 3114 20896
rect 4617 20893 4629 20896
rect 4663 20924 4675 20927
rect 5442 20924 5448 20936
rect 4663 20896 5448 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 5442 20884 5448 20896
rect 5500 20884 5506 20936
rect 10318 20884 10324 20936
rect 10376 20884 10382 20936
rect 10520 20933 10548 21100
rect 10612 21100 12434 21128
rect 10612 20933 10640 21100
rect 12406 21060 12434 21100
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 15933 21131 15991 21137
rect 15933 21128 15945 21131
rect 15252 21100 15945 21128
rect 15252 21088 15258 21100
rect 15933 21097 15945 21100
rect 15979 21097 15991 21131
rect 15933 21091 15991 21097
rect 16666 21088 16672 21140
rect 16724 21088 16730 21140
rect 26694 21128 26700 21140
rect 20916 21100 26700 21128
rect 12713 21063 12771 21069
rect 12713 21060 12725 21063
rect 12406 21032 12725 21060
rect 12713 21029 12725 21032
rect 12759 21060 12771 21063
rect 12759 21032 13216 21060
rect 12759 21029 12771 21032
rect 12713 21023 12771 21029
rect 11054 20992 11060 21004
rect 10704 20964 11060 20992
rect 10704 20933 10732 20964
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 10505 20927 10563 20933
rect 10505 20893 10517 20927
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20893 10655 20927
rect 10597 20887 10655 20893
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20893 10747 20927
rect 11146 20924 11152 20936
rect 10689 20887 10747 20893
rect 10796 20896 11152 20924
rect 4884 20859 4942 20865
rect 4884 20825 4896 20859
rect 4930 20856 4942 20859
rect 7098 20856 7104 20868
rect 4930 20828 7104 20856
rect 4930 20825 4942 20828
rect 4884 20819 4942 20825
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 9490 20816 9496 20868
rect 9548 20816 9554 20868
rect 9709 20859 9767 20865
rect 9709 20825 9721 20859
rect 9755 20856 9767 20859
rect 10336 20856 10364 20884
rect 9755 20828 10364 20856
rect 9755 20825 9767 20828
rect 9709 20819 9767 20825
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10796 20788 10824 20896
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20924 11391 20927
rect 11422 20924 11428 20936
rect 11379 20896 11428 20924
rect 11379 20893 11391 20896
rect 11333 20887 11391 20893
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 13188 20924 13216 21032
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 20916 21069 20944 21100
rect 26694 21088 26700 21100
rect 26752 21128 26758 21140
rect 27430 21128 27436 21140
rect 26752 21100 27436 21128
rect 26752 21088 26758 21100
rect 27430 21088 27436 21100
rect 27488 21088 27494 21140
rect 28261 21131 28319 21137
rect 28261 21128 28273 21131
rect 27540 21100 28273 21128
rect 20901 21063 20959 21069
rect 20901 21060 20913 21063
rect 14332 21032 20913 21060
rect 14332 21020 14338 21032
rect 20901 21029 20913 21032
rect 20947 21029 20959 21063
rect 20901 21023 20959 21029
rect 21542 21020 21548 21072
rect 21600 21060 21606 21072
rect 21600 21032 26556 21060
rect 21600 21020 21606 21032
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15473 20995 15531 21001
rect 15473 20992 15485 20995
rect 14967 20964 15485 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15473 20961 15485 20964
rect 15519 20961 15531 20995
rect 15473 20955 15531 20961
rect 15580 20964 16160 20992
rect 15580 20924 15608 20964
rect 13188 20896 15608 20924
rect 15654 20884 15660 20936
rect 15712 20884 15718 20936
rect 15749 20927 15807 20933
rect 15749 20893 15761 20927
rect 15795 20924 15807 20927
rect 15838 20924 15844 20936
rect 15795 20896 15844 20924
rect 15795 20893 15807 20896
rect 15749 20887 15807 20893
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 16025 20927 16083 20933
rect 16025 20924 16037 20927
rect 15948 20896 16037 20924
rect 11578 20859 11636 20865
rect 11578 20856 11590 20859
rect 10888 20828 11590 20856
rect 10888 20797 10916 20828
rect 11578 20825 11590 20828
rect 11624 20825 11636 20859
rect 11578 20819 11636 20825
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 14642 20856 14648 20868
rect 14516 20828 14648 20856
rect 14516 20816 14522 20828
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 9907 20760 10824 20788
rect 10873 20791 10931 20797
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10873 20757 10885 20791
rect 10919 20757 10931 20791
rect 10873 20751 10931 20757
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 12066 20788 12072 20800
rect 11112 20760 12072 20788
rect 11112 20748 11118 20760
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13872 20760 14289 20788
rect 13872 20748 13878 20760
rect 14277 20757 14289 20760
rect 14323 20757 14335 20791
rect 14277 20751 14335 20757
rect 14734 20748 14740 20800
rect 14792 20748 14798 20800
rect 15948 20788 15976 20896
rect 16025 20893 16037 20896
rect 16071 20893 16083 20927
rect 16132 20924 16160 20964
rect 16574 20952 16580 21004
rect 16632 20992 16638 21004
rect 16632 20964 16896 20992
rect 16632 20952 16638 20964
rect 16868 20933 16896 20964
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22186 20992 22192 21004
rect 22060 20964 22192 20992
rect 22060 20952 22066 20964
rect 22186 20952 22192 20964
rect 22244 20952 22250 21004
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 22462 20992 22468 21004
rect 22336 20964 22468 20992
rect 22336 20952 22342 20964
rect 22462 20952 22468 20964
rect 22520 20992 22526 21004
rect 22520 20964 23336 20992
rect 22520 20952 22526 20964
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16132 20896 16773 20924
rect 16025 20887 16083 20893
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 16776 20856 16804 20887
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 23057 20927 23115 20933
rect 23057 20924 23069 20927
rect 22480 20896 23069 20924
rect 17034 20856 17040 20868
rect 16776 20828 17040 20856
rect 17034 20816 17040 20828
rect 17092 20816 17098 20868
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 22480 20856 22508 20896
rect 23057 20893 23069 20896
rect 23103 20893 23115 20927
rect 23057 20887 23115 20893
rect 23198 20884 23204 20936
rect 23256 20884 23262 20936
rect 23308 20933 23336 20964
rect 26142 20952 26148 21004
rect 26200 20952 26206 21004
rect 23293 20927 23351 20933
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 22922 20865 22928 20868
rect 22152 20828 22508 20856
rect 22908 20859 22928 20865
rect 22152 20816 22158 20828
rect 22908 20825 22920 20859
rect 22908 20819 22928 20825
rect 22922 20816 22928 20819
rect 22980 20816 22986 20868
rect 23492 20856 23520 20887
rect 24486 20884 24492 20936
rect 24544 20924 24550 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24544 20896 24593 20924
rect 24544 20884 24550 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24946 20924 24952 20936
rect 24811 20896 24952 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 25038 20884 25044 20936
rect 25096 20884 25102 20936
rect 26418 20884 26424 20936
rect 26476 20884 26482 20936
rect 26436 20856 26464 20884
rect 23492 20828 26464 20856
rect 26528 20856 26556 21032
rect 27157 20927 27215 20933
rect 27157 20893 27169 20927
rect 27203 20924 27215 20927
rect 27540 20924 27568 21100
rect 28261 21097 28273 21100
rect 28307 21097 28319 21131
rect 28261 21091 28319 21097
rect 29638 21088 29644 21140
rect 29696 21128 29702 21140
rect 31294 21137 31300 21140
rect 31278 21131 31300 21137
rect 29696 21100 29960 21128
rect 29696 21088 29702 21100
rect 27706 21020 27712 21072
rect 27764 21020 27770 21072
rect 29932 21060 29960 21100
rect 31278 21097 31290 21131
rect 31352 21128 31358 21140
rect 31757 21131 31815 21137
rect 31352 21100 31524 21128
rect 31278 21091 31300 21097
rect 31294 21088 31300 21091
rect 31352 21088 31358 21100
rect 31386 21060 31392 21072
rect 29932 21032 31392 21060
rect 31386 21020 31392 21032
rect 31444 21020 31450 21072
rect 31496 21060 31524 21100
rect 31757 21097 31769 21131
rect 31803 21128 31815 21131
rect 32582 21128 32588 21140
rect 31803 21100 32588 21128
rect 31803 21097 31815 21100
rect 31757 21091 31815 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 35802 21088 35808 21140
rect 35860 21128 35866 21140
rect 36081 21131 36139 21137
rect 36081 21128 36093 21131
rect 35860 21100 36093 21128
rect 35860 21088 35866 21100
rect 36081 21097 36093 21100
rect 36127 21097 36139 21131
rect 36081 21091 36139 21097
rect 31846 21060 31852 21072
rect 31496 21032 31852 21060
rect 31846 21020 31852 21032
rect 31904 21020 31910 21072
rect 35894 21060 35900 21072
rect 35544 21032 35900 21060
rect 27724 20992 27752 21020
rect 27724 20964 27936 20992
rect 27203 20896 27568 20924
rect 27203 20893 27215 20896
rect 27157 20887 27215 20893
rect 27614 20884 27620 20936
rect 27672 20884 27678 20936
rect 27706 20884 27712 20936
rect 27764 20924 27770 20936
rect 27908 20933 27936 20964
rect 29362 20952 29368 21004
rect 29420 20992 29426 21004
rect 29546 20992 29552 21004
rect 29420 20964 29552 20992
rect 29420 20952 29426 20964
rect 29546 20952 29552 20964
rect 29604 20992 29610 21004
rect 29604 20964 29868 20992
rect 29604 20952 29610 20964
rect 27893 20927 27951 20933
rect 27764 20896 27809 20924
rect 27764 20884 27770 20896
rect 27893 20893 27905 20927
rect 27939 20893 27951 20927
rect 27893 20887 27951 20893
rect 27982 20884 27988 20936
rect 28040 20884 28046 20936
rect 28074 20884 28080 20936
rect 28132 20933 28138 20936
rect 28132 20924 28140 20933
rect 28132 20896 28177 20924
rect 28132 20887 28140 20896
rect 28132 20884 28138 20887
rect 28350 20884 28356 20936
rect 28408 20924 28414 20936
rect 29454 20924 29460 20936
rect 28408 20896 29460 20924
rect 28408 20884 28414 20896
rect 29454 20884 29460 20896
rect 29512 20884 29518 20936
rect 29840 20924 29868 20964
rect 30650 20952 30656 21004
rect 30708 20992 30714 21004
rect 30834 20992 30840 21004
rect 30708 20964 30840 20992
rect 30708 20952 30714 20964
rect 30834 20952 30840 20964
rect 30892 20992 30898 21004
rect 31481 20995 31539 21001
rect 31481 20992 31493 20995
rect 30892 20964 31493 20992
rect 30892 20952 30898 20964
rect 31481 20961 31493 20964
rect 31527 20961 31539 20995
rect 31481 20955 31539 20961
rect 31570 20952 31576 21004
rect 31628 20992 31634 21004
rect 34514 20992 34520 21004
rect 31628 20964 34520 20992
rect 31628 20952 31634 20964
rect 34514 20952 34520 20964
rect 34572 20992 34578 21004
rect 35544 21001 35572 21032
rect 35894 21020 35900 21032
rect 35952 21020 35958 21072
rect 35437 20995 35495 21001
rect 35437 20992 35449 20995
rect 34572 20964 35449 20992
rect 34572 20952 34578 20964
rect 35437 20961 35449 20964
rect 35483 20961 35495 20995
rect 35437 20955 35495 20961
rect 35529 20995 35587 21001
rect 35529 20961 35541 20995
rect 35575 20961 35587 20995
rect 35529 20955 35587 20961
rect 34698 20924 34704 20936
rect 29840 20896 34704 20924
rect 34698 20884 34704 20896
rect 34756 20884 34762 20936
rect 35618 20884 35624 20936
rect 35676 20924 35682 20936
rect 35805 20927 35863 20933
rect 35805 20924 35817 20927
rect 35676 20896 35817 20924
rect 35676 20884 35682 20896
rect 35805 20893 35817 20896
rect 35851 20893 35863 20927
rect 35805 20887 35863 20893
rect 35897 20927 35955 20933
rect 35897 20893 35909 20927
rect 35943 20893 35955 20927
rect 35897 20887 35955 20893
rect 31113 20859 31171 20865
rect 31113 20856 31125 20859
rect 26528 20828 28994 20856
rect 16022 20788 16028 20800
rect 15948 20760 16028 20788
rect 16022 20748 16028 20760
rect 16080 20788 16086 20800
rect 16485 20791 16543 20797
rect 16485 20788 16497 20791
rect 16080 20760 16497 20788
rect 16080 20748 16086 20760
rect 16485 20757 16497 20760
rect 16531 20757 16543 20791
rect 16485 20751 16543 20757
rect 17586 20748 17592 20800
rect 17644 20788 17650 20800
rect 23106 20788 23112 20800
rect 17644 20760 23112 20788
rect 17644 20748 17650 20760
rect 23106 20748 23112 20760
rect 23164 20748 23170 20800
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24912 20760 24961 20788
rect 24912 20748 24918 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 26878 20748 26884 20800
rect 26936 20788 26942 20800
rect 27065 20791 27123 20797
rect 27065 20788 27077 20791
rect 26936 20760 27077 20788
rect 26936 20748 26942 20760
rect 27065 20757 27077 20760
rect 27111 20757 27123 20791
rect 28966 20788 28994 20828
rect 29288 20828 31125 20856
rect 29288 20788 29316 20828
rect 31113 20825 31125 20828
rect 31159 20856 31171 20859
rect 31478 20856 31484 20868
rect 31159 20828 31484 20856
rect 31159 20825 31171 20828
rect 31113 20819 31171 20825
rect 31478 20816 31484 20828
rect 31536 20816 31542 20868
rect 35710 20816 35716 20868
rect 35768 20856 35774 20868
rect 35912 20856 35940 20887
rect 37734 20884 37740 20936
rect 37792 20924 37798 20936
rect 37829 20927 37887 20933
rect 37829 20924 37841 20927
rect 37792 20896 37841 20924
rect 37792 20884 37798 20896
rect 37829 20893 37841 20896
rect 37875 20893 37887 20927
rect 37829 20887 37887 20893
rect 35768 20828 35940 20856
rect 38105 20859 38163 20865
rect 35768 20816 35774 20828
rect 38105 20825 38117 20859
rect 38151 20856 38163 20859
rect 39022 20856 39028 20868
rect 38151 20828 39028 20856
rect 38151 20825 38163 20828
rect 38105 20819 38163 20825
rect 39022 20816 39028 20828
rect 39080 20816 39086 20868
rect 28966 20760 29316 20788
rect 27065 20751 27123 20757
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 29822 20788 29828 20800
rect 29420 20760 29828 20788
rect 29420 20748 29426 20760
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 6880 20556 7941 20584
rect 6880 20544 6886 20556
rect 7929 20553 7941 20556
rect 7975 20584 7987 20587
rect 14369 20587 14427 20593
rect 7975 20556 14320 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 9122 20516 9128 20528
rect 5592 20488 9128 20516
rect 5592 20476 5598 20488
rect 6564 20457 6592 20488
rect 9122 20476 9128 20488
rect 9180 20476 9186 20528
rect 13256 20519 13314 20525
rect 13256 20485 13268 20519
rect 13302 20516 13314 20519
rect 13814 20516 13820 20528
rect 13302 20488 13820 20516
rect 13302 20485 13314 20488
rect 13256 20479 13314 20485
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 14292 20516 14320 20556
rect 14369 20553 14381 20587
rect 14415 20584 14427 20587
rect 14458 20584 14464 20596
rect 14415 20556 14464 20584
rect 14415 20553 14427 20556
rect 14369 20547 14427 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 14792 20556 14933 20584
rect 14792 20544 14798 20556
rect 14921 20553 14933 20556
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 19702 20584 19708 20596
rect 15620 20556 19708 20584
rect 15620 20544 15626 20556
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20036 20556 20821 20584
rect 20036 20544 20042 20556
rect 20809 20553 20821 20556
rect 20855 20584 20867 20587
rect 20855 20556 27292 20584
rect 20855 20553 20867 20556
rect 20809 20547 20867 20553
rect 16666 20516 16672 20528
rect 14292 20488 16672 20516
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 19242 20516 19248 20528
rect 18524 20488 19248 20516
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6816 20451 6874 20457
rect 6816 20417 6828 20451
rect 6862 20448 6874 20451
rect 7098 20448 7104 20460
rect 6862 20420 7104 20448
rect 6862 20417 6874 20420
rect 6816 20411 6874 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20448 17463 20451
rect 17586 20448 17592 20460
rect 17451 20420 17592 20448
rect 17451 20417 17463 20420
rect 17405 20411 17463 20417
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 18524 20457 18552 20488
rect 19242 20476 19248 20488
rect 19300 20516 19306 20528
rect 19300 20488 19840 20516
rect 19300 20476 19306 20488
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 19426 20408 19432 20460
rect 19484 20408 19490 20460
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19685 20451 19743 20457
rect 19685 20448 19697 20451
rect 19576 20420 19697 20448
rect 19576 20408 19582 20420
rect 19685 20417 19697 20420
rect 19731 20417 19743 20451
rect 19812 20448 19840 20488
rect 20070 20476 20076 20528
rect 20128 20516 20134 20528
rect 22554 20516 22560 20528
rect 20128 20488 20576 20516
rect 20128 20476 20134 20488
rect 20548 20448 20576 20488
rect 22066 20488 22560 20516
rect 22066 20448 22094 20488
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 23106 20476 23112 20528
rect 23164 20516 23170 20528
rect 23164 20488 27200 20516
rect 23164 20476 23170 20488
rect 19812 20420 20484 20448
rect 20548 20420 22094 20448
rect 22373 20451 22431 20457
rect 19685 20411 19743 20417
rect 11514 20340 11520 20392
rect 11572 20380 11578 20392
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 11572 20352 13001 20380
rect 11572 20340 11578 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 15378 20340 15384 20392
rect 15436 20340 15442 20392
rect 15562 20340 15568 20392
rect 15620 20340 15626 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16356 20352 17141 20380
rect 16356 20340 16362 20352
rect 17129 20349 17141 20352
rect 17175 20380 17187 20383
rect 18322 20380 18328 20392
rect 17175 20352 18328 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 18322 20340 18328 20352
rect 18380 20340 18386 20392
rect 15930 20272 15936 20324
rect 15988 20312 15994 20324
rect 19242 20312 19248 20324
rect 15988 20284 19248 20312
rect 15988 20272 15994 20284
rect 19242 20272 19248 20284
rect 19300 20272 19306 20324
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17221 20247 17279 20253
rect 17221 20244 17233 20247
rect 17000 20216 17233 20244
rect 17000 20204 17006 20216
rect 17221 20213 17233 20216
rect 17267 20213 17279 20247
rect 17221 20207 17279 20213
rect 17589 20247 17647 20253
rect 17589 20213 17601 20247
rect 17635 20244 17647 20247
rect 19702 20244 19708 20256
rect 17635 20216 19708 20244
rect 17635 20213 17647 20216
rect 17589 20207 17647 20213
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 19794 20204 19800 20256
rect 19852 20244 19858 20256
rect 20346 20244 20352 20256
rect 19852 20216 20352 20244
rect 19852 20204 19858 20216
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 20456 20244 20484 20420
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 22738 20448 22744 20460
rect 22419 20420 22744 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 24578 20408 24584 20460
rect 24636 20408 24642 20460
rect 25038 20408 25044 20460
rect 25096 20448 25102 20460
rect 25501 20451 25559 20457
rect 25501 20448 25513 20451
rect 25096 20420 25513 20448
rect 25096 20408 25102 20420
rect 25501 20417 25513 20420
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25590 20408 25596 20460
rect 25648 20408 25654 20460
rect 27172 20457 27200 20488
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 27157 20451 27215 20457
rect 27157 20417 27169 20451
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 21048 20352 22324 20380
rect 21048 20340 21054 20352
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 22005 20315 22063 20321
rect 22005 20312 22017 20315
rect 20772 20284 22017 20312
rect 20772 20272 20778 20284
rect 22005 20281 22017 20284
rect 22051 20281 22063 20315
rect 22296 20312 22324 20352
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 24765 20383 24823 20389
rect 24765 20349 24777 20383
rect 24811 20349 24823 20383
rect 24765 20343 24823 20349
rect 22572 20312 22600 20343
rect 22296 20284 22600 20312
rect 24780 20312 24808 20343
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 25700 20380 25728 20411
rect 24912 20352 25728 20380
rect 27264 20380 27292 20556
rect 27338 20544 27344 20596
rect 27396 20544 27402 20596
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 28994 20584 29000 20596
rect 27764 20556 29000 20584
rect 27764 20544 27770 20556
rect 28994 20544 29000 20556
rect 29052 20544 29058 20596
rect 33502 20544 33508 20596
rect 33560 20544 33566 20596
rect 27356 20516 27384 20544
rect 27433 20519 27491 20525
rect 27433 20516 27445 20519
rect 27356 20488 27445 20516
rect 27433 20485 27445 20488
rect 27479 20485 27491 20519
rect 27433 20479 27491 20485
rect 28166 20476 28172 20528
rect 28224 20516 28230 20528
rect 31662 20516 31668 20528
rect 28224 20488 31668 20516
rect 28224 20476 28230 20488
rect 31662 20476 31668 20488
rect 31720 20516 31726 20528
rect 35805 20519 35863 20525
rect 31720 20488 35296 20516
rect 31720 20476 31726 20488
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20448 27583 20451
rect 27614 20448 27620 20460
rect 27571 20420 27620 20448
rect 27571 20417 27583 20420
rect 27525 20411 27583 20417
rect 27614 20408 27620 20420
rect 27672 20448 27678 20460
rect 28718 20448 28724 20460
rect 27672 20420 28724 20448
rect 27672 20408 27678 20420
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 28994 20408 29000 20460
rect 29052 20448 29058 20460
rect 29549 20451 29607 20457
rect 29549 20448 29561 20451
rect 29052 20420 29561 20448
rect 29052 20408 29058 20420
rect 29549 20417 29561 20420
rect 29595 20448 29607 20451
rect 29595 20420 30604 20448
rect 29595 20417 29607 20420
rect 29549 20411 29607 20417
rect 27890 20380 27896 20392
rect 27264 20352 27896 20380
rect 24912 20340 24918 20352
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 29273 20383 29331 20389
rect 29273 20349 29285 20383
rect 29319 20380 29331 20383
rect 29730 20380 29736 20392
rect 29319 20352 29736 20380
rect 29319 20349 29331 20352
rect 29273 20343 29331 20349
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 30576 20380 30604 20420
rect 30650 20408 30656 20460
rect 30708 20408 30714 20460
rect 30742 20408 30748 20460
rect 30800 20408 30806 20460
rect 30926 20408 30932 20460
rect 30984 20448 30990 20460
rect 31055 20451 31113 20457
rect 31055 20448 31067 20451
rect 30984 20420 31067 20448
rect 30984 20408 30990 20420
rect 31055 20417 31067 20420
rect 31101 20417 31113 20451
rect 31055 20411 31113 20417
rect 33137 20451 33195 20457
rect 33137 20417 33149 20451
rect 33183 20417 33195 20451
rect 33137 20411 33195 20417
rect 32674 20380 32680 20392
rect 30576 20352 32680 20380
rect 32674 20340 32680 20352
rect 32732 20340 32738 20392
rect 33152 20380 33180 20411
rect 33226 20408 33232 20460
rect 33284 20448 33290 20460
rect 35268 20457 35296 20488
rect 35805 20485 35817 20519
rect 35851 20516 35863 20519
rect 37734 20516 37740 20528
rect 35851 20488 37740 20516
rect 35851 20485 35863 20488
rect 35805 20479 35863 20485
rect 37734 20476 37740 20488
rect 37792 20516 37798 20528
rect 37921 20519 37979 20525
rect 37921 20516 37933 20519
rect 37792 20488 37933 20516
rect 37792 20476 37798 20488
rect 37921 20485 37933 20488
rect 37967 20485 37979 20519
rect 37921 20479 37979 20485
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 33284 20420 33333 20448
rect 33284 20408 33290 20420
rect 33321 20417 33333 20420
rect 33367 20417 33379 20451
rect 33321 20411 33379 20417
rect 35253 20451 35311 20457
rect 35253 20417 35265 20451
rect 35299 20448 35311 20451
rect 35434 20448 35440 20460
rect 35299 20420 35440 20448
rect 35299 20417 35311 20420
rect 35253 20411 35311 20417
rect 35434 20408 35440 20420
rect 35492 20408 35498 20460
rect 35529 20451 35587 20457
rect 35529 20417 35541 20451
rect 35575 20417 35587 20451
rect 35529 20411 35587 20417
rect 33502 20380 33508 20392
rect 33152 20352 33508 20380
rect 33502 20340 33508 20352
rect 33560 20340 33566 20392
rect 33962 20340 33968 20392
rect 34020 20380 34026 20392
rect 35544 20380 35572 20411
rect 35618 20408 35624 20460
rect 35676 20408 35682 20460
rect 37826 20408 37832 20460
rect 37884 20408 37890 20460
rect 34020 20352 35572 20380
rect 34020 20340 34026 20352
rect 38010 20340 38016 20392
rect 38068 20340 38074 20392
rect 24946 20312 24952 20324
rect 24780 20284 24952 20312
rect 22005 20275 22063 20281
rect 24946 20272 24952 20284
rect 25004 20272 25010 20324
rect 29365 20315 29423 20321
rect 29365 20312 29377 20315
rect 25424 20284 29377 20312
rect 25424 20244 25452 20284
rect 29365 20281 29377 20284
rect 29411 20281 29423 20315
rect 29365 20275 29423 20281
rect 31297 20315 31355 20321
rect 31297 20281 31309 20315
rect 31343 20312 31355 20315
rect 31386 20312 31392 20324
rect 31343 20284 31392 20312
rect 31343 20281 31355 20284
rect 31297 20275 31355 20281
rect 31386 20272 31392 20284
rect 31444 20272 31450 20324
rect 20456 20216 25452 20244
rect 27430 20204 27436 20256
rect 27488 20244 27494 20256
rect 27709 20247 27767 20253
rect 27709 20244 27721 20247
rect 27488 20216 27721 20244
rect 27488 20204 27494 20216
rect 27709 20213 27721 20216
rect 27755 20213 27767 20247
rect 27709 20207 27767 20213
rect 29733 20247 29791 20253
rect 29733 20213 29745 20247
rect 29779 20244 29791 20247
rect 29822 20244 29828 20256
rect 29779 20216 29828 20244
rect 29779 20213 29791 20216
rect 29733 20207 29791 20213
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30742 20204 30748 20256
rect 30800 20244 30806 20256
rect 31570 20244 31576 20256
rect 30800 20216 31576 20244
rect 30800 20204 30806 20216
rect 31570 20204 31576 20216
rect 31628 20204 31634 20256
rect 35345 20247 35403 20253
rect 35345 20213 35357 20247
rect 35391 20244 35403 20247
rect 35802 20244 35808 20256
rect 35391 20216 35808 20244
rect 35391 20213 35403 20216
rect 35345 20207 35403 20213
rect 35802 20204 35808 20216
rect 35860 20204 35866 20256
rect 37458 20204 37464 20256
rect 37516 20204 37522 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 7098 20000 7104 20052
rect 7156 20000 7162 20052
rect 15289 20043 15347 20049
rect 7208 20012 12434 20040
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 7208 19972 7236 20012
rect 5684 19944 7236 19972
rect 12406 19972 12434 20012
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 15378 20040 15384 20052
rect 15335 20012 15384 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 16666 20000 16672 20052
rect 16724 20040 16730 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 16724 20012 17141 20040
rect 16724 20000 16730 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 17586 20000 17592 20052
rect 17644 20000 17650 20052
rect 19429 20043 19487 20049
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 19518 20040 19524 20052
rect 19475 20012 19524 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 22002 20040 22008 20052
rect 21652 20012 22008 20040
rect 17402 19972 17408 19984
rect 12406 19944 17408 19972
rect 5684 19932 5690 19944
rect 17402 19932 17408 19944
rect 17460 19932 17466 19984
rect 4614 19864 4620 19916
rect 4672 19864 4678 19916
rect 9122 19864 9128 19916
rect 9180 19864 9186 19916
rect 15933 19907 15991 19913
rect 15933 19873 15945 19907
rect 15979 19904 15991 19907
rect 16022 19904 16028 19916
rect 15979 19876 16028 19904
rect 15979 19873 15991 19876
rect 15933 19867 15991 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 17218 19904 17224 19916
rect 16448 19876 17224 19904
rect 16448 19864 16454 19876
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19836 4583 19839
rect 4706 19836 4712 19848
rect 4571 19808 4712 19836
rect 4571 19805 4583 19808
rect 4525 19799 4583 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6822 19796 6828 19848
rect 6880 19796 6886 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 6972 19808 8125 19836
rect 6972 19796 6978 19808
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8938 19836 8944 19848
rect 8343 19808 8944 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 11698 19796 11704 19848
rect 11756 19796 11762 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14608 19808 14749 19836
rect 14608 19796 14614 19808
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15712 19808 15761 19836
rect 15712 19796 15718 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 17494 19836 17500 19848
rect 17451 19808 17500 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 6730 19728 6736 19780
rect 6788 19728 6794 19780
rect 9214 19728 9220 19780
rect 9272 19768 9278 19780
rect 9370 19771 9428 19777
rect 9370 19768 9382 19771
rect 9272 19740 9382 19768
rect 9272 19728 9278 19740
rect 9370 19737 9382 19740
rect 9416 19737 9428 19771
rect 9370 19731 9428 19737
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11425 19771 11483 19777
rect 11425 19768 11437 19771
rect 11020 19740 11437 19768
rect 11020 19728 11026 19740
rect 11425 19737 11437 19740
rect 11471 19737 11483 19771
rect 14826 19768 14832 19780
rect 11425 19731 11483 19737
rect 12406 19740 14832 19768
rect 4062 19660 4068 19712
rect 4120 19660 4126 19712
rect 4430 19660 4436 19712
rect 4488 19660 4494 19712
rect 6748 19700 6776 19728
rect 6822 19700 6828 19712
rect 6748 19672 6828 19700
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7984 19672 8217 19700
rect 7984 19660 7990 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 8205 19663 8263 19669
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 12406 19700 12434 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15764 19768 15792 19799
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 17604 19836 17632 20000
rect 18509 19975 18567 19981
rect 18509 19941 18521 19975
rect 18555 19972 18567 19975
rect 20990 19972 20996 19984
rect 18555 19944 20996 19972
rect 18555 19941 18567 19944
rect 18509 19935 18567 19941
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 21450 19932 21456 19984
rect 21508 19932 21514 19984
rect 17678 19864 17684 19916
rect 17736 19904 17742 19916
rect 17736 19876 18644 19904
rect 17736 19864 17742 19876
rect 18616 19845 18644 19876
rect 19702 19864 19708 19916
rect 19760 19904 19766 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19760 19876 19993 19904
rect 19760 19864 19766 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 21652 19848 21680 20012
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 24762 20040 24768 20052
rect 22520 20012 24768 20040
rect 22520 20000 22526 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 25038 20000 25044 20052
rect 25096 20000 25102 20052
rect 26510 20000 26516 20052
rect 26568 20000 26574 20052
rect 28626 20000 28632 20052
rect 28684 20000 28690 20052
rect 29822 20000 29828 20052
rect 29880 20000 29886 20052
rect 34606 20000 34612 20052
rect 34664 20040 34670 20052
rect 35158 20040 35164 20052
rect 34664 20012 35164 20040
rect 34664 20000 34670 20012
rect 35158 20000 35164 20012
rect 35216 20000 35222 20052
rect 35529 20043 35587 20049
rect 35529 20009 35541 20043
rect 35575 20040 35587 20043
rect 35618 20040 35624 20052
rect 35575 20012 35624 20040
rect 35575 20009 35587 20012
rect 35529 20003 35587 20009
rect 35618 20000 35624 20012
rect 35676 20000 35682 20052
rect 21744 19944 25452 19972
rect 18233 19839 18291 19845
rect 18233 19836 18245 19839
rect 17604 19808 18245 19836
rect 18233 19805 18245 19808
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20714 19836 20720 19848
rect 19935 19808 20720 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 15930 19768 15936 19780
rect 15764 19740 15936 19768
rect 15930 19728 15936 19740
rect 15988 19728 15994 19780
rect 17126 19728 17132 19780
rect 17184 19728 17190 19780
rect 18340 19768 18368 19799
rect 17420 19740 18368 19768
rect 18616 19768 18644 19799
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 21634 19845 21640 19848
rect 21632 19799 21640 19845
rect 21634 19796 21640 19799
rect 21692 19796 21698 19848
rect 21744 19845 21772 19944
rect 23198 19864 23204 19916
rect 23256 19864 23262 19916
rect 24670 19864 24676 19916
rect 24728 19864 24734 19916
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 19797 19771 19855 19777
rect 18616 19740 19748 19768
rect 17420 19712 17448 19740
rect 10560 19672 12434 19700
rect 14645 19703 14703 19709
rect 10560 19660 10566 19672
rect 14645 19669 14657 19703
rect 14691 19700 14703 19703
rect 14734 19700 14740 19712
rect 14691 19672 14740 19700
rect 14691 19669 14703 19672
rect 14645 19663 14703 19669
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15562 19660 15568 19712
rect 15620 19700 15626 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15620 19672 15669 19700
rect 15620 19660 15626 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 17310 19700 17316 19712
rect 16448 19672 17316 19700
rect 16448 19660 16454 19672
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17402 19660 17408 19712
rect 17460 19660 17466 19712
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 18690 19700 18696 19712
rect 18095 19672 18696 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19720 19700 19748 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 19978 19768 19984 19780
rect 19843 19740 19984 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 21821 19771 21879 19777
rect 21821 19737 21833 19771
rect 21867 19768 21879 19771
rect 21910 19768 21916 19780
rect 21867 19740 21916 19768
rect 21867 19737 21879 19740
rect 21821 19731 21879 19737
rect 21910 19728 21916 19740
rect 21968 19768 21974 19780
rect 22278 19768 22284 19780
rect 21968 19740 22284 19768
rect 21968 19728 21974 19740
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 20254 19700 20260 19712
rect 19720 19672 20260 19700
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 22480 19700 22508 19799
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 22833 19839 22891 19845
rect 22833 19836 22845 19839
rect 22704 19808 22845 19836
rect 22704 19796 22710 19808
rect 22833 19805 22845 19808
rect 22879 19805 22891 19839
rect 22833 19799 22891 19805
rect 23382 19796 23388 19848
rect 23440 19796 23446 19848
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 25424 19768 25452 19944
rect 26234 19932 26240 19984
rect 26292 19972 26298 19984
rect 26624 19975 26682 19981
rect 26624 19972 26636 19975
rect 26292 19944 26636 19972
rect 26292 19932 26298 19944
rect 26624 19941 26636 19944
rect 26670 19941 26682 19975
rect 27614 19972 27620 19984
rect 26624 19935 26682 19941
rect 26804 19944 27620 19972
rect 26421 19907 26479 19913
rect 26421 19873 26433 19907
rect 26467 19904 26479 19907
rect 26510 19904 26516 19916
rect 26467 19876 26516 19904
rect 26467 19873 26479 19876
rect 26421 19867 26479 19873
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 26804 19845 26832 19944
rect 27614 19932 27620 19944
rect 27672 19972 27678 19984
rect 27890 19972 27896 19984
rect 27672 19944 27896 19972
rect 27672 19932 27678 19944
rect 27890 19932 27896 19944
rect 27948 19932 27954 19984
rect 26988 19876 27568 19904
rect 26789 19839 26847 19845
rect 26789 19805 26801 19839
rect 26835 19805 26847 19839
rect 26789 19799 26847 19805
rect 26988 19768 27016 19876
rect 27062 19796 27068 19848
rect 27120 19836 27126 19848
rect 27249 19839 27307 19845
rect 27249 19836 27261 19839
rect 27120 19808 27261 19836
rect 27120 19796 27126 19808
rect 27249 19805 27261 19808
rect 27295 19805 27307 19839
rect 27249 19799 27307 19805
rect 27433 19839 27491 19845
rect 27433 19805 27445 19839
rect 27479 19805 27491 19839
rect 27540 19836 27568 19876
rect 28460 19876 28580 19904
rect 28166 19836 28172 19848
rect 27540 19808 28172 19836
rect 27433 19799 27491 19805
rect 25424 19740 27016 19768
rect 20680 19672 22508 19700
rect 20680 19660 20686 19672
rect 23106 19660 23112 19712
rect 23164 19700 23170 19712
rect 26145 19703 26203 19709
rect 26145 19700 26157 19703
rect 23164 19672 26157 19700
rect 23164 19660 23170 19672
rect 26145 19669 26157 19672
rect 26191 19700 26203 19703
rect 27154 19700 27160 19712
rect 26191 19672 27160 19700
rect 26191 19669 26203 19672
rect 26145 19663 26203 19669
rect 27154 19660 27160 19672
rect 27212 19700 27218 19712
rect 27448 19700 27476 19799
rect 28166 19796 28172 19808
rect 28224 19796 28230 19848
rect 27801 19771 27859 19777
rect 27801 19737 27813 19771
rect 27847 19768 27859 19771
rect 27982 19768 27988 19780
rect 27847 19740 27988 19768
rect 27847 19737 27859 19740
rect 27801 19731 27859 19737
rect 27982 19728 27988 19740
rect 28040 19728 28046 19780
rect 27212 19672 27476 19700
rect 28460 19700 28488 19876
rect 28552 19845 28580 19876
rect 28645 19845 28673 20000
rect 31481 19975 31539 19981
rect 31481 19941 31493 19975
rect 31527 19972 31539 19975
rect 31570 19972 31576 19984
rect 31527 19944 31576 19972
rect 31527 19941 31539 19944
rect 31481 19935 31539 19941
rect 31570 19932 31576 19944
rect 31628 19932 31634 19984
rect 31726 19944 35020 19972
rect 29086 19904 29092 19916
rect 28736 19876 29092 19904
rect 28736 19848 28764 19876
rect 29086 19864 29092 19876
rect 29144 19864 29150 19916
rect 30650 19864 30656 19916
rect 30708 19904 30714 19916
rect 30929 19907 30987 19913
rect 30929 19904 30941 19907
rect 30708 19876 30941 19904
rect 30708 19864 30714 19876
rect 30929 19873 30941 19876
rect 30975 19873 30987 19907
rect 30929 19867 30987 19873
rect 28537 19839 28595 19845
rect 28537 19805 28549 19839
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 28630 19839 28688 19845
rect 28630 19805 28642 19839
rect 28676 19805 28688 19839
rect 28630 19799 28688 19805
rect 28718 19796 28724 19848
rect 28776 19796 28782 19848
rect 28902 19796 28908 19848
rect 28960 19796 28966 19848
rect 28994 19796 29000 19848
rect 29052 19845 29058 19848
rect 29052 19836 29060 19845
rect 29052 19808 29097 19836
rect 29052 19799 29060 19808
rect 29052 19796 29058 19799
rect 29730 19796 29736 19848
rect 29788 19796 29794 19848
rect 29822 19796 29828 19848
rect 29880 19796 29886 19848
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 31726 19836 31754 19944
rect 32490 19864 32496 19916
rect 32548 19904 32554 19916
rect 32548 19876 32817 19904
rect 32548 19864 32554 19876
rect 31036 19808 31754 19836
rect 28813 19771 28871 19777
rect 28813 19737 28825 19771
rect 28859 19737 28871 19771
rect 29932 19768 29960 19796
rect 31036 19780 31064 19808
rect 32214 19796 32220 19848
rect 32272 19836 32278 19848
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 32272 19808 32321 19836
rect 32272 19796 32278 19808
rect 32309 19805 32321 19808
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 32398 19796 32404 19848
rect 32456 19796 32462 19848
rect 32789 19845 32817 19876
rect 33502 19864 33508 19916
rect 33560 19864 33566 19916
rect 33965 19907 34023 19913
rect 33965 19873 33977 19907
rect 34011 19904 34023 19907
rect 34422 19904 34428 19916
rect 34011 19876 34428 19904
rect 34011 19873 34023 19876
rect 33965 19867 34023 19873
rect 34422 19864 34428 19876
rect 34480 19864 34486 19916
rect 32674 19839 32732 19845
rect 32674 19836 32686 19839
rect 32508 19808 32686 19836
rect 28813 19731 28871 19737
rect 29564 19740 29960 19768
rect 28534 19700 28540 19712
rect 28460 19672 28540 19700
rect 27212 19660 27218 19672
rect 28534 19660 28540 19672
rect 28592 19660 28598 19712
rect 28626 19660 28632 19712
rect 28684 19700 28690 19712
rect 28828 19700 28856 19731
rect 28684 19672 28856 19700
rect 28684 19660 28690 19672
rect 29178 19660 29184 19712
rect 29236 19660 29242 19712
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 29564 19700 29592 19740
rect 31018 19728 31024 19780
rect 31076 19728 31082 19780
rect 31205 19771 31263 19777
rect 31205 19737 31217 19771
rect 31251 19768 31263 19771
rect 32030 19768 32036 19780
rect 31251 19740 32036 19768
rect 31251 19737 31263 19740
rect 31205 19731 31263 19737
rect 32030 19728 32036 19740
rect 32088 19768 32094 19780
rect 32508 19768 32536 19808
rect 32674 19805 32686 19808
rect 32720 19805 32732 19839
rect 32789 19839 32873 19845
rect 32789 19808 32827 19839
rect 32674 19799 32732 19805
rect 32815 19805 32827 19808
rect 32861 19805 32873 19839
rect 32815 19799 32873 19805
rect 33226 19796 33232 19848
rect 33284 19836 33290 19848
rect 33597 19839 33655 19845
rect 33597 19836 33609 19839
rect 33284 19808 33609 19836
rect 33284 19796 33290 19808
rect 33597 19805 33609 19808
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 34790 19796 34796 19848
rect 34848 19836 34854 19848
rect 34992 19845 35020 19944
rect 35066 19864 35072 19916
rect 35124 19904 35130 19916
rect 35124 19876 35388 19904
rect 35124 19864 35130 19876
rect 35360 19848 35388 19876
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 34848 19808 34897 19836
rect 34848 19796 34854 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 34978 19839 35036 19845
rect 34978 19805 34990 19839
rect 35024 19805 35036 19839
rect 34978 19799 35036 19805
rect 35250 19796 35256 19848
rect 35308 19796 35314 19848
rect 35342 19796 35348 19848
rect 35400 19845 35406 19848
rect 35400 19836 35408 19845
rect 35400 19808 35445 19836
rect 35400 19799 35408 19808
rect 35400 19796 35406 19799
rect 36722 19796 36728 19848
rect 36780 19796 36786 19848
rect 36992 19839 37050 19845
rect 36992 19805 37004 19839
rect 37038 19836 37050 19839
rect 37458 19836 37464 19848
rect 37038 19808 37464 19836
rect 37038 19805 37050 19808
rect 36992 19799 37050 19805
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 32088 19740 32536 19768
rect 32585 19771 32643 19777
rect 32088 19728 32094 19740
rect 32585 19737 32597 19771
rect 32631 19737 32643 19771
rect 32585 19731 32643 19737
rect 29512 19672 29592 19700
rect 29512 19660 29518 19672
rect 29914 19660 29920 19712
rect 29972 19700 29978 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 29972 19672 30113 19700
rect 29972 19660 29978 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 32600 19700 32628 19731
rect 35158 19728 35164 19780
rect 35216 19728 35222 19780
rect 32858 19700 32864 19712
rect 32600 19672 32864 19700
rect 30101 19663 30159 19669
rect 32858 19660 32864 19672
rect 32916 19660 32922 19712
rect 32950 19660 32956 19712
rect 33008 19660 33014 19712
rect 35268 19700 35296 19796
rect 37826 19700 37832 19712
rect 35268 19672 37832 19700
rect 37826 19660 37832 19672
rect 37884 19700 37890 19712
rect 38105 19703 38163 19709
rect 38105 19700 38117 19703
rect 37884 19672 38117 19700
rect 37884 19660 37890 19672
rect 38105 19669 38117 19672
rect 38151 19669 38163 19703
rect 38105 19663 38163 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 5626 19456 5632 19508
rect 5684 19456 5690 19508
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 7558 19496 7564 19508
rect 5767 19468 7564 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 9214 19496 9220 19508
rect 9171 19468 9220 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 9324 19468 10824 19496
rect 3688 19431 3746 19437
rect 3688 19397 3700 19431
rect 3734 19428 3746 19431
rect 4062 19428 4068 19440
rect 3734 19400 4068 19428
rect 3734 19397 3746 19400
rect 3688 19391 3746 19397
rect 4062 19388 4068 19400
rect 4120 19388 4126 19440
rect 7926 19388 7932 19440
rect 7984 19428 7990 19440
rect 9324 19428 9352 19468
rect 7984 19400 9352 19428
rect 9401 19431 9459 19437
rect 7984 19388 7990 19400
rect 3418 19320 3424 19372
rect 3476 19320 3482 19372
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 6638 19360 6644 19372
rect 4672 19332 6644 19360
rect 4672 19320 4678 19332
rect 5920 19301 5948 19332
rect 6638 19320 6644 19332
rect 6696 19360 6702 19372
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6696 19332 6837 19360
rect 6696 19320 6702 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 8478 19360 8484 19372
rect 7055 19332 8484 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19261 5963 19295
rect 9232 19292 9260 19400
rect 9401 19397 9413 19431
rect 9447 19428 9459 19431
rect 10502 19428 10508 19440
rect 9447 19400 10508 19428
rect 9447 19397 9459 19400
rect 9401 19391 9459 19397
rect 10502 19388 10508 19400
rect 10560 19388 10566 19440
rect 10796 19437 10824 19468
rect 10888 19468 13093 19496
rect 10888 19437 10916 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 13081 19459 13139 19465
rect 15105 19499 15163 19505
rect 15105 19465 15117 19499
rect 15151 19496 15163 19499
rect 15194 19496 15200 19508
rect 15151 19468 15200 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19397 10839 19431
rect 10781 19391 10839 19397
rect 10873 19431 10931 19437
rect 10873 19397 10885 19431
rect 10919 19397 10931 19431
rect 11946 19431 12004 19437
rect 11946 19428 11958 19431
rect 10873 19391 10931 19397
rect 11164 19400 11958 19428
rect 9306 19320 9312 19372
rect 9364 19320 9370 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9416 19332 9505 19360
rect 9416 19292 9444 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9674 19320 9680 19372
rect 9732 19320 9738 19372
rect 10594 19320 10600 19372
rect 10652 19320 10658 19372
rect 10962 19320 10968 19372
rect 11020 19320 11026 19372
rect 9232 19264 9444 19292
rect 5905 19255 5963 19261
rect 4430 19184 4436 19236
rect 4488 19224 4494 19236
rect 4801 19227 4859 19233
rect 4801 19224 4813 19227
rect 4488 19196 4813 19224
rect 4488 19184 4494 19196
rect 4801 19193 4813 19196
rect 4847 19224 4859 19227
rect 5442 19224 5448 19236
rect 4847 19196 5448 19224
rect 4847 19193 4859 19196
rect 4801 19187 4859 19193
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 11164 19233 11192 19400
rect 11946 19397 11958 19400
rect 11992 19397 12004 19431
rect 13096 19428 13124 19459
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 15562 19456 15568 19508
rect 15620 19456 15626 19508
rect 17494 19456 17500 19508
rect 17552 19496 17558 19508
rect 19242 19496 19248 19508
rect 17552 19468 19248 19496
rect 17552 19456 17558 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20162 19496 20168 19508
rect 20088 19468 20168 19496
rect 14645 19431 14703 19437
rect 14645 19428 14657 19431
rect 13096 19400 14657 19428
rect 11946 19391 12004 19397
rect 14645 19397 14657 19400
rect 14691 19397 14703 19431
rect 15470 19428 15476 19440
rect 14645 19391 14703 19397
rect 14844 19400 15476 19428
rect 14844 19372 14872 19400
rect 15470 19388 15476 19400
rect 15528 19388 15534 19440
rect 17512 19428 17540 19456
rect 18230 19428 18236 19440
rect 16592 19400 17540 19428
rect 17604 19400 18236 19428
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11572 19332 11713 19360
rect 11572 19320 11578 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 11149 19227 11207 19233
rect 11149 19193 11161 19227
rect 11195 19193 11207 19227
rect 11149 19187 11207 19193
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 14936 19224 14964 19323
rect 15930 19320 15936 19372
rect 15988 19320 15994 19372
rect 16592 19360 16620 19400
rect 16500 19332 16620 19360
rect 16022 19252 16028 19304
rect 16080 19252 16086 19304
rect 16209 19295 16267 19301
rect 16209 19261 16221 19295
rect 16255 19292 16267 19295
rect 16500 19292 16528 19332
rect 17310 19320 17316 19372
rect 17368 19320 17374 19372
rect 17402 19320 17408 19372
rect 17460 19320 17466 19372
rect 17604 19369 17632 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 17678 19320 17684 19372
rect 17736 19320 17742 19372
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19329 19487 19363
rect 20088 19360 20116 19468
rect 20162 19456 20168 19468
rect 20220 19496 20226 19508
rect 25133 19499 25191 19505
rect 20220 19468 23060 19496
rect 20220 19456 20226 19468
rect 21284 19437 21312 19468
rect 21269 19431 21327 19437
rect 21269 19397 21281 19431
rect 21315 19397 21327 19431
rect 21269 19391 21327 19397
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 23032 19428 23060 19468
rect 25133 19465 25145 19499
rect 25179 19496 25191 19499
rect 30926 19496 30932 19508
rect 25179 19468 30932 19496
rect 25179 19465 25191 19468
rect 25133 19459 25191 19465
rect 30926 19456 30932 19468
rect 30984 19456 30990 19508
rect 32670 19499 32728 19505
rect 32670 19465 32682 19499
rect 32716 19496 32728 19499
rect 33502 19496 33508 19508
rect 32716 19468 33508 19496
rect 32716 19465 32728 19468
rect 32670 19459 32728 19465
rect 33502 19456 33508 19468
rect 33560 19456 33566 19508
rect 35434 19456 35440 19508
rect 35492 19496 35498 19508
rect 35713 19499 35771 19505
rect 35713 19496 35725 19499
rect 35492 19468 35725 19496
rect 35492 19456 35498 19468
rect 35713 19465 35725 19468
rect 35759 19465 35771 19499
rect 35713 19459 35771 19465
rect 27062 19428 27068 19440
rect 21784 19400 22416 19428
rect 23032 19400 27068 19428
rect 21784 19388 21790 19400
rect 20158 19363 20216 19369
rect 20158 19360 20170 19363
rect 20088 19332 20170 19360
rect 19429 19323 19487 19329
rect 20158 19329 20170 19332
rect 20204 19329 20216 19363
rect 20158 19323 20216 19329
rect 17696 19292 17724 19320
rect 16255 19264 16528 19292
rect 17604 19264 17724 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 16224 19224 16252 19255
rect 17604 19224 17632 19264
rect 19058 19252 19064 19304
rect 19116 19252 19122 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19444 19292 19472 19323
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 20312 19332 20453 19360
rect 20312 19320 20318 19332
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20588 19332 20637 19360
rect 20588 19320 20594 19332
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 21174 19320 21180 19372
rect 21232 19360 21238 19372
rect 21453 19363 21511 19369
rect 21453 19360 21465 19363
rect 21232 19332 21465 19360
rect 21232 19320 21238 19332
rect 21453 19329 21465 19332
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 22278 19320 22284 19372
rect 22336 19320 22342 19372
rect 22388 19360 22416 19400
rect 27062 19388 27068 19400
rect 27120 19428 27126 19440
rect 27120 19400 27660 19428
rect 27120 19388 27126 19400
rect 22741 19363 22799 19369
rect 22741 19360 22753 19363
rect 22388 19332 22753 19360
rect 22741 19329 22753 19332
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 23014 19320 23020 19372
rect 23072 19320 23078 19372
rect 23106 19320 23112 19372
rect 23164 19320 23170 19372
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23348 19332 23397 19360
rect 23348 19320 23354 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 24578 19320 24584 19372
rect 24636 19320 24642 19372
rect 27154 19320 27160 19372
rect 27212 19320 27218 19372
rect 27632 19369 27660 19400
rect 28074 19388 28080 19440
rect 28132 19428 28138 19440
rect 28132 19400 28856 19428
rect 28132 19388 28138 19400
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 27982 19320 27988 19372
rect 28040 19360 28046 19372
rect 28828 19369 28856 19400
rect 29086 19388 29092 19440
rect 29144 19428 29150 19440
rect 29549 19431 29607 19437
rect 29549 19428 29561 19431
rect 29144 19400 29561 19428
rect 29144 19388 29150 19400
rect 29549 19397 29561 19400
rect 29595 19428 29607 19431
rect 30190 19428 30196 19440
rect 29595 19400 30196 19428
rect 29595 19397 29607 19400
rect 29549 19391 29607 19397
rect 30190 19388 30196 19400
rect 30248 19388 30254 19440
rect 31662 19388 31668 19440
rect 31720 19428 31726 19440
rect 32585 19431 32643 19437
rect 32585 19428 32597 19431
rect 31720 19400 32597 19428
rect 31720 19388 31726 19400
rect 32585 19397 32597 19400
rect 32631 19397 32643 19431
rect 32585 19391 32643 19397
rect 32769 19431 32827 19437
rect 32769 19397 32781 19431
rect 32815 19428 32827 19431
rect 32950 19428 32956 19440
rect 32815 19400 32956 19428
rect 32815 19397 32827 19400
rect 32769 19391 32827 19397
rect 32950 19388 32956 19400
rect 33008 19388 33014 19440
rect 33686 19388 33692 19440
rect 33744 19428 33750 19440
rect 36722 19428 36728 19440
rect 33744 19400 36728 19428
rect 33744 19388 33750 19400
rect 29454 19369 29460 19372
rect 28629 19363 28687 19369
rect 28629 19360 28641 19363
rect 28040 19332 28641 19360
rect 28040 19320 28046 19332
rect 28629 19329 28641 19332
rect 28675 19360 28687 19363
rect 28813 19363 28871 19369
rect 28675 19332 28764 19360
rect 28675 19329 28687 19332
rect 28629 19323 28687 19329
rect 19392 19264 19472 19292
rect 19392 19252 19398 19264
rect 20990 19252 20996 19304
rect 21048 19292 21054 19304
rect 21085 19295 21143 19301
rect 21085 19292 21097 19295
rect 21048 19264 21097 19292
rect 21048 19252 21054 19264
rect 21085 19261 21097 19264
rect 21131 19261 21143 19295
rect 21085 19255 21143 19261
rect 24857 19295 24915 19301
rect 24857 19261 24869 19295
rect 24903 19292 24915 19295
rect 25498 19292 25504 19304
rect 24903 19264 25504 19292
rect 24903 19261 24915 19264
rect 24857 19255 24915 19261
rect 25498 19252 25504 19264
rect 25556 19252 25562 19304
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 28350 19292 28356 19304
rect 27939 19264 28356 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 28350 19252 28356 19264
rect 28408 19292 28414 19304
rect 28534 19292 28540 19304
rect 28408 19264 28540 19292
rect 28408 19252 28414 19264
rect 28534 19252 28540 19264
rect 28592 19252 28598 19304
rect 24394 19224 24400 19236
rect 14884 19196 16252 19224
rect 16500 19196 17632 19224
rect 19306 19196 24400 19224
rect 14884 19184 14890 19196
rect 5258 19116 5264 19168
rect 5316 19116 5322 19168
rect 6730 19116 6736 19168
rect 6788 19156 6794 19168
rect 6917 19159 6975 19165
rect 6917 19156 6929 19159
rect 6788 19128 6929 19156
rect 6788 19116 6794 19128
rect 6917 19125 6929 19128
rect 6963 19125 6975 19159
rect 6917 19119 6975 19125
rect 14918 19116 14924 19168
rect 14976 19116 14982 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15378 19156 15384 19168
rect 15252 19128 15384 19156
rect 15252 19116 15258 19128
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16500 19156 16528 19196
rect 15896 19128 16528 19156
rect 15896 19116 15902 19128
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 17000 19128 17141 19156
rect 17000 19116 17006 19128
rect 17129 19125 17141 19128
rect 17175 19125 17187 19159
rect 17129 19119 17187 19125
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19306 19156 19334 19196
rect 24394 19184 24400 19196
rect 24452 19184 24458 19236
rect 24486 19184 24492 19236
rect 24544 19224 24550 19236
rect 27706 19224 27712 19236
rect 24544 19196 27712 19224
rect 24544 19184 24550 19196
rect 27706 19184 27712 19196
rect 27764 19184 27770 19236
rect 19116 19128 19334 19156
rect 19116 19116 19122 19128
rect 19978 19116 19984 19168
rect 20036 19116 20042 19168
rect 24762 19116 24768 19168
rect 24820 19116 24826 19168
rect 28736 19156 28764 19332
rect 28813 19329 28825 19363
rect 28859 19329 28871 19363
rect 29273 19363 29331 19369
rect 29273 19360 29285 19363
rect 28813 19323 28871 19329
rect 29104 19332 29285 19360
rect 29104 19304 29132 19332
rect 29273 19329 29285 19332
rect 29319 19329 29331 19363
rect 29273 19323 29331 19329
rect 29421 19363 29460 19369
rect 29421 19329 29433 19363
rect 29421 19323 29460 19329
rect 29454 19320 29460 19323
rect 29512 19320 29518 19372
rect 29638 19320 29644 19372
rect 29696 19320 29702 19372
rect 29730 19320 29736 19372
rect 29788 19369 29794 19372
rect 29788 19360 29796 19369
rect 32493 19363 32551 19369
rect 29788 19332 29833 19360
rect 29788 19323 29796 19332
rect 32493 19329 32505 19363
rect 32539 19360 32551 19363
rect 32674 19360 32680 19372
rect 32539 19332 32680 19360
rect 32539 19329 32551 19332
rect 32493 19323 32551 19329
rect 29788 19320 29794 19323
rect 32674 19320 32680 19332
rect 32732 19360 32738 19372
rect 33229 19363 33287 19369
rect 33229 19360 33241 19363
rect 32732 19332 33241 19360
rect 32732 19320 32738 19332
rect 33229 19329 33241 19332
rect 33275 19329 33287 19363
rect 33229 19323 33287 19329
rect 33318 19320 33324 19372
rect 33376 19320 33382 19372
rect 33502 19320 33508 19372
rect 33560 19320 33566 19372
rect 34348 19369 34376 19400
rect 36722 19388 36728 19400
rect 36780 19388 36786 19440
rect 34333 19363 34391 19369
rect 34333 19329 34345 19363
rect 34379 19329 34391 19363
rect 34333 19323 34391 19329
rect 34422 19320 34428 19372
rect 34480 19360 34486 19372
rect 34589 19363 34647 19369
rect 34589 19360 34601 19363
rect 34480 19332 34601 19360
rect 34480 19320 34486 19332
rect 34589 19329 34601 19332
rect 34635 19329 34647 19363
rect 34589 19323 34647 19329
rect 37550 19320 37556 19372
rect 37608 19360 37614 19372
rect 37829 19363 37887 19369
rect 37829 19360 37841 19363
rect 37608 19332 37841 19360
rect 37608 19320 37614 19332
rect 37829 19329 37841 19332
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 38105 19363 38163 19369
rect 38105 19329 38117 19363
rect 38151 19360 38163 19363
rect 39022 19360 39028 19372
rect 38151 19332 39028 19360
rect 38151 19329 38163 19332
rect 38105 19323 38163 19329
rect 39022 19320 39028 19332
rect 39080 19320 39086 19372
rect 29086 19252 29092 19304
rect 29144 19252 29150 19304
rect 31846 19252 31852 19304
rect 31904 19292 31910 19304
rect 31904 19264 34376 19292
rect 31904 19252 31910 19264
rect 28813 19227 28871 19233
rect 28813 19193 28825 19227
rect 28859 19224 28871 19227
rect 29822 19224 29828 19236
rect 28859 19196 29828 19224
rect 28859 19193 28871 19196
rect 28813 19187 28871 19193
rect 29822 19184 29828 19196
rect 29880 19184 29886 19236
rect 30098 19184 30104 19236
rect 30156 19224 30162 19236
rect 34146 19224 34152 19236
rect 30156 19196 34152 19224
rect 30156 19184 30162 19196
rect 34146 19184 34152 19196
rect 34204 19184 34210 19236
rect 29178 19156 29184 19168
rect 28736 19128 29184 19156
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 29270 19116 29276 19168
rect 29328 19156 29334 19168
rect 29917 19159 29975 19165
rect 29917 19156 29929 19159
rect 29328 19128 29929 19156
rect 29328 19116 29334 19128
rect 29917 19125 29929 19128
rect 29963 19125 29975 19159
rect 29917 19119 29975 19125
rect 33505 19159 33563 19165
rect 33505 19125 33517 19159
rect 33551 19156 33563 19159
rect 33594 19156 33600 19168
rect 33551 19128 33600 19156
rect 33551 19125 33563 19128
rect 33505 19119 33563 19125
rect 33594 19116 33600 19128
rect 33652 19116 33658 19168
rect 34348 19156 34376 19264
rect 35066 19156 35072 19168
rect 34348 19128 35072 19156
rect 35066 19116 35072 19128
rect 35124 19156 35130 19168
rect 35434 19156 35440 19168
rect 35124 19128 35440 19156
rect 35124 19116 35130 19128
rect 35434 19116 35440 19128
rect 35492 19116 35498 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 5626 18912 5632 18964
rect 5684 18952 5690 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 5684 18924 5825 18952
rect 5684 18912 5690 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 5813 18915 5871 18921
rect 13262 18912 13268 18964
rect 13320 18952 13326 18964
rect 15565 18955 15623 18961
rect 13320 18924 15516 18952
rect 13320 18912 13326 18924
rect 5442 18844 5448 18896
rect 5500 18884 5506 18896
rect 15488 18884 15516 18924
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 15930 18952 15936 18964
rect 15611 18924 15936 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 17126 18912 17132 18964
rect 17184 18952 17190 18964
rect 17773 18955 17831 18961
rect 17773 18952 17785 18955
rect 17184 18924 17785 18952
rect 17184 18912 17190 18924
rect 17773 18921 17785 18924
rect 17819 18921 17831 18955
rect 19886 18952 19892 18964
rect 17773 18915 17831 18921
rect 18064 18924 19892 18952
rect 18064 18884 18092 18924
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 20070 18952 20076 18964
rect 20027 18924 20076 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20070 18912 20076 18924
rect 20128 18952 20134 18964
rect 20530 18952 20536 18964
rect 20128 18924 20536 18952
rect 20128 18912 20134 18924
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 24578 18912 24584 18964
rect 24636 18912 24642 18964
rect 24765 18955 24823 18961
rect 24765 18921 24777 18955
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 5500 18856 15332 18884
rect 15488 18856 18092 18884
rect 18141 18887 18199 18893
rect 5500 18844 5506 18856
rect 6730 18776 6736 18828
rect 6788 18776 6794 18828
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 7101 18819 7159 18825
rect 7101 18816 7113 18819
rect 6972 18788 7113 18816
rect 6972 18776 6978 18788
rect 7101 18785 7113 18788
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 7374 18816 7380 18828
rect 7239 18788 7380 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 3476 18720 4445 18748
rect 3476 18708 3482 18720
rect 4433 18717 4445 18720
rect 4479 18748 4491 18751
rect 5626 18748 5632 18760
rect 4479 18720 5632 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6144 18720 6837 18748
rect 6144 18708 6150 18720
rect 6825 18717 6837 18720
rect 6871 18717 6883 18751
rect 7116 18748 7144 18779
rect 7374 18776 7380 18788
rect 7432 18816 7438 18828
rect 13354 18816 13360 18828
rect 7432 18788 13360 18816
rect 7432 18776 7438 18788
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 8662 18748 8668 18760
rect 7116 18720 8668 18748
rect 6825 18711 6883 18717
rect 8662 18708 8668 18720
rect 8720 18748 8726 18760
rect 9306 18748 9312 18760
rect 8720 18720 9312 18748
rect 8720 18708 8726 18720
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 13648 18748 13676 18779
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 15194 18748 15200 18760
rect 13648 18720 15200 18748
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 4700 18683 4758 18689
rect 4700 18649 4712 18683
rect 4746 18680 4758 18683
rect 5258 18680 5264 18692
rect 4746 18652 5264 18680
rect 4746 18649 4758 18652
rect 4700 18643 4758 18649
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 7208 18652 9260 18680
rect 6546 18572 6552 18624
rect 6604 18572 6610 18624
rect 6822 18572 6828 18624
rect 6880 18612 6886 18624
rect 7208 18612 7236 18652
rect 6880 18584 7236 18612
rect 6880 18572 6886 18584
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 8628 18584 9137 18612
rect 8628 18572 8634 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9232 18612 9260 18652
rect 9398 18640 9404 18692
rect 9456 18640 9462 18692
rect 9493 18683 9551 18689
rect 9493 18649 9505 18683
rect 9539 18680 9551 18683
rect 10318 18680 10324 18692
rect 9539 18652 10324 18680
rect 9539 18649 9551 18652
rect 9493 18643 9551 18649
rect 9508 18612 9536 18643
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 12437 18683 12495 18689
rect 12437 18649 12449 18683
rect 12483 18680 12495 18683
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 12483 18652 14657 18680
rect 12483 18649 12495 18652
rect 12437 18643 12495 18649
rect 14645 18649 14657 18652
rect 14691 18649 14703 18683
rect 15304 18680 15332 18856
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 19058 18884 19064 18896
rect 18187 18856 19064 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 19150 18844 19156 18896
rect 19208 18884 19214 18896
rect 19610 18884 19616 18896
rect 19208 18856 19616 18884
rect 19208 18844 19214 18856
rect 19610 18844 19616 18856
rect 19668 18844 19674 18896
rect 23290 18844 23296 18896
rect 23348 18884 23354 18896
rect 24780 18884 24808 18915
rect 32674 18912 32680 18964
rect 32732 18952 32738 18964
rect 33413 18955 33471 18961
rect 32732 18924 33364 18952
rect 32732 18912 32738 18924
rect 23348 18856 24808 18884
rect 33336 18884 33364 18924
rect 33413 18921 33425 18955
rect 33459 18952 33471 18955
rect 33502 18952 33508 18964
rect 33459 18924 33508 18952
rect 33459 18921 33471 18924
rect 33413 18915 33471 18921
rect 33502 18912 33508 18924
rect 33560 18912 33566 18964
rect 36078 18884 36084 18896
rect 33336 18856 36084 18884
rect 23348 18844 23354 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 17972 18788 19441 18816
rect 15470 18708 15476 18760
rect 15528 18708 15534 18760
rect 17972 18757 18000 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 30098 18816 30104 18828
rect 19429 18779 19487 18785
rect 26436 18788 30104 18816
rect 26436 18760 26464 18788
rect 30098 18776 30104 18788
rect 30156 18776 30162 18828
rect 31018 18776 31024 18828
rect 31076 18816 31082 18828
rect 31478 18816 31484 18828
rect 31076 18788 31484 18816
rect 31076 18776 31082 18788
rect 31478 18776 31484 18788
rect 31536 18816 31542 18828
rect 31536 18788 32076 18816
rect 31536 18776 31542 18788
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 16408 18720 17969 18748
rect 16408 18680 16436 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18322 18748 18328 18760
rect 18279 18720 18328 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 19797 18751 19855 18757
rect 19797 18748 19809 18751
rect 18432 18720 19809 18748
rect 15304 18652 16436 18680
rect 14645 18643 14703 18649
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 18432 18680 18460 18720
rect 19797 18717 19809 18720
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 19886 18708 19892 18760
rect 19944 18748 19950 18760
rect 20990 18748 20996 18760
rect 19944 18720 20996 18748
rect 19944 18708 19950 18720
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 22002 18748 22008 18760
rect 21499 18720 22008 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 24486 18748 24492 18760
rect 23624 18720 24492 18748
rect 23624 18708 23630 18720
rect 24486 18708 24492 18720
rect 24544 18748 24550 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24544 18720 24777 18748
rect 24544 18708 24550 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 16540 18652 18460 18680
rect 16540 18640 16546 18652
rect 18966 18640 18972 18692
rect 19024 18680 19030 18692
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 19024 18652 21373 18680
rect 19024 18640 19030 18652
rect 21361 18649 21373 18652
rect 21407 18649 21419 18683
rect 21361 18643 21419 18649
rect 24670 18640 24676 18692
rect 24728 18680 24734 18692
rect 24964 18680 24992 18711
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 26418 18708 26424 18760
rect 26476 18708 26482 18760
rect 26510 18708 26516 18760
rect 26568 18748 26574 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 26568 18720 28181 18748
rect 26568 18708 26574 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 24728 18652 24992 18680
rect 26329 18683 26387 18689
rect 24728 18640 24734 18652
rect 26329 18649 26341 18683
rect 26375 18680 26387 18683
rect 27246 18680 27252 18692
rect 26375 18652 27252 18680
rect 26375 18649 26387 18652
rect 26329 18643 26387 18649
rect 27246 18640 27252 18652
rect 27304 18640 27310 18692
rect 9232 18584 9536 18612
rect 9125 18575 9183 18581
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 12989 18615 13047 18621
rect 12989 18612 13001 18615
rect 12768 18584 13001 18612
rect 12768 18572 12774 18584
rect 12989 18581 13001 18584
rect 13035 18581 13047 18615
rect 12989 18575 13047 18581
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 13357 18615 13415 18621
rect 13357 18612 13369 18615
rect 13320 18584 13369 18612
rect 13320 18572 13326 18584
rect 13357 18581 13369 18584
rect 13403 18581 13415 18615
rect 13357 18575 13415 18581
rect 13449 18615 13507 18621
rect 13449 18581 13461 18615
rect 13495 18612 13507 18615
rect 14277 18615 14335 18621
rect 14277 18612 14289 18615
rect 13495 18584 14289 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 14277 18581 14289 18584
rect 14323 18581 14335 18615
rect 14277 18575 14335 18581
rect 14737 18615 14795 18621
rect 14737 18581 14749 18615
rect 14783 18612 14795 18615
rect 16758 18612 16764 18624
rect 14783 18584 16764 18612
rect 14783 18581 14795 18584
rect 14737 18575 14795 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 19613 18615 19671 18621
rect 19613 18581 19625 18615
rect 19659 18612 19671 18615
rect 20622 18612 20628 18624
rect 19659 18584 20628 18612
rect 19659 18581 19671 18584
rect 19613 18575 19671 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 26697 18615 26755 18621
rect 26697 18581 26709 18615
rect 26743 18612 26755 18615
rect 27890 18612 27896 18624
rect 26743 18584 27896 18612
rect 26743 18581 26755 18584
rect 26697 18575 26755 18581
rect 27890 18572 27896 18584
rect 27948 18572 27954 18624
rect 27982 18572 27988 18624
rect 28040 18572 28046 18624
rect 28184 18612 28212 18711
rect 28534 18708 28540 18760
rect 28592 18708 28598 18760
rect 30834 18708 30840 18760
rect 30892 18708 30898 18760
rect 31294 18708 31300 18760
rect 31352 18708 31358 18760
rect 31846 18708 31852 18760
rect 31904 18708 31910 18760
rect 32048 18757 32076 18788
rect 32490 18776 32496 18828
rect 32548 18816 32554 18828
rect 37737 18819 37795 18825
rect 32548 18788 33272 18816
rect 32548 18776 32554 18788
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 32272 18720 32781 18748
rect 32272 18708 32278 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 32917 18751 32975 18757
rect 32917 18717 32929 18751
rect 32963 18748 32975 18751
rect 32963 18717 32996 18748
rect 32917 18711 32996 18717
rect 28258 18640 28264 18692
rect 28316 18640 28322 18692
rect 28353 18683 28411 18689
rect 28353 18649 28365 18683
rect 28399 18680 28411 18683
rect 28718 18680 28724 18692
rect 28399 18652 28724 18680
rect 28399 18649 28411 18652
rect 28353 18643 28411 18649
rect 28718 18640 28724 18652
rect 28776 18680 28782 18692
rect 29730 18680 29736 18692
rect 28776 18652 29736 18680
rect 28776 18640 28782 18652
rect 29730 18640 29736 18652
rect 29788 18640 29794 18692
rect 32309 18683 32367 18689
rect 32309 18649 32321 18683
rect 32355 18680 32367 18683
rect 32674 18680 32680 18692
rect 32355 18652 32680 18680
rect 32355 18649 32367 18652
rect 32309 18643 32367 18649
rect 28994 18612 29000 18624
rect 28184 18584 29000 18612
rect 28994 18572 29000 18584
rect 29052 18572 29058 18624
rect 32214 18572 32220 18624
rect 32272 18612 32278 18624
rect 32324 18612 32352 18643
rect 32674 18640 32680 18652
rect 32732 18640 32738 18692
rect 32272 18584 32352 18612
rect 32968 18612 32996 18711
rect 33042 18708 33048 18760
rect 33100 18708 33106 18760
rect 33244 18757 33272 18788
rect 37737 18785 37749 18819
rect 37783 18816 37795 18819
rect 38010 18816 38016 18828
rect 37783 18788 38016 18816
rect 37783 18785 37795 18788
rect 37737 18779 37795 18785
rect 38010 18776 38016 18788
rect 38068 18776 38074 18828
rect 33234 18751 33292 18757
rect 33234 18717 33246 18751
rect 33280 18717 33292 18751
rect 35526 18748 35532 18760
rect 33234 18711 33292 18717
rect 33336 18720 35532 18748
rect 33134 18640 33140 18692
rect 33192 18680 33198 18692
rect 33336 18680 33364 18720
rect 35526 18708 35532 18720
rect 35584 18708 35590 18760
rect 37461 18683 37519 18689
rect 37461 18680 37473 18683
rect 33192 18652 33364 18680
rect 35360 18652 37473 18680
rect 33192 18640 33198 18652
rect 35360 18624 35388 18652
rect 37461 18649 37473 18652
rect 37507 18680 37519 18683
rect 38102 18680 38108 18692
rect 37507 18652 38108 18680
rect 37507 18649 37519 18652
rect 37461 18643 37519 18649
rect 38102 18640 38108 18652
rect 38160 18640 38166 18692
rect 35342 18612 35348 18624
rect 32968 18584 35348 18612
rect 32272 18572 32278 18584
rect 35342 18572 35348 18584
rect 35400 18572 35406 18624
rect 36998 18572 37004 18624
rect 37056 18612 37062 18624
rect 37093 18615 37151 18621
rect 37093 18612 37105 18615
rect 37056 18584 37105 18612
rect 37056 18572 37062 18584
rect 37093 18581 37105 18584
rect 37139 18581 37151 18615
rect 37093 18575 37151 18581
rect 37550 18572 37556 18624
rect 37608 18572 37614 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 10962 18408 10968 18420
rect 9364 18380 10968 18408
rect 9364 18368 9370 18380
rect 9122 18340 9128 18352
rect 8312 18312 9128 18340
rect 8312 18284 8340 18312
rect 9122 18300 9128 18312
rect 9180 18300 9186 18352
rect 10594 18340 10600 18352
rect 10152 18312 10600 18340
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 8570 18281 8576 18284
rect 8564 18272 8576 18281
rect 8531 18244 8576 18272
rect 8564 18235 8576 18244
rect 8570 18232 8576 18235
rect 8628 18232 8634 18284
rect 10152 18281 10180 18312
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10318 18232 10324 18284
rect 10376 18232 10382 18284
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 10704 18272 10732 18380
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 15838 18408 15844 18420
rect 13280 18380 15844 18408
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 12069 18343 12127 18349
rect 12069 18340 12081 18343
rect 11756 18312 12081 18340
rect 11756 18300 11762 18312
rect 12069 18309 12081 18312
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 10551 18244 10732 18272
rect 12345 18275 12403 18281
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 12345 18235 12403 18241
rect 12544 18244 13185 18272
rect 10428 18204 10456 18235
rect 10594 18204 10600 18216
rect 10428 18176 10600 18204
rect 10594 18164 10600 18176
rect 10652 18204 10658 18216
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 10652 18176 12173 18204
rect 10652 18164 10658 18176
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12360 18204 12388 18235
rect 12360 18176 12480 18204
rect 12161 18167 12219 18173
rect 9398 18096 9404 18148
rect 9456 18136 9462 18148
rect 9677 18139 9735 18145
rect 9677 18136 9689 18139
rect 9456 18108 9689 18136
rect 9456 18096 9462 18108
rect 9677 18105 9689 18108
rect 9723 18136 9735 18139
rect 9723 18108 12388 18136
rect 9723 18105 9735 18108
rect 9677 18099 9735 18105
rect 12360 18080 12388 18108
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 11238 18068 11244 18080
rect 10735 18040 11244 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 12342 18028 12348 18080
rect 12400 18028 12406 18080
rect 12452 18068 12480 18176
rect 12544 18145 12572 18244
rect 13173 18241 13185 18244
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 13280 18204 13308 18380
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 18966 18368 18972 18420
rect 19024 18368 19030 18420
rect 19061 18411 19119 18417
rect 19061 18377 19073 18411
rect 19107 18408 19119 18411
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19107 18380 19809 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 20180 18380 21036 18408
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 16206 18340 16212 18352
rect 13504 18312 16212 18340
rect 13504 18300 13510 18312
rect 16206 18300 16212 18312
rect 16264 18340 16270 18352
rect 16853 18343 16911 18349
rect 16853 18340 16865 18343
rect 16264 18312 16865 18340
rect 16264 18300 16270 18312
rect 16853 18309 16865 18312
rect 16899 18309 16911 18343
rect 20180 18340 20208 18380
rect 16853 18303 16911 18309
rect 19306 18312 20208 18340
rect 20257 18343 20315 18349
rect 13354 18232 13360 18284
rect 13412 18272 13418 18284
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 13412 18244 14749 18272
rect 13412 18232 13418 18244
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 13280 18176 13400 18204
rect 13372 18145 13400 18176
rect 13446 18164 13452 18216
rect 13504 18164 13510 18216
rect 14752 18204 14780 18235
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14884 18244 14933 18272
rect 14884 18232 14890 18244
rect 14921 18241 14933 18244
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 19306 18272 19334 18312
rect 20257 18309 20269 18343
rect 20303 18340 20315 18343
rect 20622 18340 20628 18352
rect 20303 18312 20628 18340
rect 20303 18309 20315 18312
rect 20257 18303 20315 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 21008 18349 21036 18380
rect 21266 18368 21272 18420
rect 21324 18408 21330 18420
rect 21453 18411 21511 18417
rect 21453 18408 21465 18411
rect 21324 18380 21465 18408
rect 21324 18368 21330 18380
rect 21453 18377 21465 18380
rect 21499 18377 21511 18411
rect 21453 18371 21511 18377
rect 22002 18368 22008 18420
rect 22060 18368 22066 18420
rect 24854 18368 24860 18420
rect 24912 18368 24918 18420
rect 28258 18368 28264 18420
rect 28316 18408 28322 18420
rect 28316 18380 29316 18408
rect 28316 18368 28322 18380
rect 20993 18343 21051 18349
rect 20993 18309 21005 18343
rect 21039 18340 21051 18343
rect 22830 18340 22836 18352
rect 21039 18312 22836 18340
rect 21039 18309 21051 18312
rect 20993 18303 21051 18309
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 23658 18340 23664 18352
rect 23400 18312 23664 18340
rect 16816 18244 19334 18272
rect 20165 18275 20223 18281
rect 16816 18232 16822 18244
rect 20165 18241 20177 18275
rect 20211 18272 20223 18275
rect 20438 18272 20444 18284
rect 20211 18244 20444 18272
rect 20211 18241 20223 18244
rect 20165 18235 20223 18241
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 21266 18232 21272 18284
rect 21324 18232 21330 18284
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22152 18244 22201 18272
rect 22152 18232 22158 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22370 18272 22376 18284
rect 22327 18244 22376 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18232 22526 18284
rect 23106 18232 23112 18284
rect 23164 18272 23170 18284
rect 23290 18272 23296 18284
rect 23164 18244 23296 18272
rect 23164 18232 23170 18244
rect 23290 18232 23296 18244
rect 23348 18232 23354 18284
rect 23400 18281 23428 18312
rect 23658 18300 23664 18312
rect 23716 18340 23722 18352
rect 24670 18340 24676 18352
rect 23716 18312 24676 18340
rect 23716 18300 23722 18312
rect 24670 18300 24676 18312
rect 24728 18300 24734 18352
rect 27890 18300 27896 18352
rect 27948 18340 27954 18352
rect 29288 18340 29316 18380
rect 29546 18368 29552 18420
rect 29604 18408 29610 18420
rect 29641 18411 29699 18417
rect 29641 18408 29653 18411
rect 29604 18380 29653 18408
rect 29604 18368 29610 18380
rect 29641 18377 29653 18380
rect 29687 18377 29699 18411
rect 29641 18371 29699 18377
rect 33226 18368 33232 18420
rect 33284 18368 33290 18420
rect 36633 18411 36691 18417
rect 36633 18377 36645 18411
rect 36679 18408 36691 18411
rect 37550 18408 37556 18420
rect 36679 18380 37556 18408
rect 36679 18377 36691 18380
rect 36633 18371 36691 18377
rect 37550 18368 37556 18380
rect 37608 18368 37614 18420
rect 27948 18312 29224 18340
rect 29288 18312 29776 18340
rect 27948 18300 27954 18312
rect 23385 18275 23443 18281
rect 23385 18241 23397 18275
rect 23431 18241 23443 18275
rect 23385 18235 23443 18241
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 23753 18275 23811 18281
rect 23753 18241 23765 18275
rect 23799 18272 23811 18275
rect 24581 18275 24639 18281
rect 24581 18272 24593 18275
rect 23799 18244 24593 18272
rect 23799 18241 23811 18244
rect 23753 18235 23811 18241
rect 24581 18241 24593 18244
rect 24627 18272 24639 18275
rect 24762 18272 24768 18284
rect 24627 18244 24768 18272
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 24762 18232 24768 18244
rect 24820 18272 24826 18284
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 24820 18244 25329 18272
rect 24820 18232 24826 18244
rect 25317 18241 25329 18244
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 17126 18204 17132 18216
rect 14752 18176 17132 18204
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 17586 18164 17592 18216
rect 17644 18164 17650 18216
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19978 18204 19984 18216
rect 19291 18176 19984 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20349 18207 20407 18213
rect 20349 18204 20361 18207
rect 20312 18176 20361 18204
rect 20312 18164 20318 18176
rect 20349 18173 20361 18176
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 21082 18164 21088 18216
rect 21140 18164 21146 18216
rect 23584 18204 23612 18232
rect 22664 18176 23612 18204
rect 12529 18139 12587 18145
rect 12529 18105 12541 18139
rect 12575 18105 12587 18139
rect 13357 18139 13415 18145
rect 12529 18099 12587 18105
rect 12636 18108 13124 18136
rect 12636 18068 12664 18108
rect 12452 18040 12664 18068
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 12989 18071 13047 18077
rect 12989 18068 13001 18071
rect 12952 18040 13001 18068
rect 12952 18028 12958 18040
rect 12989 18037 13001 18040
rect 13035 18037 13047 18071
rect 13096 18068 13124 18108
rect 13357 18105 13369 18139
rect 13403 18105 13415 18139
rect 14826 18136 14832 18148
rect 13357 18099 13415 18105
rect 13464 18108 14832 18136
rect 13464 18068 13492 18108
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 16022 18096 16028 18148
rect 16080 18136 16086 18148
rect 22664 18136 22692 18176
rect 24210 18164 24216 18216
rect 24268 18164 24274 18216
rect 24673 18207 24731 18213
rect 24673 18173 24685 18207
rect 24719 18204 24731 18207
rect 24854 18204 24860 18216
rect 24719 18176 24860 18204
rect 24719 18173 24731 18176
rect 24673 18167 24731 18173
rect 24854 18164 24860 18176
rect 24912 18204 24918 18216
rect 25516 18204 25544 18235
rect 25590 18232 25596 18284
rect 25648 18232 25654 18284
rect 28169 18275 28227 18281
rect 28169 18241 28181 18275
rect 28215 18272 28227 18275
rect 28902 18272 28908 18284
rect 28215 18244 28908 18272
rect 28215 18241 28227 18244
rect 28169 18235 28227 18241
rect 28902 18232 28908 18244
rect 28960 18232 28966 18284
rect 29196 18281 29224 18312
rect 29181 18275 29239 18281
rect 29181 18241 29193 18275
rect 29227 18241 29239 18275
rect 29643 18275 29701 18281
rect 29643 18272 29655 18275
rect 29181 18235 29239 18241
rect 29288 18244 29655 18272
rect 24912 18176 25544 18204
rect 24912 18164 24918 18176
rect 27798 18164 27804 18216
rect 27856 18204 27862 18216
rect 28077 18207 28135 18213
rect 28077 18204 28089 18207
rect 27856 18176 28089 18204
rect 27856 18164 27862 18176
rect 28077 18173 28089 18176
rect 28123 18173 28135 18207
rect 28077 18167 28135 18173
rect 28350 18164 28356 18216
rect 28408 18204 28414 18216
rect 29086 18204 29092 18216
rect 28408 18176 29092 18204
rect 28408 18164 28414 18176
rect 29086 18164 29092 18176
rect 29144 18204 29150 18216
rect 29288 18204 29316 18244
rect 29643 18241 29655 18244
rect 29689 18241 29701 18275
rect 29643 18235 29701 18241
rect 29144 18176 29316 18204
rect 29144 18164 29150 18176
rect 16080 18108 21128 18136
rect 16080 18096 16086 18108
rect 13096 18040 13492 18068
rect 12989 18031 13047 18037
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 14700 18040 14749 18068
rect 14700 18028 14706 18040
rect 14737 18037 14749 18040
rect 14783 18037 14795 18071
rect 14737 18031 14795 18037
rect 18598 18028 18604 18080
rect 18656 18028 18662 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20496 18040 21005 18068
rect 20496 18028 20502 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 21100 18068 21128 18108
rect 22388 18108 22692 18136
rect 21266 18068 21272 18080
rect 21100 18040 21272 18068
rect 20993 18031 21051 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 22388 18077 22416 18108
rect 22830 18096 22836 18148
rect 22888 18136 22894 18148
rect 28442 18136 28448 18148
rect 22888 18108 28448 18136
rect 22888 18096 22894 18108
rect 28442 18096 28448 18108
rect 28500 18096 28506 18148
rect 29270 18096 29276 18148
rect 29328 18096 29334 18148
rect 29748 18136 29776 18312
rect 33594 18300 33600 18352
rect 33652 18300 33658 18352
rect 35250 18300 35256 18352
rect 35308 18300 35314 18352
rect 35342 18300 35348 18352
rect 35400 18300 35406 18352
rect 33413 18275 33471 18281
rect 33413 18241 33425 18275
rect 33459 18272 33471 18275
rect 33502 18272 33508 18284
rect 33459 18244 33508 18272
rect 33459 18241 33471 18244
rect 33413 18235 33471 18241
rect 33502 18232 33508 18244
rect 33560 18232 33566 18284
rect 34790 18232 34796 18284
rect 34848 18272 34854 18284
rect 34977 18275 35035 18281
rect 34977 18272 34989 18275
rect 34848 18244 34989 18272
rect 34848 18232 34854 18244
rect 34977 18241 34989 18244
rect 35023 18241 35035 18275
rect 34977 18235 35035 18241
rect 34992 18204 35020 18235
rect 35066 18232 35072 18284
rect 35124 18232 35130 18284
rect 35434 18232 35440 18284
rect 35492 18281 35498 18284
rect 35492 18272 35500 18281
rect 35492 18244 35537 18272
rect 35492 18235 35500 18244
rect 35492 18232 35498 18235
rect 35894 18232 35900 18284
rect 35952 18272 35958 18284
rect 36081 18275 36139 18281
rect 36081 18272 36093 18275
rect 35952 18244 36093 18272
rect 35952 18232 35958 18244
rect 36081 18241 36093 18244
rect 36127 18241 36139 18275
rect 36081 18235 36139 18241
rect 36354 18232 36360 18284
rect 36412 18232 36418 18284
rect 36449 18275 36507 18281
rect 36449 18241 36461 18275
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 36464 18204 36492 18235
rect 37826 18232 37832 18284
rect 37884 18232 37890 18284
rect 34992 18176 35480 18204
rect 35452 18148 35480 18176
rect 35636 18176 36492 18204
rect 38105 18207 38163 18213
rect 29748 18108 31708 18136
rect 31680 18080 31708 18108
rect 35434 18096 35440 18148
rect 35492 18096 35498 18148
rect 35636 18145 35664 18176
rect 38105 18173 38117 18207
rect 38151 18204 38163 18207
rect 39022 18204 39028 18216
rect 38151 18176 39028 18204
rect 38151 18173 38163 18176
rect 38105 18167 38163 18173
rect 39022 18164 39028 18176
rect 39080 18164 39086 18216
rect 35621 18139 35679 18145
rect 35621 18105 35633 18139
rect 35667 18105 35679 18139
rect 35621 18099 35679 18105
rect 22373 18071 22431 18077
rect 22373 18037 22385 18071
rect 22419 18037 22431 18071
rect 22373 18031 22431 18037
rect 24578 18028 24584 18080
rect 24636 18068 24642 18080
rect 24946 18068 24952 18080
rect 24636 18040 24952 18068
rect 24636 18028 24642 18040
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25314 18028 25320 18080
rect 25372 18028 25378 18080
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 27801 18071 27859 18077
rect 27801 18068 27813 18071
rect 27672 18040 27813 18068
rect 27672 18028 27678 18040
rect 27801 18037 27813 18040
rect 27847 18037 27859 18071
rect 27801 18031 27859 18037
rect 29825 18071 29883 18077
rect 29825 18037 29837 18071
rect 29871 18068 29883 18071
rect 30190 18068 30196 18080
rect 29871 18040 30196 18068
rect 29871 18037 29883 18040
rect 29825 18031 29883 18037
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 31662 18028 31668 18080
rect 31720 18068 31726 18080
rect 33318 18068 33324 18080
rect 31720 18040 33324 18068
rect 31720 18028 31726 18040
rect 33318 18028 33324 18040
rect 33376 18028 33382 18080
rect 35802 18028 35808 18080
rect 35860 18068 35866 18080
rect 36173 18071 36231 18077
rect 36173 18068 36185 18071
rect 35860 18040 36185 18068
rect 35860 18028 35866 18040
rect 36173 18037 36185 18040
rect 36219 18037 36231 18071
rect 36173 18031 36231 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 7374 17824 7380 17876
rect 7432 17824 7438 17876
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 10594 17864 10600 17876
rect 10183 17836 10600 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 17126 17824 17132 17876
rect 17184 17824 17190 17876
rect 23109 17867 23167 17873
rect 17328 17836 22094 17864
rect 12250 17756 12256 17808
rect 12308 17796 12314 17808
rect 17037 17799 17095 17805
rect 17037 17796 17049 17799
rect 12308 17768 17049 17796
rect 12308 17756 12314 17768
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 5997 17663 6055 17669
rect 5997 17660 6009 17663
rect 5684 17632 6009 17660
rect 5684 17620 5690 17632
rect 5997 17629 6009 17632
rect 6043 17660 6055 17663
rect 8294 17660 8300 17672
rect 6043 17632 8300 17660
rect 6043 17629 6055 17632
rect 5997 17623 6055 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 11238 17620 11244 17672
rect 11296 17669 11302 17672
rect 11296 17660 11308 17669
rect 11296 17632 11341 17660
rect 11296 17623 11308 17632
rect 11296 17620 11302 17623
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 14384 17669 14412 17768
rect 17037 17765 17049 17768
rect 17083 17796 17095 17799
rect 17218 17796 17224 17808
rect 17083 17768 17224 17796
rect 17083 17765 17095 17768
rect 17037 17759 17095 17765
rect 17218 17756 17224 17768
rect 17276 17756 17282 17808
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 15703 17700 16681 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 17328 17728 17356 17836
rect 20070 17756 20076 17808
rect 20128 17796 20134 17808
rect 21545 17799 21603 17805
rect 21545 17796 21557 17799
rect 20128 17768 21557 17796
rect 20128 17756 20134 17768
rect 21545 17765 21557 17768
rect 21591 17765 21603 17799
rect 22066 17796 22094 17836
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 24210 17864 24216 17876
rect 23155 17836 24216 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 24210 17824 24216 17836
rect 24268 17824 24274 17876
rect 24302 17824 24308 17876
rect 24360 17864 24366 17876
rect 29089 17867 29147 17873
rect 24360 17836 27752 17864
rect 24360 17824 24366 17836
rect 22370 17796 22376 17808
rect 22066 17768 22376 17796
rect 21545 17759 21603 17765
rect 22370 17756 22376 17768
rect 22428 17796 22434 17808
rect 24228 17796 24256 17824
rect 25590 17796 25596 17808
rect 22428 17768 23244 17796
rect 24228 17768 25596 17796
rect 22428 17756 22434 17768
rect 16669 17691 16727 17697
rect 16868 17700 17356 17728
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17629 14427 17663
rect 14369 17623 14427 17629
rect 14462 17663 14520 17669
rect 14462 17629 14474 17663
rect 14508 17629 14520 17663
rect 14462 17623 14520 17629
rect 6264 17595 6322 17601
rect 6264 17561 6276 17595
rect 6310 17592 6322 17595
rect 6546 17592 6552 17604
rect 6310 17564 6552 17592
rect 6310 17561 6322 17564
rect 6264 17555 6322 17561
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 14476 17592 14504 17623
rect 14642 17620 14648 17672
rect 14700 17620 14706 17672
rect 14734 17620 14740 17672
rect 14792 17620 14798 17672
rect 14826 17620 14832 17672
rect 14884 17669 14890 17672
rect 14884 17663 14933 17669
rect 14884 17629 14887 17663
rect 14921 17660 14933 17663
rect 16868 17660 16896 17700
rect 18598 17688 18604 17740
rect 18656 17688 18662 17740
rect 18690 17688 18696 17740
rect 18748 17688 18754 17740
rect 23216 17728 23244 17768
rect 24029 17731 24087 17737
rect 18800 17700 22140 17728
rect 14921 17632 16896 17660
rect 14921 17629 14933 17632
rect 14884 17623 14933 17629
rect 14884 17620 14890 17623
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17218 17660 17224 17672
rect 17092 17632 17224 17660
rect 17092 17620 17098 17632
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17660 17463 17663
rect 17494 17660 17500 17672
rect 17451 17632 17500 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18800 17660 18828 17700
rect 17920 17632 18828 17660
rect 17920 17620 17926 17632
rect 21634 17620 21640 17672
rect 21692 17669 21698 17672
rect 22112 17669 22140 17700
rect 23216 17700 23888 17728
rect 21692 17663 21735 17669
rect 21723 17629 21735 17663
rect 21692 17623 21735 17629
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 22097 17663 22155 17669
rect 21867 17632 22048 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 21692 17620 21698 17623
rect 13872 17564 14504 17592
rect 15841 17595 15899 17601
rect 13872 17552 13878 17564
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 17126 17592 17132 17604
rect 15887 17564 17132 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 18104 17564 18521 17592
rect 18104 17552 18110 17564
rect 18509 17561 18521 17564
rect 18555 17592 18567 17595
rect 19242 17592 19248 17604
rect 18555 17564 19248 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 21910 17552 21916 17604
rect 21968 17552 21974 17604
rect 22020 17592 22048 17632
rect 22097 17629 22109 17663
rect 22143 17660 22155 17663
rect 23017 17663 23075 17669
rect 22143 17632 22876 17660
rect 22143 17629 22155 17632
rect 22097 17623 22155 17629
rect 22848 17592 22876 17632
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23106 17660 23112 17672
rect 23063 17632 23112 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 23216 17669 23244 17700
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17629 23259 17663
rect 23201 17623 23259 17629
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23860 17669 23888 17700
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24854 17728 24860 17740
rect 24075 17700 24860 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 24964 17737 24992 17768
rect 25590 17756 25596 17768
rect 25648 17756 25654 17808
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17697 25007 17731
rect 27724 17728 27752 17836
rect 29089 17833 29101 17867
rect 29135 17864 29147 17867
rect 32950 17864 32956 17876
rect 29135 17836 32956 17864
rect 29135 17833 29147 17836
rect 29089 17827 29147 17833
rect 32950 17824 32956 17836
rect 33008 17824 33014 17876
rect 38102 17824 38108 17876
rect 38160 17824 38166 17876
rect 31665 17799 31723 17805
rect 31665 17796 31677 17799
rect 31220 17768 31677 17796
rect 29454 17728 29460 17740
rect 27724 17700 29460 17728
rect 24949 17691 25007 17697
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 30653 17731 30711 17737
rect 30653 17697 30665 17731
rect 30699 17728 30711 17731
rect 31110 17728 31116 17740
rect 30699 17700 31116 17728
rect 30699 17697 30711 17700
rect 30653 17691 30711 17697
rect 31110 17688 31116 17700
rect 31168 17688 31174 17740
rect 31220 17737 31248 17768
rect 31665 17765 31677 17768
rect 31711 17765 31723 17799
rect 31665 17759 31723 17765
rect 31205 17731 31263 17737
rect 31205 17697 31217 17731
rect 31251 17697 31263 17731
rect 32490 17728 32496 17740
rect 31205 17691 31263 17697
rect 31864 17700 32496 17728
rect 31864 17672 31892 17700
rect 32490 17688 32496 17700
rect 32548 17688 32554 17740
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23348 17632 23673 17660
rect 23348 17620 23354 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 24302 17660 24308 17672
rect 23891 17632 24308 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 24302 17620 24308 17632
rect 24360 17620 24366 17672
rect 24578 17620 24584 17672
rect 24636 17660 24642 17672
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24636 17632 24685 17660
rect 24636 17620 24642 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 24762 17620 24768 17672
rect 24820 17620 24826 17672
rect 27453 17663 27511 17669
rect 27453 17629 27465 17663
rect 27499 17660 27511 17663
rect 27614 17660 27620 17672
rect 27499 17632 27620 17660
rect 27499 17629 27511 17632
rect 27453 17623 27511 17629
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 27706 17620 27712 17672
rect 27764 17620 27770 17672
rect 27798 17620 27804 17672
rect 27856 17660 27862 17672
rect 28721 17663 28779 17669
rect 28721 17660 28733 17663
rect 27856 17632 28733 17660
rect 27856 17620 27862 17632
rect 28721 17629 28733 17632
rect 28767 17629 28779 17663
rect 28721 17623 28779 17629
rect 30466 17620 30472 17672
rect 30524 17660 30530 17672
rect 30837 17663 30895 17669
rect 30837 17660 30849 17663
rect 30524 17632 30849 17660
rect 30524 17620 30530 17632
rect 30837 17629 30849 17632
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 31846 17620 31852 17672
rect 31904 17620 31910 17672
rect 32217 17663 32275 17669
rect 32217 17629 32229 17663
rect 32263 17660 32275 17663
rect 32582 17660 32588 17672
rect 32263 17632 32588 17660
rect 32263 17629 32275 17632
rect 32217 17623 32275 17629
rect 32582 17620 32588 17632
rect 32640 17620 32646 17672
rect 36722 17620 36728 17672
rect 36780 17620 36786 17672
rect 36998 17669 37004 17672
rect 36992 17660 37004 17669
rect 36959 17632 37004 17660
rect 36992 17623 37004 17632
rect 36998 17620 37004 17623
rect 37056 17620 37062 17672
rect 23750 17592 23756 17604
rect 22020 17564 22094 17592
rect 22848 17564 23756 17592
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 12621 17527 12679 17533
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 13078 17524 13084 17536
rect 12667 17496 13084 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 15010 17484 15016 17536
rect 15068 17484 15074 17536
rect 15746 17484 15752 17536
rect 15804 17484 15810 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 16172 17496 16221 17524
rect 16172 17484 16178 17496
rect 16209 17493 16221 17496
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 22066 17524 22094 17564
rect 23750 17552 23756 17564
rect 23808 17552 23814 17604
rect 26418 17592 26424 17604
rect 23952 17564 26424 17592
rect 23952 17524 23980 17564
rect 26418 17552 26424 17564
rect 26476 17552 26482 17604
rect 28902 17552 28908 17604
rect 28960 17552 28966 17604
rect 30742 17552 30748 17604
rect 30800 17592 30806 17604
rect 31941 17595 31999 17601
rect 31941 17592 31953 17595
rect 30800 17564 31953 17592
rect 30800 17552 30806 17564
rect 31941 17561 31953 17564
rect 31987 17561 31999 17595
rect 31941 17555 31999 17561
rect 32033 17595 32091 17601
rect 32033 17561 32045 17595
rect 32079 17592 32091 17595
rect 32306 17592 32312 17604
rect 32079 17564 32312 17592
rect 32079 17561 32091 17564
rect 32033 17555 32091 17561
rect 32306 17552 32312 17564
rect 32364 17592 32370 17604
rect 32858 17592 32864 17604
rect 32364 17564 32864 17592
rect 32364 17552 32370 17564
rect 32858 17552 32864 17564
rect 32916 17592 32922 17604
rect 33042 17592 33048 17604
rect 32916 17564 33048 17592
rect 32916 17552 32922 17564
rect 33042 17552 33048 17564
rect 33100 17552 33106 17604
rect 22066 17496 23980 17524
rect 25130 17484 25136 17536
rect 25188 17484 25194 17536
rect 26234 17484 26240 17536
rect 26292 17524 26298 17536
rect 26329 17527 26387 17533
rect 26329 17524 26341 17527
rect 26292 17496 26341 17524
rect 26292 17484 26298 17496
rect 26329 17493 26341 17496
rect 26375 17493 26387 17527
rect 28920 17524 28948 17552
rect 30837 17527 30895 17533
rect 30837 17524 30849 17527
rect 28920 17496 30849 17524
rect 26329 17487 26387 17493
rect 30837 17493 30849 17496
rect 30883 17493 30895 17527
rect 30837 17487 30895 17493
rect 30926 17484 30932 17536
rect 30984 17524 30990 17536
rect 34882 17524 34888 17536
rect 30984 17496 34888 17524
rect 30984 17484 30990 17496
rect 34882 17484 34888 17496
rect 34940 17484 34946 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12299 17292 12434 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 8481 17255 8539 17261
rect 8481 17252 8493 17255
rect 8444 17224 8493 17252
rect 8444 17212 8450 17224
rect 8481 17221 8493 17224
rect 8527 17221 8539 17255
rect 8481 17215 8539 17221
rect 8573 17255 8631 17261
rect 8573 17221 8585 17255
rect 8619 17252 8631 17255
rect 10502 17252 10508 17264
rect 8619 17224 10508 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 10502 17212 10508 17224
rect 10560 17212 10566 17264
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 11204 17224 11897 17252
rect 11204 17212 11210 17224
rect 11885 17221 11897 17224
rect 11931 17221 11943 17255
rect 11885 17215 11943 17221
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12406 17252 12434 17292
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 15804 17292 16037 17320
rect 15804 17280 15810 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 30285 17323 30343 17329
rect 16025 17283 16083 17289
rect 16132 17292 28764 17320
rect 12958 17255 13016 17261
rect 12958 17252 12970 17255
rect 12023 17224 12204 17252
rect 12406 17224 12970 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8312 17116 8340 17147
rect 8662 17144 8668 17196
rect 8720 17144 8726 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 8938 17116 8944 17128
rect 8312 17088 8944 17116
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 11716 17048 11744 17147
rect 12066 17144 12072 17196
rect 12124 17144 12130 17196
rect 12176 17184 12204 17224
rect 12958 17221 12970 17224
rect 13004 17221 13016 17255
rect 12958 17215 13016 17221
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 16132 17252 16160 17292
rect 19426 17252 19432 17264
rect 13136 17224 16160 17252
rect 17972 17224 19432 17252
rect 13136 17212 13142 17224
rect 12176 17156 14136 17184
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12400 17088 12725 17116
rect 12400 17076 12406 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 11716 17020 12434 17048
rect 8846 16940 8852 16992
rect 8904 16940 8910 16992
rect 12406 16980 12434 17020
rect 13078 16980 13084 16992
rect 12406 16952 13084 16980
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 14108 16989 14136 17156
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 15068 17156 15853 17184
rect 15068 17144 15074 17156
rect 15841 17153 15853 17156
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 17972 17193 18000 17224
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 18230 17193 18236 17196
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 15988 17156 17969 17184
rect 15988 17144 15994 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 18224 17184 18236 17193
rect 18191 17156 18236 17184
rect 17957 17147 18015 17153
rect 18224 17147 18236 17156
rect 18230 17144 18236 17147
rect 18288 17144 18294 17196
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 18984 17156 19993 17184
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17116 15623 17119
rect 17862 17116 17868 17128
rect 15611 17088 17868 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 17586 17048 17592 17060
rect 15712 17020 17592 17048
rect 15712 17008 15718 17020
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 16206 16980 16212 16992
rect 14139 16952 16212 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 17218 16940 17224 16992
rect 17276 16980 17282 16992
rect 18984 16980 19012 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 20272 17184 20300 17292
rect 22554 17212 22560 17264
rect 22612 17212 22618 17264
rect 22773 17255 22831 17261
rect 22773 17221 22785 17255
rect 22819 17252 22831 17255
rect 23290 17252 23296 17264
rect 22819 17224 23296 17252
rect 22819 17221 22831 17224
rect 22773 17215 22831 17221
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 23658 17212 23664 17264
rect 23716 17252 23722 17264
rect 23753 17255 23811 17261
rect 23753 17252 23765 17255
rect 23716 17224 23765 17252
rect 23716 17212 23722 17224
rect 23753 17221 23765 17224
rect 23799 17221 23811 17255
rect 23753 17215 23811 17221
rect 23842 17212 23848 17264
rect 23900 17252 23906 17264
rect 25222 17252 25228 17264
rect 23900 17224 25228 17252
rect 23900 17212 23906 17224
rect 20211 17156 20300 17184
rect 22572 17184 22600 17212
rect 23385 17187 23443 17193
rect 23385 17184 23397 17187
rect 22572 17156 23397 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 23385 17153 23397 17156
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 23584 17116 23612 17147
rect 24026 17144 24032 17196
rect 24084 17184 24090 17196
rect 24578 17184 24584 17196
rect 24084 17156 24584 17184
rect 24084 17144 24090 17156
rect 24578 17144 24584 17156
rect 24636 17144 24642 17196
rect 24688 17193 24716 17224
rect 25222 17212 25228 17224
rect 25280 17212 25286 17264
rect 28074 17212 28080 17264
rect 28132 17252 28138 17264
rect 28626 17252 28632 17264
rect 28132 17224 28632 17252
rect 28132 17212 28138 17224
rect 28626 17212 28632 17224
rect 28684 17212 28690 17264
rect 28736 17261 28764 17292
rect 30285 17289 30297 17323
rect 30331 17320 30343 17323
rect 30926 17320 30932 17332
rect 30331 17292 30932 17320
rect 30331 17289 30343 17292
rect 30285 17283 30343 17289
rect 30926 17280 30932 17292
rect 30984 17280 30990 17332
rect 31757 17323 31815 17329
rect 31036 17292 31524 17320
rect 28721 17255 28779 17261
rect 28721 17221 28733 17255
rect 28767 17221 28779 17255
rect 28721 17215 28779 17221
rect 29822 17212 29828 17264
rect 29880 17252 29886 17264
rect 30009 17255 30067 17261
rect 30009 17252 30021 17255
rect 29880 17224 30021 17252
rect 29880 17212 29886 17224
rect 30009 17221 30021 17224
rect 30055 17221 30067 17255
rect 30009 17215 30067 17221
rect 30374 17212 30380 17264
rect 30432 17252 30438 17264
rect 30650 17252 30656 17264
rect 30432 17224 30656 17252
rect 30432 17212 30438 17224
rect 30650 17212 30656 17224
rect 30708 17252 30714 17264
rect 31036 17252 31064 17292
rect 30708 17224 31064 17252
rect 30708 17212 30714 17224
rect 31110 17212 31116 17264
rect 31168 17252 31174 17264
rect 31496 17261 31524 17292
rect 31757 17289 31769 17323
rect 31803 17320 31815 17323
rect 33296 17323 33354 17329
rect 31803 17292 32904 17320
rect 31803 17289 31815 17292
rect 31757 17283 31815 17289
rect 31389 17255 31447 17261
rect 31389 17252 31401 17255
rect 31168 17224 31401 17252
rect 31168 17212 31174 17224
rect 31389 17221 31401 17224
rect 31435 17221 31447 17255
rect 31389 17215 31447 17221
rect 31481 17255 31539 17261
rect 31481 17221 31493 17255
rect 31527 17221 31539 17255
rect 31481 17215 31539 17221
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 25130 17144 25136 17196
rect 25188 17144 25194 17196
rect 25314 17144 25320 17196
rect 25372 17144 25378 17196
rect 27982 17144 27988 17196
rect 28040 17184 28046 17196
rect 28353 17187 28411 17193
rect 28353 17184 28365 17187
rect 28040 17156 28365 17184
rect 28040 17144 28046 17156
rect 28353 17153 28365 17156
rect 28399 17153 28411 17187
rect 28353 17147 28411 17153
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28818 17187 28876 17193
rect 28818 17184 28830 17187
rect 28500 17156 28545 17184
rect 28736 17156 28830 17184
rect 28500 17144 28506 17156
rect 23348 17088 23612 17116
rect 23348 17076 23354 17088
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 27246 17116 27252 17128
rect 26384 17088 27252 17116
rect 26384 17076 26390 17088
rect 27246 17076 27252 17088
rect 27304 17116 27310 17128
rect 28258 17116 28264 17128
rect 27304 17088 28264 17116
rect 27304 17076 27310 17088
rect 28258 17076 28264 17088
rect 28316 17116 28322 17128
rect 28736 17116 28764 17156
rect 28818 17153 28830 17156
rect 28864 17153 28876 17187
rect 28818 17147 28876 17153
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29638 17184 29644 17196
rect 29052 17156 29644 17184
rect 29052 17144 29058 17156
rect 29638 17144 29644 17156
rect 29696 17184 29702 17196
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 29696 17156 29745 17184
rect 29696 17144 29702 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17184 30159 17187
rect 30834 17184 30840 17196
rect 30147 17156 30840 17184
rect 30147 17153 30159 17156
rect 30101 17147 30159 17153
rect 28316 17088 28764 17116
rect 29932 17116 29960 17147
rect 30834 17144 30840 17156
rect 30892 17144 30898 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 30944 17156 31217 17184
rect 30374 17116 30380 17128
rect 29932 17088 30380 17116
rect 28316 17076 28322 17088
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 19300 17020 19349 17048
rect 19300 17008 19306 17020
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 19337 17011 19395 17017
rect 22925 17051 22983 17057
rect 22925 17017 22937 17051
rect 22971 17048 22983 17051
rect 23106 17048 23112 17060
rect 22971 17020 23112 17048
rect 22971 17017 22983 17020
rect 22925 17011 22983 17017
rect 23106 17008 23112 17020
rect 23164 17008 23170 17060
rect 28442 17008 28448 17060
rect 28500 17048 28506 17060
rect 30944 17048 30972 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 31573 17187 31631 17193
rect 31573 17153 31585 17187
rect 31619 17184 31631 17187
rect 31846 17184 31852 17196
rect 31619 17156 31852 17184
rect 31619 17153 31631 17156
rect 31573 17147 31631 17153
rect 31846 17144 31852 17156
rect 31904 17144 31910 17196
rect 32876 17193 32904 17292
rect 33296 17289 33308 17323
rect 33342 17320 33354 17323
rect 33686 17320 33692 17332
rect 33342 17292 33692 17320
rect 33342 17289 33354 17292
rect 33296 17283 33354 17289
rect 33686 17280 33692 17292
rect 33744 17280 33750 17332
rect 35161 17255 35219 17261
rect 35161 17221 35173 17255
rect 35207 17252 35219 17255
rect 37734 17252 37740 17264
rect 35207 17224 37740 17252
rect 35207 17221 35219 17224
rect 35161 17215 35219 17221
rect 37734 17212 37740 17224
rect 37792 17252 37798 17264
rect 37792 17224 37872 17252
rect 37792 17212 37798 17224
rect 32861 17187 32919 17193
rect 32861 17153 32873 17187
rect 32907 17153 32919 17187
rect 32861 17147 32919 17153
rect 33042 17144 33048 17196
rect 33100 17184 33106 17196
rect 33413 17187 33471 17193
rect 33413 17184 33425 17187
rect 33100 17156 33425 17184
rect 33100 17144 33106 17156
rect 33413 17153 33425 17156
rect 33459 17153 33471 17187
rect 33413 17147 33471 17153
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 34514 17184 34520 17196
rect 33735 17156 34520 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 34514 17144 34520 17156
rect 34572 17144 34578 17196
rect 34609 17187 34667 17193
rect 34609 17153 34621 17187
rect 34655 17184 34667 17187
rect 34698 17184 34704 17196
rect 34655 17156 34704 17184
rect 34655 17153 34667 17156
rect 34609 17147 34667 17153
rect 34698 17144 34704 17156
rect 34756 17144 34762 17196
rect 34882 17144 34888 17196
rect 34940 17144 34946 17196
rect 34977 17187 35035 17193
rect 34977 17153 34989 17187
rect 35023 17153 35035 17187
rect 34977 17147 35035 17153
rect 32122 17076 32128 17128
rect 32180 17116 32186 17128
rect 32180 17088 32798 17116
rect 32180 17076 32186 17088
rect 34790 17076 34796 17128
rect 34848 17116 34854 17128
rect 34992 17116 35020 17147
rect 35710 17144 35716 17196
rect 35768 17144 35774 17196
rect 35986 17144 35992 17196
rect 36044 17144 36050 17196
rect 36078 17144 36084 17196
rect 36136 17144 36142 17196
rect 37844 17193 37872 17224
rect 37829 17187 37887 17193
rect 37829 17153 37841 17187
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 34848 17088 35020 17116
rect 38105 17119 38163 17125
rect 34848 17076 34854 17088
rect 38105 17085 38117 17119
rect 38151 17116 38163 17119
rect 39022 17116 39028 17128
rect 38151 17088 39028 17116
rect 38151 17085 38163 17088
rect 38105 17079 38163 17085
rect 39022 17076 39028 17088
rect 39080 17076 39086 17128
rect 34701 17051 34759 17057
rect 28500 17020 34652 17048
rect 28500 17008 28506 17020
rect 17276 16952 19012 16980
rect 19797 16983 19855 16989
rect 17276 16940 17282 16952
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 19978 16980 19984 16992
rect 19843 16952 19984 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 19978 16940 19984 16952
rect 20036 16940 20042 16992
rect 22738 16940 22744 16992
rect 22796 16940 22802 16992
rect 25593 16983 25651 16989
rect 25593 16949 25605 16983
rect 25639 16980 25651 16983
rect 26142 16980 26148 16992
rect 25639 16952 26148 16980
rect 25639 16949 25651 16952
rect 25593 16943 25651 16949
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 28997 16983 29055 16989
rect 28997 16949 29009 16983
rect 29043 16980 29055 16983
rect 29454 16980 29460 16992
rect 29043 16952 29460 16980
rect 29043 16949 29055 16952
rect 28997 16943 29055 16949
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 34624 16980 34652 17020
rect 34701 17017 34713 17051
rect 34747 17048 34759 17051
rect 35802 17048 35808 17060
rect 34747 17020 35808 17048
rect 34747 17017 34759 17020
rect 34701 17011 34759 17017
rect 35802 17008 35808 17020
rect 35860 17008 35866 17060
rect 36265 17051 36323 17057
rect 36265 17017 36277 17051
rect 36311 17048 36323 17051
rect 37826 17048 37832 17060
rect 36311 17020 37832 17048
rect 36311 17017 36323 17020
rect 36265 17011 36323 17017
rect 37826 17008 37832 17020
rect 37884 17008 37890 17060
rect 35710 16980 35716 16992
rect 34624 16952 35716 16980
rect 35710 16940 35716 16952
rect 35768 16940 35774 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 9490 16776 9496 16788
rect 8812 16748 9496 16776
rect 8812 16736 8818 16748
rect 9490 16736 9496 16748
rect 9548 16776 9554 16788
rect 15654 16776 15660 16788
rect 9548 16748 15660 16776
rect 9548 16736 9554 16748
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 22738 16776 22744 16788
rect 16264 16748 22744 16776
rect 16264 16736 16270 16748
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 27522 16736 27528 16788
rect 27580 16776 27586 16788
rect 30466 16776 30472 16788
rect 27580 16748 30472 16776
rect 27580 16736 27586 16748
rect 30466 16736 30472 16748
rect 30524 16736 30530 16788
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 34885 16779 34943 16785
rect 34885 16776 34897 16779
rect 34848 16748 34897 16776
rect 34848 16736 34854 16748
rect 34885 16745 34897 16748
rect 34931 16745 34943 16779
rect 34885 16739 34943 16745
rect 12897 16711 12955 16717
rect 12897 16677 12909 16711
rect 12943 16708 12955 16711
rect 13078 16708 13084 16720
rect 12943 16680 13084 16708
rect 12943 16677 12955 16680
rect 12897 16671 12955 16677
rect 13078 16668 13084 16680
rect 13136 16668 13142 16720
rect 17126 16668 17132 16720
rect 17184 16708 17190 16720
rect 17221 16711 17279 16717
rect 17221 16708 17233 16711
rect 17184 16680 17233 16708
rect 17184 16668 17190 16680
rect 17221 16677 17233 16680
rect 17267 16708 17279 16711
rect 19150 16708 19156 16720
rect 17267 16680 19156 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 19150 16668 19156 16680
rect 19208 16668 19214 16720
rect 19242 16668 19248 16720
rect 19300 16708 19306 16720
rect 26697 16711 26755 16717
rect 19300 16680 26188 16708
rect 19300 16668 19306 16680
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 8294 16640 8300 16652
rect 7699 16612 8300 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 9122 16600 9128 16652
rect 9180 16600 9186 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9381 16575 9439 16581
rect 9381 16572 9393 16575
rect 8904 16544 9393 16572
rect 8904 16532 8910 16544
rect 9381 16541 9393 16544
rect 9427 16541 9439 16575
rect 9381 16535 9439 16541
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11532 16572 11560 16603
rect 15838 16600 15844 16652
rect 15896 16600 15902 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 19484 16612 21281 16640
rect 19484 16600 19490 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21634 16600 21640 16652
rect 21692 16640 21698 16652
rect 21692 16612 22140 16640
rect 21692 16600 21698 16612
rect 12342 16572 12348 16584
rect 11112 16544 12348 16572
rect 11112 16532 11118 16544
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 16114 16581 16120 16584
rect 16108 16572 16120 16581
rect 16075 16544 16120 16572
rect 16108 16535 16120 16544
rect 16114 16532 16120 16535
rect 16172 16532 16178 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 19306 16544 21465 16572
rect 5896 16507 5954 16513
rect 5896 16473 5908 16507
rect 5942 16504 5954 16507
rect 6546 16504 6552 16516
rect 5942 16476 6552 16504
rect 5942 16473 5954 16476
rect 5896 16467 5954 16473
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 8386 16464 8392 16516
rect 8444 16464 8450 16516
rect 11784 16507 11842 16513
rect 8496 16476 10640 16504
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16436 7067 16439
rect 8496 16436 8524 16476
rect 7055 16408 8524 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 10502 16396 10508 16448
rect 10560 16396 10566 16448
rect 10612 16436 10640 16476
rect 11784 16473 11796 16507
rect 11830 16504 11842 16507
rect 12250 16504 12256 16516
rect 11830 16476 12256 16504
rect 11830 16473 11842 16476
rect 11784 16467 11842 16473
rect 12250 16464 12256 16476
rect 12308 16464 12314 16516
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 19306 16504 19334 16544
rect 21453 16541 21465 16544
rect 21499 16572 21511 16575
rect 21542 16572 21548 16584
rect 21499 16544 21548 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 21542 16532 21548 16544
rect 21600 16532 21606 16584
rect 21910 16532 21916 16584
rect 21968 16532 21974 16584
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 22112 16572 22140 16612
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 23477 16643 23535 16649
rect 23477 16640 23489 16643
rect 23440 16612 23489 16640
rect 23440 16600 23446 16612
rect 23477 16609 23489 16612
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 22373 16575 22431 16581
rect 22373 16572 22385 16575
rect 22112 16544 22385 16572
rect 22005 16535 22063 16541
rect 22373 16541 22385 16544
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 15344 16476 19334 16504
rect 22020 16504 22048 16535
rect 22738 16532 22744 16584
rect 22796 16572 22802 16584
rect 26160 16581 26188 16680
rect 26697 16677 26709 16711
rect 26743 16708 26755 16711
rect 26743 16680 30144 16708
rect 26743 16677 26755 16680
rect 26697 16671 26755 16677
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 27522 16640 27528 16652
rect 26292 16612 27528 16640
rect 26292 16600 26298 16612
rect 23201 16575 23259 16581
rect 23201 16572 23213 16575
rect 22796 16544 23213 16572
rect 22796 16532 22802 16544
rect 23201 16541 23213 16544
rect 23247 16541 23259 16575
rect 23201 16535 23259 16541
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26326 16532 26332 16584
rect 26384 16532 26390 16584
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 27448 16581 27476 16612
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 28092 16612 28672 16640
rect 27341 16575 27399 16581
rect 27341 16572 27353 16575
rect 26568 16544 27353 16572
rect 26568 16532 26574 16544
rect 27341 16541 27353 16544
rect 27387 16541 27399 16575
rect 27341 16535 27399 16541
rect 27433 16575 27491 16581
rect 27433 16541 27445 16575
rect 27479 16541 27491 16575
rect 27433 16535 27491 16541
rect 22020 16476 22094 16504
rect 15344 16464 15350 16476
rect 12158 16436 12164 16448
rect 10612 16408 12164 16436
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 22066 16436 22094 16476
rect 23290 16464 23296 16516
rect 23348 16504 23354 16516
rect 23385 16507 23443 16513
rect 23385 16504 23397 16507
rect 23348 16476 23397 16504
rect 23348 16464 23354 16476
rect 23385 16473 23397 16476
rect 23431 16473 23443 16507
rect 26234 16504 26240 16516
rect 23385 16467 23443 16473
rect 23768 16476 26240 16504
rect 23768 16436 23796 16476
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 26418 16504 26424 16516
rect 26344 16476 26424 16504
rect 22066 16408 23796 16436
rect 23842 16396 23848 16448
rect 23900 16436 23906 16448
rect 26344 16436 26372 16476
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 27356 16504 27384 16535
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 27709 16575 27767 16581
rect 27709 16572 27721 16575
rect 27672 16544 27721 16572
rect 27672 16532 27678 16544
rect 27709 16541 27721 16544
rect 27755 16572 27767 16575
rect 28092 16572 28120 16612
rect 27755 16544 28120 16572
rect 27755 16541 27767 16544
rect 27709 16535 27767 16541
rect 28166 16532 28172 16584
rect 28224 16532 28230 16584
rect 28258 16532 28264 16584
rect 28316 16572 28322 16584
rect 28353 16575 28411 16581
rect 28353 16572 28365 16575
rect 28316 16544 28365 16572
rect 28316 16532 28322 16544
rect 28353 16541 28365 16544
rect 28399 16541 28411 16575
rect 28353 16535 28411 16541
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 27525 16507 27583 16513
rect 27356 16476 27476 16504
rect 23900 16408 26372 16436
rect 27157 16439 27215 16445
rect 23900 16396 23906 16408
rect 27157 16405 27169 16439
rect 27203 16436 27215 16439
rect 27338 16436 27344 16448
rect 27203 16408 27344 16436
rect 27203 16405 27215 16408
rect 27157 16399 27215 16405
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 27448 16436 27476 16476
rect 27525 16473 27537 16507
rect 27571 16504 27583 16507
rect 28074 16504 28080 16516
rect 27571 16476 28080 16504
rect 27571 16473 27583 16476
rect 27525 16467 27583 16473
rect 28074 16464 28080 16476
rect 28132 16464 28138 16516
rect 28442 16464 28448 16516
rect 28500 16464 28506 16516
rect 28552 16436 28580 16535
rect 28644 16504 28672 16612
rect 29270 16600 29276 16652
rect 29328 16640 29334 16652
rect 29822 16640 29828 16652
rect 29328 16612 29828 16640
rect 29328 16600 29334 16612
rect 29822 16600 29828 16612
rect 29880 16600 29886 16652
rect 29178 16532 29184 16584
rect 29236 16572 29242 16584
rect 29730 16572 29736 16584
rect 29236 16544 29736 16572
rect 29236 16532 29242 16544
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30006 16532 30012 16584
rect 30064 16532 30070 16584
rect 30116 16581 30144 16680
rect 33336 16680 33732 16708
rect 30282 16600 30288 16652
rect 30340 16600 30346 16652
rect 30374 16600 30380 16652
rect 30432 16640 30438 16652
rect 30432 16612 31340 16640
rect 30432 16600 30438 16612
rect 31312 16584 31340 16612
rect 32416 16612 32720 16640
rect 30101 16575 30159 16581
rect 30101 16541 30113 16575
rect 30147 16541 30159 16575
rect 30101 16535 30159 16541
rect 30926 16532 30932 16584
rect 30984 16532 30990 16584
rect 31018 16532 31024 16584
rect 31076 16572 31082 16584
rect 31113 16575 31171 16581
rect 31113 16572 31125 16575
rect 31076 16544 31125 16572
rect 31076 16532 31082 16544
rect 31113 16541 31125 16544
rect 31159 16541 31171 16575
rect 31113 16535 31171 16541
rect 31294 16532 31300 16584
rect 31352 16532 31358 16584
rect 31938 16532 31944 16584
rect 31996 16572 32002 16584
rect 32033 16575 32091 16581
rect 32033 16572 32045 16575
rect 31996 16544 32045 16572
rect 31996 16532 32002 16544
rect 32033 16541 32045 16544
rect 32079 16541 32091 16575
rect 32033 16535 32091 16541
rect 32181 16575 32239 16581
rect 32181 16541 32193 16575
rect 32227 16572 32239 16575
rect 32227 16541 32260 16572
rect 32181 16535 32260 16541
rect 30742 16504 30748 16516
rect 28644 16476 30748 16504
rect 30742 16464 30748 16476
rect 30800 16504 30806 16516
rect 31205 16507 31263 16513
rect 31205 16504 31217 16507
rect 30800 16476 31217 16504
rect 30800 16464 30806 16476
rect 31205 16473 31217 16476
rect 31251 16473 31263 16507
rect 31205 16467 31263 16473
rect 27448 16408 28580 16436
rect 28721 16439 28779 16445
rect 28721 16405 28733 16439
rect 28767 16436 28779 16439
rect 28994 16436 29000 16448
rect 28767 16408 29000 16436
rect 28767 16405 28779 16408
rect 28721 16399 28779 16405
rect 28994 16396 29000 16408
rect 29052 16396 29058 16448
rect 31481 16439 31539 16445
rect 31481 16405 31493 16439
rect 31527 16436 31539 16439
rect 32030 16436 32036 16448
rect 31527 16408 32036 16436
rect 31527 16405 31539 16408
rect 31481 16399 31539 16405
rect 32030 16396 32036 16408
rect 32088 16396 32094 16448
rect 32232 16436 32260 16535
rect 32306 16532 32312 16584
rect 32364 16532 32370 16584
rect 32416 16581 32444 16612
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 32490 16532 32496 16584
rect 32548 16581 32554 16584
rect 32548 16572 32556 16581
rect 32692 16572 32720 16612
rect 33336 16572 33364 16680
rect 33594 16600 33600 16652
rect 33652 16600 33658 16652
rect 32548 16544 32593 16572
rect 32692 16544 33364 16572
rect 32548 16535 32556 16544
rect 32548 16532 32554 16535
rect 33502 16532 33508 16584
rect 33560 16532 33566 16584
rect 33704 16572 33732 16680
rect 33870 16600 33876 16652
rect 33928 16600 33934 16652
rect 35268 16612 35664 16640
rect 34698 16572 34704 16584
rect 33704 16544 34704 16572
rect 34698 16532 34704 16544
rect 34756 16532 34762 16584
rect 35066 16581 35072 16584
rect 35064 16572 35072 16581
rect 35027 16544 35072 16572
rect 35064 16535 35072 16544
rect 35066 16532 35072 16535
rect 35124 16532 35130 16584
rect 35268 16572 35296 16612
rect 35381 16575 35439 16581
rect 35381 16572 35393 16575
rect 35176 16544 35296 16572
rect 35176 16513 35204 16544
rect 35360 16541 35393 16572
rect 35427 16541 35439 16575
rect 35360 16535 35439 16541
rect 35529 16575 35587 16581
rect 35529 16541 35541 16575
rect 35575 16541 35587 16575
rect 35636 16572 35664 16612
rect 36722 16600 36728 16652
rect 36780 16600 36786 16652
rect 37550 16572 37556 16584
rect 35636 16544 37556 16572
rect 35529 16535 35587 16541
rect 35161 16507 35219 16513
rect 35161 16504 35173 16507
rect 32600 16476 35173 16504
rect 32600 16436 32628 16476
rect 35161 16473 35173 16476
rect 35207 16473 35219 16507
rect 35161 16467 35219 16473
rect 35250 16464 35256 16516
rect 35308 16464 35314 16516
rect 32232 16408 32628 16436
rect 32677 16439 32735 16445
rect 32677 16405 32689 16439
rect 32723 16436 32735 16439
rect 33042 16436 33048 16448
rect 32723 16408 33048 16436
rect 32723 16405 32735 16408
rect 32677 16399 32735 16405
rect 33042 16396 33048 16408
rect 33100 16396 33106 16448
rect 34606 16396 34612 16448
rect 34664 16436 34670 16448
rect 35360 16436 35388 16535
rect 35544 16504 35572 16535
rect 37550 16532 37556 16544
rect 37608 16532 37614 16584
rect 35452 16476 35572 16504
rect 36992 16507 37050 16513
rect 35452 16448 35480 16476
rect 36992 16473 37004 16507
rect 37038 16504 37050 16507
rect 37458 16504 37464 16516
rect 37038 16476 37464 16504
rect 37038 16473 37050 16476
rect 36992 16467 37050 16473
rect 37458 16464 37464 16476
rect 37516 16464 37522 16516
rect 34664 16408 35388 16436
rect 34664 16396 34670 16408
rect 35434 16396 35440 16448
rect 35492 16396 35498 16448
rect 38102 16396 38108 16448
rect 38160 16396 38166 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 6546 16192 6552 16244
rect 6604 16192 6610 16244
rect 6914 16192 6920 16244
rect 6972 16192 6978 16244
rect 7006 16192 7012 16244
rect 7064 16192 7070 16244
rect 7926 16192 7932 16244
rect 7984 16192 7990 16244
rect 8938 16192 8944 16244
rect 8996 16192 9002 16244
rect 10686 16232 10692 16244
rect 9048 16204 10692 16232
rect 7024 16096 7052 16192
rect 7870 16099 7928 16105
rect 7870 16096 7882 16099
rect 7024 16068 7882 16096
rect 7870 16065 7882 16068
rect 7916 16065 7928 16099
rect 7870 16059 7928 16065
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8343 16068 8524 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6696 16000 7205 16028
rect 6696 15988 6702 16000
rect 7193 15997 7205 16000
rect 7239 16028 7251 16031
rect 8312 16028 8340 16059
rect 7239 16000 8340 16028
rect 8389 16031 8447 16037
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8496 16028 8524 16068
rect 8662 16056 8668 16108
rect 8720 16096 8726 16108
rect 9048 16105 9076 16204
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 21600 16204 23060 16232
rect 21600 16192 21606 16204
rect 11054 16164 11060 16176
rect 9784 16136 11060 16164
rect 9784 16105 9812 16136
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 15933 16167 15991 16173
rect 15933 16133 15945 16167
rect 15979 16164 15991 16167
rect 16022 16164 16028 16176
rect 15979 16136 16028 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 16022 16124 16028 16136
rect 16080 16124 16086 16176
rect 22554 16164 22560 16176
rect 19720 16136 22560 16164
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 8720 16068 8861 16096
rect 8720 16056 8726 16068
rect 8849 16065 8861 16068
rect 8895 16065 8907 16099
rect 8849 16059 8907 16065
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16065 9091 16099
rect 9033 16059 9091 16065
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 10036 16099 10094 16105
rect 10036 16065 10048 16099
rect 10082 16096 10094 16099
rect 10410 16096 10416 16108
rect 10082 16068 10416 16096
rect 10082 16065 10094 16068
rect 10036 16059 10094 16065
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 11514 16056 11520 16108
rect 11572 16096 11578 16108
rect 12986 16096 12992 16108
rect 11572 16068 12992 16096
rect 11572 16056 11578 16068
rect 12986 16056 12992 16068
rect 13044 16096 13050 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13044 16068 14289 16096
rect 13044 16056 13050 16068
rect 14277 16065 14289 16068
rect 14323 16096 14335 16099
rect 15838 16096 15844 16108
rect 14323 16068 15844 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 16908 16068 17233 16096
rect 16908 16056 16914 16068
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 9490 16028 9496 16040
rect 8496 16000 9496 16028
rect 8389 15991 8447 15997
rect 7742 15852 7748 15904
rect 7800 15852 7806 15904
rect 8404 15892 8432 15991
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 17328 16028 17356 16059
rect 17494 16056 17500 16108
rect 17552 16056 17558 16108
rect 19720 16105 19748 16136
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 22649 16167 22707 16173
rect 22649 16133 22661 16167
rect 22695 16164 22707 16167
rect 22738 16164 22744 16176
rect 22695 16136 22744 16164
rect 22695 16133 22707 16136
rect 22649 16127 22707 16133
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 22922 16173 22928 16176
rect 22865 16167 22928 16173
rect 22865 16133 22877 16167
rect 22911 16133 22928 16167
rect 22865 16127 22928 16133
rect 22922 16124 22928 16127
rect 22980 16124 22986 16176
rect 23032 16164 23060 16204
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 25682 16232 25688 16244
rect 23164 16204 25688 16232
rect 23164 16192 23170 16204
rect 25682 16192 25688 16204
rect 25740 16192 25746 16244
rect 31021 16235 31079 16241
rect 31021 16201 31033 16235
rect 31067 16201 31079 16235
rect 31021 16195 31079 16201
rect 24305 16167 24363 16173
rect 24305 16164 24317 16167
rect 23032 16136 24317 16164
rect 24305 16133 24317 16136
rect 24351 16164 24363 16167
rect 24394 16164 24400 16176
rect 24351 16136 24400 16164
rect 24351 16133 24363 16136
rect 24305 16127 24363 16133
rect 24394 16124 24400 16136
rect 24452 16124 24458 16176
rect 25958 16124 25964 16176
rect 26016 16124 26022 16176
rect 27614 16164 27620 16176
rect 27080 16136 27620 16164
rect 19978 16105 19984 16108
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16065 19763 16099
rect 19972 16096 19984 16105
rect 19939 16068 19984 16096
rect 19705 16059 19763 16065
rect 19972 16059 19984 16068
rect 19978 16056 19984 16059
rect 20036 16056 20042 16108
rect 21266 16056 21272 16108
rect 21324 16096 21330 16108
rect 21324 16068 24440 16096
rect 21324 16056 21330 16068
rect 17862 16028 17868 16040
rect 15580 16000 17868 16028
rect 10704 15932 12434 15960
rect 8478 15892 8484 15904
rect 8404 15864 8484 15892
rect 8478 15852 8484 15864
rect 8536 15892 8542 15904
rect 10704 15892 10732 15932
rect 8536 15864 10732 15892
rect 8536 15852 8542 15864
rect 11146 15852 11152 15904
rect 11204 15852 11210 15904
rect 12406 15892 12434 15932
rect 15580 15892 15608 16000
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 23014 16028 23020 16040
rect 22066 16000 23020 16028
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 22066 15960 22094 16000
rect 23014 15988 23020 16000
rect 23072 15988 23078 16040
rect 24412 16037 24440 16068
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25682 16096 25688 16108
rect 25096 16068 25688 16096
rect 25096 16056 25102 16068
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 27080 16096 27108 16136
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 30466 16124 30472 16176
rect 30524 16124 30530 16176
rect 25823 16068 27108 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 15997 24271 16031
rect 24213 15991 24271 15997
rect 24397 16031 24455 16037
rect 24397 15997 24409 16031
rect 24443 16028 24455 16031
rect 25792 16028 25820 16059
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 27212 16068 27261 16096
rect 27212 16056 27218 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27338 16056 27344 16108
rect 27396 16056 27402 16108
rect 27430 16056 27436 16108
rect 27488 16056 27494 16108
rect 27522 16056 27528 16108
rect 27580 16056 27586 16108
rect 28810 16056 28816 16108
rect 28868 16056 28874 16108
rect 28902 16056 28908 16108
rect 28960 16056 28966 16108
rect 28994 16056 29000 16108
rect 29052 16056 29058 16108
rect 29086 16056 29092 16108
rect 29144 16056 29150 16108
rect 30374 16056 30380 16108
rect 30432 16056 30438 16108
rect 30745 16099 30803 16105
rect 30745 16065 30757 16099
rect 30791 16096 30803 16099
rect 30926 16096 30932 16108
rect 30791 16068 30932 16096
rect 30791 16065 30803 16068
rect 30745 16059 30803 16065
rect 30926 16056 30932 16068
rect 30984 16056 30990 16108
rect 31036 16096 31064 16195
rect 31110 16192 31116 16244
rect 31168 16232 31174 16244
rect 32490 16232 32496 16244
rect 31168 16204 32496 16232
rect 31168 16192 31174 16204
rect 32490 16192 32496 16204
rect 32548 16192 32554 16244
rect 33502 16192 33508 16244
rect 33560 16192 33566 16244
rect 35066 16232 35072 16244
rect 34440 16204 35072 16232
rect 32030 16124 32036 16176
rect 32088 16164 32094 16176
rect 34440 16164 34468 16204
rect 35066 16192 35072 16204
rect 35124 16232 35130 16244
rect 35805 16235 35863 16241
rect 35124 16204 35664 16232
rect 35124 16192 35130 16204
rect 32088 16136 32444 16164
rect 32088 16124 32094 16136
rect 32416 16105 32444 16136
rect 32692 16136 34468 16164
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 31036 16068 32321 16096
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 32401 16099 32459 16105
rect 32401 16065 32413 16099
rect 32447 16065 32459 16099
rect 32401 16059 32459 16065
rect 32582 16056 32588 16108
rect 32640 16056 32646 16108
rect 32692 16105 32720 16136
rect 34514 16124 34520 16176
rect 34572 16164 34578 16176
rect 35529 16167 35587 16173
rect 35529 16164 35541 16167
rect 34572 16136 35541 16164
rect 34572 16124 34578 16136
rect 35529 16133 35541 16136
rect 35575 16133 35587 16167
rect 35529 16127 35587 16133
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 24443 16000 25820 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 23382 15960 23388 15972
rect 20772 15932 22094 15960
rect 22848 15932 23388 15960
rect 20772 15920 20778 15932
rect 12406 15864 15608 15892
rect 17678 15852 17684 15904
rect 17736 15852 17742 15904
rect 22848 15901 22876 15932
rect 23382 15920 23388 15932
rect 23440 15920 23446 15972
rect 24026 15920 24032 15972
rect 24084 15960 24090 15972
rect 24228 15960 24256 15991
rect 30834 15988 30840 16040
rect 30892 15988 30898 16040
rect 31754 15988 31760 16040
rect 31812 16028 31818 16040
rect 32692 16028 32720 16059
rect 33042 16056 33048 16108
rect 33100 16096 33106 16108
rect 33321 16099 33379 16105
rect 33321 16096 33333 16099
rect 33100 16068 33333 16096
rect 33100 16056 33106 16068
rect 33321 16065 33333 16068
rect 33367 16065 33379 16099
rect 33321 16059 33379 16065
rect 33686 16056 33692 16108
rect 33744 16056 33750 16108
rect 35161 16099 35219 16105
rect 35161 16065 35173 16099
rect 35207 16065 35219 16099
rect 35161 16059 35219 16065
rect 35254 16099 35312 16105
rect 35254 16065 35266 16099
rect 35300 16065 35312 16099
rect 35254 16059 35312 16065
rect 31812 16000 32720 16028
rect 31812 15988 31818 16000
rect 34974 15988 34980 16040
rect 35032 16028 35038 16040
rect 35167 16028 35195 16059
rect 35032 16000 35195 16028
rect 35268 16028 35296 16059
rect 35342 16056 35348 16108
rect 35400 16105 35406 16108
rect 35400 16099 35449 16105
rect 35400 16065 35403 16099
rect 35437 16065 35449 16099
rect 35400 16059 35449 16065
rect 35400 16056 35406 16059
rect 35544 16028 35572 16127
rect 35636 16105 35664 16204
rect 35805 16201 35817 16235
rect 35851 16232 35863 16235
rect 36078 16232 36084 16244
rect 35851 16204 36084 16232
rect 35851 16201 35863 16204
rect 35805 16195 35863 16201
rect 36078 16192 36084 16204
rect 36136 16192 36142 16244
rect 37458 16192 37464 16244
rect 37516 16192 37522 16244
rect 37826 16192 37832 16244
rect 37884 16232 37890 16244
rect 37921 16235 37979 16241
rect 37921 16232 37933 16235
rect 37884 16204 37933 16232
rect 37884 16192 37890 16204
rect 37921 16201 37933 16204
rect 37967 16201 37979 16235
rect 37921 16195 37979 16201
rect 35626 16099 35684 16105
rect 35626 16065 35638 16099
rect 35672 16065 35684 16099
rect 35626 16059 35684 16065
rect 37829 16099 37887 16105
rect 37829 16065 37841 16099
rect 37875 16096 37887 16099
rect 38102 16096 38108 16108
rect 37875 16068 38108 16096
rect 37875 16065 37887 16068
rect 37829 16059 37887 16065
rect 37844 16028 37872 16059
rect 38102 16056 38108 16068
rect 38160 16056 38166 16108
rect 35268 16000 35388 16028
rect 35544 16000 37872 16028
rect 35032 15988 35038 16000
rect 25038 15960 25044 15972
rect 24084 15932 25044 15960
rect 24084 15920 24090 15932
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15892 21143 15895
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 21131 15864 22845 15892
rect 21131 15861 21143 15864
rect 21085 15855 21143 15861
rect 22833 15861 22845 15864
rect 22879 15861 22891 15895
rect 22833 15855 22891 15861
rect 23017 15895 23075 15901
rect 23017 15861 23029 15895
rect 23063 15892 23075 15895
rect 24394 15892 24400 15904
rect 23063 15864 24400 15892
rect 23063 15861 23075 15864
rect 23017 15855 23075 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 24765 15895 24823 15901
rect 24765 15861 24777 15895
rect 24811 15892 24823 15895
rect 25222 15892 25228 15904
rect 24811 15864 25228 15892
rect 24811 15861 24823 15864
rect 24765 15855 24823 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 25958 15852 25964 15904
rect 26016 15852 26022 15904
rect 27709 15895 27767 15901
rect 27709 15861 27721 15895
rect 27755 15892 27767 15895
rect 28074 15892 28080 15904
rect 27755 15864 28080 15892
rect 27755 15861 27767 15864
rect 27709 15855 27767 15861
rect 28074 15852 28080 15864
rect 28132 15852 28138 15904
rect 29273 15895 29331 15901
rect 29273 15861 29285 15895
rect 29319 15892 29331 15895
rect 29546 15892 29552 15904
rect 29319 15864 29552 15892
rect 29319 15861 29331 15864
rect 29273 15855 29331 15861
rect 29546 15852 29552 15864
rect 29604 15852 29610 15904
rect 31478 15852 31484 15904
rect 31536 15892 31542 15904
rect 32858 15892 32864 15904
rect 31536 15864 32864 15892
rect 31536 15852 31542 15864
rect 32858 15852 32864 15864
rect 32916 15852 32922 15904
rect 32950 15852 32956 15904
rect 33008 15892 33014 15904
rect 33689 15895 33747 15901
rect 33689 15892 33701 15895
rect 33008 15864 33701 15892
rect 33008 15852 33014 15864
rect 33689 15861 33701 15864
rect 33735 15861 33747 15895
rect 33689 15855 33747 15861
rect 33778 15852 33784 15904
rect 33836 15892 33842 15904
rect 35360 15892 35388 16000
rect 38010 15988 38016 16040
rect 38068 15988 38074 16040
rect 33836 15864 35388 15892
rect 33836 15852 33842 15864
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 6457 15691 6515 15697
rect 6457 15657 6469 15691
rect 6503 15688 6515 15691
rect 8478 15688 8484 15700
rect 6503 15660 8484 15688
rect 6503 15657 6515 15660
rect 6457 15651 6515 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 10410 15648 10416 15700
rect 10468 15648 10474 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 13446 15688 13452 15700
rect 10827 15660 13452 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 27154 15648 27160 15700
rect 27212 15648 27218 15700
rect 28810 15648 28816 15700
rect 28868 15688 28874 15700
rect 29089 15691 29147 15697
rect 29089 15688 29101 15691
rect 28868 15660 29101 15688
rect 28868 15648 28874 15660
rect 29089 15657 29101 15660
rect 29135 15657 29147 15691
rect 34698 15688 34704 15700
rect 29089 15651 29147 15657
rect 29196 15660 34704 15688
rect 11698 15580 11704 15632
rect 11756 15620 11762 15632
rect 11793 15623 11851 15629
rect 11793 15620 11805 15623
rect 11756 15592 11805 15620
rect 11756 15580 11762 15592
rect 11793 15589 11805 15592
rect 11839 15589 11851 15623
rect 16853 15623 16911 15629
rect 11793 15583 11851 15589
rect 12406 15592 16252 15620
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11146 15552 11152 15564
rect 10919 15524 11152 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 11146 15512 11152 15524
rect 11204 15552 11210 15564
rect 12406 15552 12434 15592
rect 11204 15524 12434 15552
rect 11204 15512 11210 15524
rect 12986 15512 12992 15564
rect 13044 15512 13050 15564
rect 7581 15487 7639 15493
rect 7581 15453 7593 15487
rect 7627 15484 7639 15487
rect 7742 15484 7748 15496
rect 7627 15456 7748 15484
rect 7627 15453 7639 15456
rect 7581 15447 7639 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7834 15444 7840 15496
rect 7892 15444 7898 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10284 15456 10609 15484
rect 10284 15444 10290 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 11790 15444 11796 15496
rect 11848 15444 11854 15496
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 11992 15456 13737 15484
rect 11992 15428 12020 15456
rect 13725 15453 13737 15456
rect 13771 15484 13783 15487
rect 14274 15484 14280 15496
rect 13771 15456 14280 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 16224 15493 16252 15592
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 18414 15620 18420 15632
rect 16899 15592 18420 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 18414 15580 18420 15592
rect 18472 15580 18478 15632
rect 18506 15580 18512 15632
rect 18564 15580 18570 15632
rect 20254 15580 20260 15632
rect 20312 15620 20318 15632
rect 21453 15623 21511 15629
rect 21453 15620 21465 15623
rect 20312 15592 21465 15620
rect 20312 15580 20318 15592
rect 21453 15589 21465 15592
rect 21499 15589 21511 15623
rect 21453 15583 21511 15589
rect 26418 15580 26424 15632
rect 26476 15620 26482 15632
rect 29196 15620 29224 15660
rect 34698 15648 34704 15660
rect 34756 15648 34762 15700
rect 35621 15691 35679 15697
rect 35621 15657 35633 15691
rect 35667 15688 35679 15691
rect 35986 15688 35992 15700
rect 35667 15660 35992 15688
rect 35667 15657 35679 15660
rect 35621 15651 35679 15657
rect 35986 15648 35992 15660
rect 36044 15648 36050 15700
rect 30834 15620 30840 15632
rect 26476 15592 29224 15620
rect 29288 15592 30840 15620
rect 26476 15580 26482 15592
rect 17589 15555 17647 15561
rect 17589 15552 17601 15555
rect 16868 15524 17601 15552
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 8386 15376 8392 15428
rect 8444 15416 8450 15428
rect 11974 15416 11980 15428
rect 8444 15388 11980 15416
rect 8444 15376 8450 15388
rect 11974 15376 11980 15388
rect 12032 15376 12038 15428
rect 16132 15416 16160 15447
rect 16868 15428 16896 15524
rect 17589 15521 17601 15524
rect 17635 15552 17647 15555
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 17635 15524 19625 15552
rect 17635 15521 17647 15524
rect 17589 15515 17647 15521
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 29288 15552 29316 15592
rect 30834 15580 30840 15592
rect 30892 15580 30898 15632
rect 38010 15620 38016 15632
rect 31680 15592 38016 15620
rect 19613 15515 19671 15521
rect 27080 15524 29316 15552
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 16850 15416 16856 15428
rect 12084 15388 16856 15416
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 12084 15348 12112 15388
rect 16850 15376 16856 15388
rect 16908 15376 16914 15428
rect 16960 15416 16988 15447
rect 17862 15444 17868 15496
rect 17920 15444 17926 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18647 15456 19441 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15484 19763 15487
rect 20346 15484 20352 15496
rect 19751 15456 20352 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 17494 15416 17500 15428
rect 16960 15388 17500 15416
rect 17494 15376 17500 15388
rect 17552 15416 17558 15428
rect 18616 15416 18644 15447
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 20530 15444 20536 15496
rect 20588 15444 20594 15496
rect 21634 15493 21640 15496
rect 21632 15484 21640 15493
rect 21595 15456 21640 15484
rect 21632 15447 21640 15456
rect 21634 15444 21640 15447
rect 21692 15444 21698 15496
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15484 21787 15487
rect 21775 15456 21956 15484
rect 21775 15453 21787 15456
rect 21729 15447 21787 15453
rect 17552 15388 18644 15416
rect 17552 15376 17558 15388
rect 21818 15376 21824 15428
rect 21876 15376 21882 15428
rect 21928 15416 21956 15456
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22980 15456 23029 15484
rect 22980 15444 22986 15456
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 23290 15444 23296 15496
rect 23348 15444 23354 15496
rect 24854 15444 24860 15496
rect 24912 15444 24918 15496
rect 25038 15444 25044 15496
rect 25096 15444 25102 15496
rect 25866 15444 25872 15496
rect 25924 15484 25930 15496
rect 27080 15493 27108 15524
rect 30374 15512 30380 15564
rect 30432 15512 30438 15564
rect 31478 15512 31484 15564
rect 31536 15512 31542 15564
rect 31680 15561 31708 15592
rect 31665 15555 31723 15561
rect 31665 15521 31677 15555
rect 31711 15521 31723 15555
rect 31665 15515 31723 15521
rect 35434 15512 35440 15564
rect 35492 15512 35498 15564
rect 37734 15512 37740 15564
rect 37792 15552 37798 15564
rect 37936 15561 37964 15592
rect 38010 15580 38016 15592
rect 38068 15580 38074 15632
rect 37829 15555 37887 15561
rect 37829 15552 37841 15555
rect 37792 15524 37841 15552
rect 37792 15512 37798 15524
rect 37829 15521 37841 15524
rect 37875 15521 37887 15555
rect 37829 15515 37887 15521
rect 37921 15555 37979 15561
rect 37921 15521 37933 15555
rect 37967 15521 37979 15555
rect 37921 15515 37979 15521
rect 27065 15487 27123 15493
rect 27065 15484 27077 15487
rect 25924 15456 27077 15484
rect 25924 15444 25930 15456
rect 27065 15453 27077 15456
rect 27111 15453 27123 15487
rect 27065 15447 27123 15453
rect 27249 15487 27307 15493
rect 27249 15453 27261 15487
rect 27295 15484 27307 15487
rect 27522 15484 27528 15496
rect 27295 15456 27528 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 27522 15444 27528 15456
rect 27580 15484 27586 15496
rect 28997 15487 29055 15493
rect 28997 15484 29009 15487
rect 27580 15456 29009 15484
rect 27580 15444 27586 15456
rect 28997 15453 29009 15456
rect 29043 15484 29055 15487
rect 29086 15484 29092 15496
rect 29043 15456 29092 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 29178 15444 29184 15496
rect 29236 15444 29242 15496
rect 30561 15487 30619 15493
rect 30561 15453 30573 15487
rect 30607 15484 30619 15487
rect 32214 15484 32220 15496
rect 30607 15456 32220 15484
rect 30607 15453 30619 15456
rect 30561 15447 30619 15453
rect 32214 15444 32220 15456
rect 32272 15444 32278 15496
rect 35342 15444 35348 15496
rect 35400 15444 35406 15496
rect 23385 15419 23443 15425
rect 21928 15388 22094 15416
rect 11848 15320 12112 15348
rect 11848 15308 11854 15320
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 20714 15348 20720 15360
rect 12216 15320 20720 15348
rect 12216 15308 12222 15320
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 22066 15348 22094 15388
rect 23385 15385 23397 15419
rect 23431 15416 23443 15419
rect 24486 15416 24492 15428
rect 23431 15388 24492 15416
rect 23431 15385 23443 15388
rect 23385 15379 23443 15385
rect 24486 15376 24492 15388
rect 24544 15376 24550 15428
rect 28442 15416 28448 15428
rect 24872 15388 28448 15416
rect 24872 15348 24900 15388
rect 28442 15376 28448 15388
rect 28500 15376 28506 15428
rect 31389 15419 31447 15425
rect 31389 15385 31401 15419
rect 31435 15416 31447 15419
rect 31435 15388 31754 15416
rect 31435 15385 31447 15388
rect 31389 15379 31447 15385
rect 31726 15360 31754 15388
rect 34974 15376 34980 15428
rect 35032 15376 35038 15428
rect 35066 15376 35072 15428
rect 35124 15376 35130 15428
rect 37550 15376 37556 15428
rect 37608 15416 37614 15428
rect 37737 15419 37795 15425
rect 37737 15416 37749 15419
rect 37608 15388 37749 15416
rect 37608 15376 37614 15388
rect 37737 15385 37749 15388
rect 37783 15385 37795 15419
rect 37737 15379 37795 15385
rect 22066 15320 24900 15348
rect 24949 15351 25007 15357
rect 24949 15317 24961 15351
rect 24995 15348 25007 15351
rect 25406 15348 25412 15360
rect 24995 15320 25412 15348
rect 24995 15317 25007 15320
rect 24949 15311 25007 15317
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 31018 15308 31024 15360
rect 31076 15308 31082 15360
rect 31726 15320 31760 15360
rect 31754 15308 31760 15320
rect 31812 15348 31818 15360
rect 32582 15348 32588 15360
rect 31812 15320 32588 15348
rect 31812 15308 31818 15320
rect 32582 15308 32588 15320
rect 32640 15308 32646 15360
rect 32858 15308 32864 15360
rect 32916 15348 32922 15360
rect 35710 15348 35716 15360
rect 32916 15320 35716 15348
rect 32916 15308 32922 15320
rect 35710 15308 35716 15320
rect 35768 15308 35774 15360
rect 37182 15308 37188 15360
rect 37240 15348 37246 15360
rect 37369 15351 37427 15357
rect 37369 15348 37381 15351
rect 37240 15320 37381 15348
rect 37240 15308 37246 15320
rect 37369 15317 37381 15320
rect 37415 15317 37427 15351
rect 37369 15311 37427 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9916 15116 9965 15144
rect 9916 15104 9922 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 14550 15144 14556 15156
rect 13955 15116 14556 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 22080 15147 22138 15153
rect 22080 15144 22092 15147
rect 18104 15116 22092 15144
rect 18104 15104 18110 15116
rect 22080 15113 22092 15116
rect 22126 15113 22138 15147
rect 23842 15144 23848 15156
rect 22080 15107 22138 15113
rect 22572 15116 23848 15144
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 8941 15079 8999 15085
rect 8941 15076 8953 15079
rect 7892 15048 8953 15076
rect 7892 15036 7898 15048
rect 8941 15045 8953 15048
rect 8987 15076 8999 15079
rect 9122 15076 9128 15088
rect 8987 15048 9128 15076
rect 8987 15045 8999 15048
rect 8941 15039 8999 15045
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 11974 15036 11980 15088
rect 12032 15036 12038 15088
rect 15286 15036 15292 15088
rect 15344 15076 15350 15088
rect 16482 15076 16488 15088
rect 15344 15048 16488 15076
rect 15344 15036 15350 15048
rect 16482 15036 16488 15048
rect 16540 15076 16546 15088
rect 16540 15048 17540 15076
rect 16540 15036 16546 15048
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8386 15008 8392 15020
rect 8159 14980 8392 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 9858 14968 9864 15020
rect 9916 14968 9922 15020
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13320 14980 13553 15008
rect 13320 14968 13326 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16390 15008 16396 15020
rect 15979 14980 16396 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9548 14912 10057 14940
rect 9548 14900 9554 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12342 14940 12348 14952
rect 12124 14912 12348 14940
rect 12124 14900 12130 14912
rect 12342 14900 12348 14912
rect 12400 14940 12406 14952
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 12400 14912 12725 14940
rect 12400 14900 12406 14912
rect 12713 14909 12725 14912
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 12952 14912 13461 14940
rect 12952 14900 12958 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16206 14940 16212 14952
rect 16163 14912 16212 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 17144 14940 17172 14971
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17310 14968 17316 15020
rect 17368 14968 17374 15020
rect 17512 15017 17540 15048
rect 18414 15036 18420 15088
rect 18472 15076 18478 15088
rect 18782 15076 18788 15088
rect 18472 15048 18788 15076
rect 18472 15036 18478 15048
rect 18782 15036 18788 15048
rect 18840 15076 18846 15088
rect 19245 15079 19303 15085
rect 19245 15076 19257 15079
rect 18840 15048 19257 15076
rect 18840 15036 18846 15048
rect 19245 15045 19257 15048
rect 19291 15045 19303 15079
rect 19245 15039 19303 15045
rect 21910 15036 21916 15088
rect 21968 15076 21974 15088
rect 22465 15079 22523 15085
rect 22465 15076 22477 15079
rect 21968 15048 22477 15076
rect 21968 15036 21974 15048
rect 22465 15045 22477 15048
rect 22511 15045 22523 15079
rect 22465 15039 22523 15045
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17828 14980 18889 15008
rect 17828 14968 17834 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 21634 14968 21640 15020
rect 21692 15008 21698 15020
rect 22229 15011 22287 15017
rect 22229 15008 22241 15011
rect 21692 14980 22241 15008
rect 21692 14968 21698 14980
rect 22229 14977 22241 14980
rect 22275 14977 22287 15011
rect 22229 14971 22287 14977
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 22572 15008 22600 15116
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 23937 15147 23995 15153
rect 23937 15113 23949 15147
rect 23983 15144 23995 15147
rect 24854 15144 24860 15156
rect 23983 15116 24860 15144
rect 23983 15113 23995 15116
rect 23937 15107 23995 15113
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 27430 15104 27436 15156
rect 27488 15144 27494 15156
rect 27488 15116 28672 15144
rect 27488 15104 27494 15116
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 22664 15048 25697 15076
rect 22664 15017 22692 15048
rect 25685 15045 25697 15048
rect 25731 15076 25743 15079
rect 25731 15048 28304 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 22419 14980 22600 15008
rect 22649 15011 22707 15017
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22649 14977 22661 15011
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 18230 14940 18236 14952
rect 17144 14912 18236 14940
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 18463 14912 20116 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 18046 14872 18052 14884
rect 17552 14844 18052 14872
rect 17552 14832 17558 14844
rect 18046 14832 18052 14844
rect 18104 14832 18110 14884
rect 18138 14832 18144 14884
rect 18196 14872 18202 14884
rect 18432 14872 18460 14903
rect 18196 14844 18460 14872
rect 18196 14832 18202 14844
rect 19978 14832 19984 14884
rect 20036 14832 20042 14884
rect 20088 14872 20116 14912
rect 20346 14900 20352 14952
rect 20404 14900 20410 14952
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 22664 14940 22692 14971
rect 23198 14968 23204 15020
rect 23256 15008 23262 15020
rect 23566 15008 23572 15020
rect 23256 14980 23572 15008
rect 23256 14968 23262 14980
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 24394 14968 24400 15020
rect 24452 14968 24458 15020
rect 25406 14968 25412 15020
rect 25464 14968 25470 15020
rect 25590 14968 25596 15020
rect 25648 14968 25654 15020
rect 25829 15011 25887 15017
rect 25829 15008 25841 15011
rect 25700 14980 25841 15008
rect 20680 14912 22692 14940
rect 24136 14940 24164 14968
rect 24946 14940 24952 14952
rect 24136 14912 24952 14940
rect 20680 14900 20686 14912
rect 24946 14900 24952 14912
rect 25004 14900 25010 14952
rect 25038 14900 25044 14952
rect 25096 14940 25102 14952
rect 25700 14940 25728 14980
rect 25829 14977 25841 14980
rect 25875 15008 25887 15011
rect 26234 15008 26240 15020
rect 25875 14980 26240 15008
rect 25875 14977 25887 14980
rect 25829 14971 25887 14977
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 25096 14912 25728 14940
rect 27157 14943 27215 14949
rect 25096 14900 25102 14912
rect 27157 14909 27169 14943
rect 27203 14940 27215 14943
rect 27522 14940 27528 14952
rect 27203 14912 27528 14940
rect 27203 14909 27215 14912
rect 27157 14903 27215 14909
rect 27522 14900 27528 14912
rect 27580 14900 27586 14952
rect 27709 14943 27767 14949
rect 27709 14909 27721 14943
rect 27755 14940 27767 14943
rect 28169 14943 28227 14949
rect 28169 14940 28181 14943
rect 27755 14912 28181 14940
rect 27755 14909 27767 14912
rect 27709 14903 27767 14909
rect 28169 14909 28181 14912
rect 28215 14909 28227 14943
rect 28169 14903 28227 14909
rect 27617 14875 27675 14881
rect 27617 14872 27629 14875
rect 20088 14844 27629 14872
rect 27617 14841 27629 14844
rect 27663 14841 27675 14875
rect 27617 14835 27675 14841
rect 9490 14764 9496 14816
rect 9548 14764 9554 14816
rect 15749 14807 15807 14813
rect 15749 14773 15761 14807
rect 15795 14804 15807 14807
rect 16206 14804 16212 14816
rect 15795 14776 16212 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16853 14807 16911 14813
rect 16853 14773 16865 14807
rect 16899 14804 16911 14807
rect 16942 14804 16948 14816
rect 16899 14776 16948 14804
rect 16899 14773 16911 14776
rect 16853 14767 16911 14773
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 17957 14807 18015 14813
rect 17957 14804 17969 14807
rect 17920 14776 17969 14804
rect 17920 14764 17926 14776
rect 17957 14773 17969 14776
rect 18003 14773 18015 14807
rect 17957 14767 18015 14773
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 20162 14804 20168 14816
rect 19935 14776 20168 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 23106 14804 23112 14816
rect 20404 14776 23112 14804
rect 20404 14764 20410 14776
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 24305 14807 24363 14813
rect 24305 14773 24317 14807
rect 24351 14804 24363 14807
rect 24486 14804 24492 14816
rect 24351 14776 24492 14804
rect 24351 14773 24363 14776
rect 24305 14767 24363 14773
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 28166 14804 28172 14816
rect 26007 14776 28172 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 28166 14764 28172 14776
rect 28224 14764 28230 14816
rect 28276 14804 28304 15048
rect 28350 14968 28356 15020
rect 28408 14968 28414 15020
rect 28644 15017 28672 15116
rect 31754 15104 31760 15156
rect 31812 15104 31818 15156
rect 34974 15144 34980 15156
rect 33244 15116 34980 15144
rect 30644 15079 30702 15085
rect 30644 15045 30656 15079
rect 30690 15076 30702 15079
rect 31018 15076 31024 15088
rect 30690 15048 31024 15076
rect 30690 15045 30702 15048
rect 30644 15039 30702 15045
rect 31018 15036 31024 15048
rect 31076 15036 31082 15088
rect 31294 15036 31300 15088
rect 31352 15076 31358 15088
rect 33244 15085 33272 15116
rect 34974 15104 34980 15116
rect 35032 15144 35038 15156
rect 35434 15144 35440 15156
rect 35032 15116 35440 15144
rect 35032 15104 35038 15116
rect 35434 15104 35440 15116
rect 35492 15104 35498 15156
rect 33229 15079 33287 15085
rect 33229 15076 33241 15079
rect 31352 15048 33241 15076
rect 31352 15036 31358 15048
rect 33229 15045 33241 15048
rect 33275 15045 33287 15079
rect 33229 15039 33287 15045
rect 33870 15036 33876 15088
rect 33928 15076 33934 15088
rect 34854 15079 34912 15085
rect 34854 15076 34866 15079
rect 33928 15048 34866 15076
rect 33928 15036 33934 15048
rect 34854 15045 34866 15048
rect 34900 15045 34912 15079
rect 34854 15039 34912 15045
rect 38102 15036 38108 15088
rect 38160 15036 38166 15088
rect 28537 15011 28595 15017
rect 28537 14977 28549 15011
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 14977 28687 15011
rect 28629 14971 28687 14977
rect 28552 14940 28580 14971
rect 30926 14968 30932 15020
rect 30984 15008 30990 15020
rect 33597 15011 33655 15017
rect 33597 15008 33609 15011
rect 30984 14980 33609 15008
rect 30984 14968 30990 14980
rect 33597 14977 33609 14980
rect 33643 15008 33655 15011
rect 35342 15008 35348 15020
rect 33643 14980 35348 15008
rect 33643 14977 33655 14980
rect 33597 14971 33655 14977
rect 35342 14968 35348 14980
rect 35400 14968 35406 15020
rect 35710 14968 35716 15020
rect 35768 15008 35774 15020
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 35768 14980 37841 15008
rect 35768 14968 35774 14980
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 28994 14940 29000 14952
rect 28552 14912 29000 14940
rect 28994 14900 29000 14912
rect 29052 14940 29058 14952
rect 29638 14940 29644 14952
rect 29052 14912 29644 14940
rect 29052 14900 29058 14912
rect 29638 14900 29644 14912
rect 29696 14900 29702 14952
rect 30374 14900 30380 14952
rect 30432 14900 30438 14952
rect 32214 14900 32220 14952
rect 32272 14940 32278 14952
rect 33321 14943 33379 14949
rect 33321 14940 33333 14943
rect 32272 14912 33333 14940
rect 32272 14900 32278 14912
rect 33321 14909 33333 14912
rect 33367 14909 33379 14943
rect 33321 14903 33379 14909
rect 33410 14900 33416 14952
rect 33468 14940 33474 14952
rect 33689 14943 33747 14949
rect 33689 14940 33701 14943
rect 33468 14912 33701 14940
rect 33468 14900 33474 14912
rect 33689 14909 33701 14912
rect 33735 14909 33747 14943
rect 33689 14903 33747 14909
rect 34609 14943 34667 14949
rect 34609 14909 34621 14943
rect 34655 14909 34667 14943
rect 34609 14903 34667 14909
rect 33873 14875 33931 14881
rect 33873 14841 33885 14875
rect 33919 14872 33931 14875
rect 33962 14872 33968 14884
rect 33919 14844 33968 14872
rect 33919 14841 33931 14844
rect 33873 14835 33931 14841
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 34514 14804 34520 14816
rect 28276 14776 34520 14804
rect 34514 14764 34520 14776
rect 34572 14764 34578 14816
rect 34624 14804 34652 14903
rect 35710 14804 35716 14816
rect 34624 14776 35716 14804
rect 35710 14764 35716 14776
rect 35768 14764 35774 14816
rect 35986 14764 35992 14816
rect 36044 14764 36050 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 12894 14600 12900 14612
rect 12759 14572 12900 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13262 14560 13268 14612
rect 13320 14560 13326 14612
rect 17218 14560 17224 14612
rect 17276 14560 17282 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18288 14572 18705 14600
rect 18288 14560 18294 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 24394 14560 24400 14612
rect 24452 14600 24458 14612
rect 24857 14603 24915 14609
rect 24857 14600 24869 14603
rect 24452 14572 24869 14600
rect 24452 14560 24458 14572
rect 24857 14569 24869 14572
rect 24903 14569 24915 14603
rect 24857 14563 24915 14569
rect 25225 14603 25283 14609
rect 25225 14569 25237 14603
rect 25271 14600 25283 14603
rect 25590 14600 25596 14612
rect 25271 14572 25596 14600
rect 25271 14569 25283 14572
rect 25225 14563 25283 14569
rect 25590 14560 25596 14572
rect 25648 14560 25654 14612
rect 27157 14603 27215 14609
rect 27157 14569 27169 14603
rect 27203 14600 27215 14603
rect 27338 14600 27344 14612
rect 27203 14572 27344 14600
rect 27203 14569 27215 14572
rect 27157 14563 27215 14569
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 27522 14560 27528 14612
rect 27580 14600 27586 14612
rect 29270 14600 29276 14612
rect 27580 14572 29276 14600
rect 27580 14560 27586 14572
rect 29270 14560 29276 14572
rect 29328 14560 29334 14612
rect 31662 14560 31668 14612
rect 31720 14600 31726 14612
rect 35986 14600 35992 14612
rect 31720 14572 35992 14600
rect 31720 14560 31754 14572
rect 35986 14560 35992 14572
rect 36044 14560 36050 14612
rect 36081 14603 36139 14609
rect 36081 14569 36093 14603
rect 36127 14600 36139 14603
rect 36354 14600 36360 14612
rect 36127 14572 36360 14600
rect 36127 14569 36139 14572
rect 36081 14563 36139 14569
rect 36354 14560 36360 14572
rect 36412 14560 36418 14612
rect 37550 14560 37556 14612
rect 37608 14600 37614 14612
rect 38289 14603 38347 14609
rect 38289 14600 38301 14603
rect 37608 14572 38301 14600
rect 37608 14560 37614 14572
rect 38289 14569 38301 14572
rect 38335 14569 38347 14603
rect 38289 14563 38347 14569
rect 13354 14492 13360 14544
rect 13412 14492 13418 14544
rect 21358 14492 21364 14544
rect 21416 14532 21422 14544
rect 21453 14535 21511 14541
rect 21453 14532 21465 14535
rect 21416 14504 21465 14532
rect 21416 14492 21422 14504
rect 21453 14501 21465 14504
rect 21499 14501 21511 14535
rect 21453 14495 21511 14501
rect 26234 14492 26240 14544
rect 26292 14532 26298 14544
rect 31294 14532 31300 14544
rect 26292 14504 31300 14532
rect 26292 14492 26298 14504
rect 31294 14492 31300 14504
rect 31352 14492 31358 14544
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10560 14436 11529 14464
rect 10560 14424 10566 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 17862 14424 17868 14476
rect 17920 14424 17926 14476
rect 20162 14424 20168 14476
rect 20220 14424 20226 14476
rect 24946 14424 24952 14476
rect 25004 14424 25010 14476
rect 25314 14424 25320 14476
rect 25372 14464 25378 14476
rect 31726 14464 31754 14560
rect 32950 14492 32956 14544
rect 33008 14492 33014 14544
rect 34514 14492 34520 14544
rect 34572 14532 34578 14544
rect 35618 14532 35624 14544
rect 34572 14504 35624 14532
rect 34572 14492 34578 14504
rect 35618 14492 35624 14504
rect 35676 14492 35682 14544
rect 25372 14436 31754 14464
rect 32677 14467 32735 14473
rect 25372 14424 25378 14436
rect 32677 14433 32689 14467
rect 32723 14464 32735 14467
rect 33042 14464 33048 14476
rect 32723 14436 33048 14464
rect 32723 14433 32735 14436
rect 32677 14427 32735 14433
rect 33042 14424 33048 14436
rect 33100 14424 33106 14476
rect 35434 14424 35440 14476
rect 35492 14424 35498 14476
rect 35710 14424 35716 14476
rect 35768 14464 35774 14476
rect 36909 14467 36967 14473
rect 36909 14464 36921 14467
rect 35768 14436 36921 14464
rect 35768 14424 35774 14436
rect 36909 14433 36921 14436
rect 36955 14433 36967 14467
rect 36909 14427 36967 14433
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11790 14396 11796 14408
rect 11655 14368 11796 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14396 12863 14399
rect 14182 14396 14188 14408
rect 12851 14368 14188 14396
rect 12851 14365 12863 14368
rect 12805 14359 12863 14365
rect 12069 14331 12127 14337
rect 12069 14297 12081 14331
rect 12115 14328 12127 14331
rect 12250 14328 12256 14340
rect 12115 14300 12256 14328
rect 12115 14297 12127 14300
rect 12069 14291 12127 14297
rect 12250 14288 12256 14300
rect 12308 14328 12314 14340
rect 12636 14328 12664 14359
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 17586 14356 17592 14408
rect 17644 14356 17650 14408
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 12894 14328 12900 14340
rect 12308 14300 12434 14328
rect 12636 14300 12900 14328
rect 12308 14288 12314 14300
rect 12406 14260 12434 14300
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13725 14331 13783 14337
rect 13725 14297 13737 14331
rect 13771 14328 13783 14331
rect 13998 14328 14004 14340
rect 13771 14300 14004 14328
rect 13771 14297 13783 14300
rect 13725 14291 13783 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 15102 14288 15108 14340
rect 15160 14288 15166 14340
rect 15470 14288 15476 14340
rect 15528 14288 15534 14340
rect 17604 14328 17632 14356
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 17604 14300 17693 14328
rect 17681 14297 17693 14300
rect 17727 14328 17739 14331
rect 18506 14328 18512 14340
rect 17727 14300 18512 14328
rect 17727 14297 17739 14300
rect 17681 14291 17739 14297
rect 18506 14288 18512 14300
rect 18564 14328 18570 14340
rect 18708 14328 18736 14359
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18840 14368 18889 14396
rect 18840 14356 18846 14368
rect 18877 14365 18889 14368
rect 18923 14396 18935 14399
rect 18966 14396 18972 14408
rect 18923 14368 18972 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 21634 14405 21640 14408
rect 21632 14396 21640 14405
rect 21595 14368 21640 14396
rect 21632 14359 21640 14368
rect 21634 14356 21640 14359
rect 21692 14356 21698 14408
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 21910 14396 21916 14408
rect 21867 14368 21916 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 23934 14356 23940 14408
rect 23992 14396 23998 14408
rect 24394 14396 24400 14408
rect 23992 14368 24400 14396
rect 23992 14356 23998 14368
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 24486 14356 24492 14408
rect 24544 14396 24550 14408
rect 24857 14399 24915 14405
rect 24857 14396 24869 14399
rect 24544 14368 24869 14396
rect 24544 14356 24550 14368
rect 24857 14365 24869 14368
rect 24903 14365 24915 14399
rect 24857 14359 24915 14365
rect 18564 14300 20116 14328
rect 18564 14288 18570 14300
rect 15194 14260 15200 14272
rect 12406 14232 15200 14260
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17276 14232 17601 14260
rect 17276 14220 17282 14232
rect 17589 14229 17601 14232
rect 17635 14260 17647 14263
rect 17770 14260 17776 14272
rect 17635 14232 17776 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 18932 14232 19625 14260
rect 18932 14220 18938 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 19978 14220 19984 14272
rect 20036 14220 20042 14272
rect 20088 14269 20116 14300
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 22020 14328 22048 14356
rect 23753 14331 23811 14337
rect 23753 14328 23765 14331
rect 21048 14300 22048 14328
rect 23492 14300 23765 14328
rect 21048 14288 21054 14300
rect 23492 14272 23520 14300
rect 23753 14297 23765 14300
rect 23799 14297 23811 14331
rect 24872 14328 24900 14359
rect 26602 14356 26608 14408
rect 26660 14396 26666 14408
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 26660 14368 27077 14396
rect 26660 14356 26666 14368
rect 27065 14365 27077 14368
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 27154 14356 27160 14408
rect 27212 14396 27218 14408
rect 30650 14396 30656 14408
rect 27212 14368 30656 14396
rect 27212 14356 27218 14368
rect 30650 14356 30656 14368
rect 30708 14356 30714 14408
rect 35342 14356 35348 14408
rect 35400 14396 35406 14408
rect 37182 14405 37188 14408
rect 35805 14399 35863 14405
rect 35805 14396 35817 14399
rect 35400 14368 35817 14396
rect 35400 14356 35406 14368
rect 35805 14365 35817 14368
rect 35851 14365 35863 14399
rect 35805 14359 35863 14365
rect 35897 14399 35955 14405
rect 35897 14365 35909 14399
rect 35943 14365 35955 14399
rect 37176 14396 37188 14405
rect 37143 14368 37188 14396
rect 35897 14359 35955 14365
rect 37176 14359 37188 14368
rect 29822 14328 29828 14340
rect 24872 14300 29828 14328
rect 23753 14291 23811 14297
rect 29822 14288 29828 14300
rect 29880 14288 29886 14340
rect 35526 14328 35532 14340
rect 29932 14300 35532 14328
rect 20073 14263 20131 14269
rect 20073 14229 20085 14263
rect 20119 14260 20131 14263
rect 20806 14260 20812 14272
rect 20119 14232 20812 14260
rect 20119 14229 20131 14232
rect 20073 14223 20131 14229
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 21082 14220 21088 14272
rect 21140 14260 21146 14272
rect 23474 14260 23480 14272
rect 21140 14232 23480 14260
rect 21140 14220 21146 14232
rect 23474 14220 23480 14232
rect 23532 14220 23538 14272
rect 23569 14263 23627 14269
rect 23569 14229 23581 14263
rect 23615 14260 23627 14263
rect 24210 14260 24216 14272
rect 23615 14232 24216 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 28994 14260 29000 14272
rect 25004 14232 29000 14260
rect 25004 14220 25010 14232
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 29086 14220 29092 14272
rect 29144 14260 29150 14272
rect 29932 14260 29960 14300
rect 35526 14288 35532 14300
rect 35584 14288 35590 14340
rect 35618 14288 35624 14340
rect 35676 14328 35682 14340
rect 35912 14328 35940 14359
rect 37182 14356 37188 14359
rect 37240 14356 37246 14408
rect 35676 14300 35940 14328
rect 35676 14288 35682 14300
rect 29144 14232 29960 14260
rect 33137 14263 33195 14269
rect 29144 14220 29150 14232
rect 33137 14229 33149 14263
rect 33183 14260 33195 14263
rect 33686 14260 33692 14272
rect 33183 14232 33692 14260
rect 33183 14229 33195 14232
rect 33137 14223 33195 14229
rect 33686 14220 33692 14232
rect 33744 14220 33750 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9217 14059 9275 14065
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 9858 14056 9864 14068
rect 9263 14028 9864 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 13170 14056 13176 14068
rect 12207 14028 13176 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 17368 14028 17509 14056
rect 17368 14016 17374 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 18874 14056 18880 14068
rect 17497 14019 17555 14025
rect 18616 14028 18880 14056
rect 8104 13991 8162 13997
rect 8104 13957 8116 13991
rect 8150 13988 8162 13991
rect 9490 13988 9496 14000
rect 8150 13960 9496 13988
rect 8150 13957 8162 13960
rect 8104 13951 8162 13957
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 9876 13988 9904 14016
rect 9876 13960 10732 13988
rect 7834 13880 7840 13932
rect 7892 13880 7898 13932
rect 10410 13880 10416 13932
rect 10468 13880 10474 13932
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 10704 13852 10732 13960
rect 11790 13948 11796 14000
rect 11848 13948 11854 14000
rect 13081 13991 13139 13997
rect 13081 13957 13093 13991
rect 13127 13988 13139 13991
rect 14182 13988 14188 14000
rect 13127 13960 14188 13988
rect 13127 13957 13139 13960
rect 13081 13951 13139 13957
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 15470 13948 15476 14000
rect 15528 13988 15534 14000
rect 16853 13991 16911 13997
rect 16853 13988 16865 13991
rect 15528 13960 16865 13988
rect 15528 13948 15534 13960
rect 16853 13957 16865 13960
rect 16899 13988 16911 13991
rect 18138 13988 18144 14000
rect 16899 13960 18144 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 18230 13948 18236 14000
rect 18288 13988 18294 14000
rect 18288 13960 18552 13988
rect 18288 13948 18294 13960
rect 11808 13920 11836 13948
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11808 13892 11989 13920
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 13998 13920 14004 13932
rect 13495 13892 14004 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 10704 13824 11805 13852
rect 11793 13821 11805 13824
rect 11839 13852 11851 13855
rect 11882 13852 11888 13864
rect 11839 13824 11888 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12894 13812 12900 13864
rect 12952 13812 12958 13864
rect 13004 13852 13032 13883
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14550 13880 14556 13932
rect 14608 13920 14614 13932
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 14608 13892 14749 13920
rect 14608 13880 14614 13892
rect 14737 13889 14749 13892
rect 14783 13920 14795 13923
rect 15102 13920 15108 13932
rect 14783 13892 15108 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 17092 13892 17325 13920
rect 17092 13880 17098 13892
rect 17313 13889 17325 13892
rect 17359 13920 17371 13923
rect 17494 13920 17500 13932
rect 17359 13892 17500 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 17770 13880 17776 13932
rect 17828 13920 17834 13932
rect 18524 13929 18552 13960
rect 18616 13929 18644 14028
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 24118 14056 24124 14068
rect 23523 14028 24124 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 25225 14059 25283 14065
rect 25225 14025 25237 14059
rect 25271 14056 25283 14059
rect 30926 14056 30932 14068
rect 25271 14028 30932 14056
rect 25271 14025 25283 14028
rect 25225 14019 25283 14025
rect 30926 14016 30932 14028
rect 30984 14016 30990 14068
rect 19337 13991 19395 13997
rect 19337 13988 19349 13991
rect 18708 13960 19349 13988
rect 18708 13929 18736 13960
rect 19337 13957 19349 13960
rect 19383 13957 19395 13991
rect 19978 13988 19984 14000
rect 19337 13951 19395 13957
rect 19628 13960 19984 13988
rect 18509 13923 18567 13929
rect 17828 13892 18368 13920
rect 17828 13880 17834 13892
rect 13354 13852 13360 13864
rect 13004 13824 13360 13852
rect 13354 13812 13360 13824
rect 13412 13852 13418 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 13412 13824 14381 13852
rect 13412 13812 13418 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 15010 13812 15016 13864
rect 15068 13812 15074 13864
rect 17218 13812 17224 13864
rect 17276 13812 17282 13864
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 18233 13855 18291 13861
rect 18233 13852 18245 13855
rect 17460 13824 18245 13852
rect 17460 13812 17466 13824
rect 18233 13821 18245 13824
rect 18279 13821 18291 13855
rect 18340 13852 18368 13892
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18693 13923 18751 13929
rect 18693 13889 18705 13923
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 18874 13880 18880 13932
rect 18932 13880 18938 13932
rect 19628 13929 19656 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 22741 13991 22799 13997
rect 22741 13957 22753 13991
rect 22787 13988 22799 13991
rect 22787 13960 24256 13988
rect 22787 13957 22799 13960
rect 22741 13951 22799 13957
rect 24228 13932 24256 13960
rect 25590 13948 25596 14000
rect 25648 13988 25654 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25648 13960 25881 13988
rect 25648 13948 25654 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 18984 13892 19625 13920
rect 18984 13852 19012 13892
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 20070 13920 20076 13932
rect 19613 13883 19671 13889
rect 19904 13892 20076 13920
rect 18340 13824 19012 13852
rect 18233 13815 18291 13821
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19484 13824 19533 13852
rect 19484 13812 19490 13824
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 19904 13852 19932 13892
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22925 13923 22983 13929
rect 22695 13892 22876 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 19567 13824 19932 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 20346 13852 20352 13864
rect 20036 13824 20352 13852
rect 20036 13812 20042 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 10781 13787 10839 13793
rect 10781 13753 10793 13787
rect 10827 13784 10839 13787
rect 13814 13784 13820 13796
rect 10827 13756 13820 13784
rect 10827 13753 10839 13756
rect 10781 13747 10839 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 13909 13787 13967 13793
rect 13909 13753 13921 13787
rect 13955 13784 13967 13787
rect 15838 13784 15844 13796
rect 13955 13756 15844 13784
rect 13955 13753 13967 13756
rect 13909 13747 13967 13753
rect 15838 13744 15844 13756
rect 15896 13744 15902 13796
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10962 13716 10968 13728
rect 10284 13688 10968 13716
rect 10284 13676 10290 13688
rect 10962 13676 10968 13688
rect 11020 13716 11026 13728
rect 15562 13716 15568 13728
rect 11020 13688 15568 13716
rect 11020 13676 11026 13688
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 22848 13716 22876 13892
rect 22925 13889 22937 13923
rect 22971 13920 22983 13923
rect 23474 13920 23480 13932
rect 22971 13892 23480 13920
rect 22971 13889 22983 13892
rect 22925 13883 22983 13889
rect 23474 13880 23480 13892
rect 23532 13880 23538 13932
rect 23750 13880 23756 13932
rect 23808 13880 23814 13932
rect 24026 13880 24032 13932
rect 24084 13880 24090 13932
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24268 13892 25053 13920
rect 24268 13880 24274 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 25682 13880 25688 13932
rect 25740 13920 25746 13932
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 25740 13892 25789 13920
rect 25740 13880 25746 13892
rect 25777 13889 25789 13892
rect 25823 13889 25835 13923
rect 25884 13920 25912 13951
rect 26050 13948 26056 14000
rect 26108 13948 26114 14000
rect 27982 13948 27988 14000
rect 28040 13948 28046 14000
rect 28442 13948 28448 14000
rect 28500 13948 28506 14000
rect 28534 13948 28540 14000
rect 28592 13988 28598 14000
rect 29086 13988 29092 14000
rect 28592 13960 29092 13988
rect 28592 13948 28598 13960
rect 29086 13948 29092 13960
rect 29144 13948 29150 14000
rect 29638 13948 29644 14000
rect 29696 13988 29702 14000
rect 35618 13988 35624 14000
rect 29696 13960 35624 13988
rect 29696 13948 29702 13960
rect 27154 13920 27160 13932
rect 25884 13892 27160 13920
rect 25777 13883 25835 13889
rect 23615 13855 23673 13861
rect 23615 13852 23627 13855
rect 22940 13824 23627 13852
rect 22940 13793 22968 13824
rect 23615 13821 23627 13824
rect 23661 13821 23673 13855
rect 23615 13815 23673 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24302 13852 24308 13864
rect 24167 13824 24308 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 24581 13855 24639 13861
rect 24581 13821 24593 13855
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 22925 13787 22983 13793
rect 22925 13753 22937 13787
rect 22971 13753 22983 13787
rect 22925 13747 22983 13753
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 24486 13784 24492 13796
rect 23348 13756 24492 13784
rect 23348 13744 23354 13756
rect 24486 13744 24492 13756
rect 24544 13744 24550 13796
rect 23658 13716 23664 13728
rect 22848 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13716 23722 13728
rect 24596 13716 24624 13815
rect 24854 13812 24860 13864
rect 24912 13852 24918 13864
rect 24949 13855 25007 13861
rect 24949 13852 24961 13855
rect 24912 13824 24961 13852
rect 24912 13812 24918 13824
rect 24949 13821 24961 13824
rect 24995 13821 25007 13855
rect 25792 13852 25820 13883
rect 27154 13880 27160 13892
rect 27212 13880 27218 13932
rect 27709 13923 27767 13929
rect 27709 13889 27721 13923
rect 27755 13889 27767 13923
rect 27709 13883 27767 13889
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 27430 13852 27436 13864
rect 25792 13824 27436 13852
rect 24949 13815 25007 13821
rect 27430 13812 27436 13824
rect 27488 13852 27494 13864
rect 27724 13852 27752 13883
rect 27488 13824 27752 13852
rect 27816 13852 27844 13883
rect 27890 13880 27896 13932
rect 27948 13920 27954 13932
rect 28813 13923 28871 13929
rect 28813 13920 28825 13923
rect 27948 13892 28825 13920
rect 27948 13880 27954 13892
rect 28813 13889 28825 13892
rect 28859 13889 28871 13923
rect 28813 13883 28871 13889
rect 28534 13852 28540 13864
rect 27816 13824 28540 13852
rect 27488 13812 27494 13824
rect 28534 13812 28540 13824
rect 28592 13812 28598 13864
rect 28828 13852 28856 13883
rect 28994 13880 29000 13932
rect 29052 13880 29058 13932
rect 29454 13880 29460 13932
rect 29512 13880 29518 13932
rect 30024 13929 30052 13960
rect 35618 13948 35624 13960
rect 35676 13948 35682 14000
rect 30009 13923 30067 13929
rect 30009 13889 30021 13923
rect 30055 13889 30067 13923
rect 30009 13883 30067 13889
rect 30098 13880 30104 13932
rect 30156 13880 30162 13932
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 31294 13880 31300 13932
rect 31352 13880 31358 13932
rect 33226 13880 33232 13932
rect 33284 13880 33290 13932
rect 29730 13852 29736 13864
rect 28828 13824 29736 13852
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 31018 13812 31024 13864
rect 31076 13812 31082 13864
rect 31757 13855 31815 13861
rect 31757 13821 31769 13855
rect 31803 13852 31815 13855
rect 32306 13852 32312 13864
rect 31803 13824 32312 13852
rect 31803 13821 31815 13824
rect 31757 13815 31815 13821
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 33321 13855 33379 13861
rect 33321 13821 33333 13855
rect 33367 13852 33379 13855
rect 33594 13852 33600 13864
rect 33367 13824 33600 13852
rect 33367 13821 33379 13824
rect 33321 13815 33379 13821
rect 33594 13812 33600 13824
rect 33652 13812 33658 13864
rect 38286 13812 38292 13864
rect 38344 13812 38350 13864
rect 28813 13787 28871 13793
rect 28813 13753 28825 13787
rect 28859 13784 28871 13787
rect 28902 13784 28908 13796
rect 28859 13756 28908 13784
rect 28859 13753 28871 13756
rect 28813 13747 28871 13753
rect 28902 13744 28908 13756
rect 28960 13744 28966 13796
rect 29917 13787 29975 13793
rect 29917 13753 29929 13787
rect 29963 13753 29975 13787
rect 29917 13747 29975 13753
rect 23716 13688 24624 13716
rect 23716 13676 23722 13688
rect 25590 13676 25596 13728
rect 25648 13716 25654 13728
rect 26053 13719 26111 13725
rect 26053 13716 26065 13719
rect 25648 13688 26065 13716
rect 25648 13676 25654 13688
rect 26053 13685 26065 13688
rect 26099 13685 26111 13719
rect 26053 13679 26111 13685
rect 27982 13676 27988 13728
rect 28040 13676 28046 13728
rect 29932 13716 29960 13747
rect 30006 13716 30012 13728
rect 29932 13688 30012 13716
rect 30006 13676 30012 13688
rect 30064 13676 30070 13728
rect 33505 13719 33563 13725
rect 33505 13685 33517 13719
rect 33551 13716 33563 13719
rect 34790 13716 34796 13728
rect 33551 13688 34796 13716
rect 33551 13685 33563 13688
rect 33505 13679 33563 13685
rect 34790 13676 34796 13688
rect 34848 13676 34854 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15068 13484 15485 13512
rect 15068 13472 15074 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 22462 13512 22468 13524
rect 15473 13475 15531 13481
rect 15672 13484 22468 13512
rect 10502 13404 10508 13456
rect 10560 13404 10566 13456
rect 15028 13444 15056 13472
rect 14384 13416 15056 13444
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 14384 13385 14412 13416
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15286 13376 15292 13388
rect 14967 13348 15292 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10192 13280 12434 13308
rect 10192 13268 10198 13280
rect 12406 13240 12434 13280
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 15672 13240 15700 13484
rect 22462 13472 22468 13484
rect 22520 13512 22526 13524
rect 23290 13512 23296 13524
rect 22520 13484 23296 13512
rect 22520 13472 22526 13484
rect 23290 13472 23296 13484
rect 23348 13472 23354 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23750 13512 23756 13524
rect 23523 13484 23756 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 26326 13472 26332 13524
rect 26384 13512 26390 13524
rect 29178 13512 29184 13524
rect 26384 13484 29184 13512
rect 26384 13472 26390 13484
rect 29178 13472 29184 13484
rect 29236 13472 29242 13524
rect 31018 13472 31024 13524
rect 31076 13512 31082 13524
rect 31205 13515 31263 13521
rect 31205 13512 31217 13515
rect 31076 13484 31217 13512
rect 31076 13472 31082 13484
rect 31205 13481 31217 13484
rect 31251 13481 31263 13515
rect 31205 13475 31263 13481
rect 33045 13515 33103 13521
rect 33045 13481 33057 13515
rect 33091 13512 33103 13515
rect 33226 13512 33232 13524
rect 33091 13484 33232 13512
rect 33091 13481 33103 13484
rect 33045 13475 33103 13481
rect 33226 13472 33232 13484
rect 33284 13472 33290 13524
rect 28629 13447 28687 13453
rect 15856 13416 25084 13444
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 15856 13376 15884 13416
rect 16574 13376 16580 13388
rect 15804 13348 15884 13376
rect 15804 13336 15810 13348
rect 15856 13317 15884 13348
rect 16224 13348 16580 13376
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 16114 13268 16120 13320
rect 16172 13268 16178 13320
rect 16224 13317 16252 13348
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 16485 13271 16543 13277
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 16807 13280 17325 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 12406 13212 15700 13240
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14553 13175 14611 13181
rect 14553 13172 14565 13175
rect 14056 13144 14565 13172
rect 14056 13132 14062 13144
rect 14553 13141 14565 13144
rect 14599 13141 14611 13175
rect 14553 13135 14611 13141
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 16500 13172 16528 13271
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 17788 13317 17816 13416
rect 21358 13376 21364 13388
rect 21008 13348 21364 13376
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 20806 13268 20812 13320
rect 20864 13268 20870 13320
rect 21008 13317 21036 13348
rect 21358 13336 21364 13348
rect 21416 13376 21422 13388
rect 21416 13348 21680 13376
rect 21416 13336 21422 13348
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21324 13280 21465 13308
rect 21324 13268 21330 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 21542 13268 21548 13320
rect 21600 13268 21606 13320
rect 21652 13308 21680 13348
rect 21726 13336 21732 13388
rect 21784 13336 21790 13388
rect 23658 13336 23664 13388
rect 23716 13336 23722 13388
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13376 23811 13379
rect 24210 13376 24216 13388
rect 23799 13348 24216 13376
rect 23799 13345 23811 13348
rect 23753 13339 23811 13345
rect 24210 13336 24216 13348
rect 24268 13336 24274 13388
rect 25056 13385 25084 13416
rect 28629 13413 28641 13447
rect 28675 13444 28687 13447
rect 29638 13444 29644 13456
rect 28675 13416 29644 13444
rect 28675 13413 28687 13416
rect 28629 13407 28687 13413
rect 29638 13404 29644 13416
rect 29696 13404 29702 13456
rect 30285 13447 30343 13453
rect 30285 13413 30297 13447
rect 30331 13444 30343 13447
rect 30331 13416 30880 13444
rect 30331 13413 30343 13416
rect 30285 13407 30343 13413
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 25593 13379 25651 13385
rect 25593 13345 25605 13379
rect 25639 13376 25651 13379
rect 25958 13376 25964 13388
rect 25639 13348 25964 13376
rect 25639 13345 25651 13348
rect 25593 13339 25651 13345
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 26053 13379 26111 13385
rect 26053 13345 26065 13379
rect 26099 13376 26111 13379
rect 26602 13376 26608 13388
rect 26099 13348 26608 13376
rect 26099 13345 26111 13348
rect 26053 13339 26111 13345
rect 26602 13336 26608 13348
rect 26660 13376 26666 13388
rect 26660 13348 27752 13376
rect 26660 13336 26666 13348
rect 22002 13308 22008 13320
rect 21652 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23532 13280 23857 13308
rect 23532 13268 23538 13280
rect 23845 13277 23857 13280
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13308 23995 13311
rect 24026 13308 24032 13320
rect 23983 13280 24032 13308
rect 23983 13277 23995 13280
rect 23937 13271 23995 13277
rect 17512 13240 17540 13268
rect 19518 13240 19524 13252
rect 17512 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 22370 13240 22376 13252
rect 20947 13212 22376 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 22370 13200 22376 13212
rect 22428 13200 22434 13252
rect 23860 13240 23888 13271
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24486 13268 24492 13320
rect 24544 13308 24550 13320
rect 24544 13280 25820 13308
rect 24544 13268 24550 13280
rect 24762 13240 24768 13252
rect 23860 13212 24768 13240
rect 24762 13200 24768 13212
rect 24820 13200 24826 13252
rect 25792 13240 25820 13280
rect 25866 13268 25872 13320
rect 25924 13268 25930 13320
rect 26436 13280 26740 13308
rect 26436 13240 26464 13280
rect 25792 13212 26464 13240
rect 26510 13200 26516 13252
rect 26568 13200 26574 13252
rect 26712 13240 26740 13280
rect 26786 13268 26792 13320
rect 26844 13308 26850 13320
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 26844 13280 27169 13308
rect 26844 13268 26850 13280
rect 27157 13277 27169 13280
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 27246 13268 27252 13320
rect 27304 13268 27310 13320
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 27356 13280 27537 13308
rect 27356 13240 27384 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 27617 13311 27675 13317
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27724 13308 27752 13348
rect 27982 13336 27988 13388
rect 28040 13376 28046 13388
rect 28445 13379 28503 13385
rect 28445 13376 28457 13379
rect 28040 13348 28457 13376
rect 28040 13336 28046 13348
rect 28445 13345 28457 13348
rect 28491 13345 28503 13379
rect 28445 13339 28503 13345
rect 29822 13336 29828 13388
rect 29880 13336 29886 13388
rect 30852 13385 30880 13416
rect 32950 13404 32956 13456
rect 33008 13404 33014 13456
rect 30837 13379 30895 13385
rect 30837 13345 30849 13379
rect 30883 13345 30895 13379
rect 30837 13339 30895 13345
rect 32585 13379 32643 13385
rect 32585 13345 32597 13379
rect 32631 13376 32643 13379
rect 32858 13376 32864 13388
rect 32631 13348 32864 13376
rect 32631 13345 32643 13348
rect 32585 13339 32643 13345
rect 32858 13336 32864 13348
rect 32916 13336 32922 13388
rect 34606 13336 34612 13388
rect 34664 13376 34670 13388
rect 35710 13376 35716 13388
rect 34664 13348 35716 13376
rect 34664 13336 34670 13348
rect 35710 13336 35716 13348
rect 35768 13336 35774 13388
rect 28721 13311 28779 13317
rect 28721 13308 28733 13311
rect 27724 13280 28733 13308
rect 27617 13271 27675 13277
rect 28721 13277 28733 13280
rect 28767 13277 28779 13311
rect 28721 13271 28779 13277
rect 26712 13212 27384 13240
rect 27430 13200 27436 13252
rect 27488 13240 27494 13252
rect 27632 13240 27660 13271
rect 29086 13268 29092 13320
rect 29144 13308 29150 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29144 13280 29929 13308
rect 29144 13268 29150 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 30926 13268 30932 13320
rect 30984 13268 30990 13320
rect 33226 13268 33232 13320
rect 33284 13308 33290 13320
rect 33505 13311 33563 13317
rect 33505 13308 33517 13311
rect 33284 13280 33517 13308
rect 33284 13268 33290 13280
rect 33505 13277 33517 13280
rect 33551 13277 33563 13311
rect 33505 13271 33563 13277
rect 33686 13268 33692 13320
rect 33744 13268 33750 13320
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 35969 13311 36027 13317
rect 35969 13308 35981 13311
rect 34848 13280 35981 13308
rect 34848 13268 34854 13280
rect 35969 13277 35981 13280
rect 36015 13277 36027 13311
rect 35969 13271 36027 13277
rect 27488 13212 27660 13240
rect 27488 13200 27494 13212
rect 15712 13144 16528 13172
rect 21729 13175 21787 13181
rect 15712 13132 15718 13144
rect 21729 13141 21741 13175
rect 21775 13172 21787 13175
rect 22186 13172 22192 13184
rect 21775 13144 22192 13172
rect 21775 13141 21787 13144
rect 21729 13135 21787 13141
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 28261 13175 28319 13181
rect 28261 13172 28273 13175
rect 22520 13144 28273 13172
rect 22520 13132 22526 13144
rect 28261 13141 28273 13144
rect 28307 13141 28319 13175
rect 28261 13135 28319 13141
rect 33597 13175 33655 13181
rect 33597 13141 33609 13175
rect 33643 13172 33655 13175
rect 33778 13172 33784 13184
rect 33643 13144 33784 13172
rect 33643 13141 33655 13144
rect 33597 13135 33655 13141
rect 33778 13132 33784 13144
rect 33836 13132 33842 13184
rect 35802 13132 35808 13184
rect 35860 13172 35866 13184
rect 37093 13175 37151 13181
rect 37093 13172 37105 13175
rect 35860 13144 37105 13172
rect 35860 13132 35866 13144
rect 37093 13141 37105 13144
rect 37139 13141 37151 13175
rect 37093 13135 37151 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 12894 12928 12900 12980
rect 12952 12968 12958 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 12952 12940 13461 12968
rect 12952 12928 12958 12940
rect 13449 12937 13461 12940
rect 13495 12937 13507 12971
rect 13449 12931 13507 12937
rect 21266 12928 21272 12980
rect 21324 12968 21330 12980
rect 22462 12968 22468 12980
rect 21324 12940 22468 12968
rect 21324 12928 21330 12940
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 23569 12971 23627 12977
rect 23569 12937 23581 12971
rect 23615 12968 23627 12971
rect 23658 12968 23664 12980
rect 23615 12940 23664 12968
rect 23615 12937 23627 12940
rect 23569 12931 23627 12937
rect 23658 12928 23664 12940
rect 23716 12928 23722 12980
rect 27246 12928 27252 12980
rect 27304 12968 27310 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 27304 12940 28549 12968
rect 27304 12928 27310 12940
rect 28537 12937 28549 12940
rect 28583 12937 28595 12971
rect 28537 12931 28595 12937
rect 34698 12928 34704 12980
rect 34756 12968 34762 12980
rect 35069 12971 35127 12977
rect 35069 12968 35081 12971
rect 34756 12940 35081 12968
rect 34756 12928 34762 12940
rect 35069 12937 35081 12940
rect 35115 12937 35127 12971
rect 35069 12931 35127 12937
rect 7834 12900 7840 12912
rect 7392 12872 7840 12900
rect 7392 12841 7420 12872
rect 7834 12860 7840 12872
rect 7892 12860 7898 12912
rect 13262 12900 13268 12912
rect 9324 12872 13268 12900
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7644 12835 7702 12841
rect 7644 12801 7656 12835
rect 7690 12832 7702 12835
rect 9324 12832 9352 12872
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 15470 12860 15476 12912
rect 15528 12860 15534 12912
rect 15562 12860 15568 12912
rect 15620 12900 15626 12912
rect 16114 12900 16120 12912
rect 15620 12872 16120 12900
rect 15620 12860 15626 12872
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 21100 12872 22017 12900
rect 7690 12804 9352 12832
rect 7690 12801 7702 12804
rect 7644 12795 7702 12801
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12832 12403 12835
rect 12710 12832 12716 12844
rect 12391 12804 12716 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 10410 12764 10416 12776
rect 9815 12736 10416 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 9324 12696 9352 12727
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 12084 12764 12112 12795
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12832 13599 12835
rect 13630 12832 13636 12844
rect 13587 12804 13636 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 12894 12764 12900 12776
rect 12084 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13170 12724 13176 12776
rect 13228 12764 13234 12776
rect 13372 12764 13400 12795
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 15252 12804 15301 12832
rect 15252 12792 15258 12804
rect 15289 12801 15301 12804
rect 15335 12801 15347 12835
rect 16574 12832 16580 12844
rect 15289 12795 15347 12801
rect 15396 12804 16580 12832
rect 15396 12764 15424 12804
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17368 12804 17417 12832
rect 17368 12792 17374 12804
rect 17405 12801 17417 12804
rect 17451 12832 17463 12835
rect 17678 12832 17684 12844
rect 17451 12804 17684 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 17678 12792 17684 12804
rect 17736 12792 17742 12844
rect 21100 12841 21128 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 26510 12900 26516 12912
rect 22005 12863 22063 12869
rect 22296 12872 26516 12900
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 21174 12792 21180 12844
rect 21232 12792 21238 12844
rect 21358 12792 21364 12844
rect 21416 12832 21422 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 21416 12804 21465 12832
rect 21416 12792 21422 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 13228 12736 15424 12764
rect 13228 12724 13234 12736
rect 17218 12724 17224 12776
rect 17276 12724 17282 12776
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 22296 12764 22324 12872
rect 26510 12860 26516 12872
rect 26568 12860 26574 12912
rect 34606 12900 34612 12912
rect 26620 12872 28028 12900
rect 26620 12844 26648 12872
rect 22370 12792 22376 12844
rect 22428 12792 22434 12844
rect 22462 12792 22468 12844
rect 22520 12792 22526 12844
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12832 23719 12835
rect 23934 12832 23940 12844
rect 23707 12804 23940 12832
rect 23707 12801 23719 12804
rect 23661 12795 23719 12801
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 25590 12792 25596 12844
rect 25648 12792 25654 12844
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12832 25927 12835
rect 26602 12832 26608 12844
rect 25915 12804 26608 12832
rect 25915 12801 25927 12804
rect 25869 12795 25927 12801
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 27890 12792 27896 12844
rect 27948 12792 27954 12844
rect 28000 12841 28028 12872
rect 33704 12872 34612 12900
rect 27985 12835 28043 12841
rect 27985 12801 27997 12835
rect 28031 12832 28043 12835
rect 28445 12835 28503 12841
rect 28445 12832 28457 12835
rect 28031 12804 28457 12832
rect 28031 12801 28043 12804
rect 27985 12795 28043 12801
rect 28445 12801 28457 12804
rect 28491 12801 28503 12835
rect 28445 12795 28503 12801
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12832 28687 12835
rect 29362 12832 29368 12844
rect 28675 12804 29368 12832
rect 28675 12801 28687 12804
rect 28629 12795 28687 12801
rect 29362 12792 29368 12804
rect 29420 12792 29426 12844
rect 33134 12792 33140 12844
rect 33192 12832 33198 12844
rect 33704 12841 33732 12872
rect 34606 12860 34612 12872
rect 34664 12860 34670 12912
rect 33689 12835 33747 12841
rect 33689 12832 33701 12835
rect 33192 12804 33701 12832
rect 33192 12792 33198 12804
rect 33689 12801 33701 12804
rect 33735 12801 33747 12835
rect 33689 12795 33747 12801
rect 33778 12792 33784 12844
rect 33836 12832 33842 12844
rect 33945 12835 34003 12841
rect 33945 12832 33957 12835
rect 33836 12804 33957 12832
rect 33836 12792 33842 12804
rect 33945 12801 33957 12804
rect 33991 12801 34003 12835
rect 33945 12795 34003 12801
rect 17552 12736 22324 12764
rect 25777 12767 25835 12773
rect 17552 12724 17558 12736
rect 25777 12733 25789 12767
rect 25823 12764 25835 12767
rect 26326 12764 26332 12776
rect 25823 12736 26332 12764
rect 25823 12733 25835 12736
rect 25777 12727 25835 12733
rect 26326 12724 26332 12736
rect 26384 12724 26390 12776
rect 27709 12767 27767 12773
rect 27709 12733 27721 12767
rect 27755 12764 27767 12767
rect 27798 12764 27804 12776
rect 27755 12736 27804 12764
rect 27755 12733 27767 12736
rect 27709 12727 27767 12733
rect 27798 12724 27804 12736
rect 27856 12724 27862 12776
rect 8803 12668 9352 12696
rect 15013 12699 15071 12705
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 15286 12696 15292 12708
rect 15059 12668 15292 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 17236 12696 17264 12724
rect 17678 12696 17684 12708
rect 17236 12668 17684 12696
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 21361 12699 21419 12705
rect 21361 12665 21373 12699
rect 21407 12696 21419 12699
rect 21910 12696 21916 12708
rect 21407 12668 21916 12696
rect 21407 12665 21419 12668
rect 21361 12659 21419 12665
rect 21910 12656 21916 12668
rect 21968 12696 21974 12708
rect 21968 12668 25544 12696
rect 21968 12656 21974 12668
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11112 12600 12081 12628
rect 11112 12588 11118 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17589 12631 17647 12637
rect 17589 12628 17601 12631
rect 17276 12600 17601 12628
rect 17276 12588 17282 12600
rect 17589 12597 17601 12600
rect 17635 12628 17647 12631
rect 17862 12628 17868 12640
rect 17635 12600 17868 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 20901 12631 20959 12637
rect 20901 12597 20913 12631
rect 20947 12628 20959 12631
rect 20990 12628 20996 12640
rect 20947 12600 20996 12628
rect 20947 12597 20959 12600
rect 20901 12591 20959 12597
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 25409 12631 25467 12637
rect 25409 12628 25421 12631
rect 21692 12600 25421 12628
rect 21692 12588 21698 12600
rect 25409 12597 25421 12600
rect 25455 12597 25467 12631
rect 25516 12628 25544 12668
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 25516 12600 27537 12628
rect 25409 12591 25467 12597
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27525 12591 27583 12597
rect 38286 12588 38292 12640
rect 38344 12588 38350 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 10962 12384 10968 12436
rect 11020 12384 11026 12436
rect 14829 12427 14887 12433
rect 14829 12393 14841 12427
rect 14875 12424 14887 12427
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 14875 12396 16865 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 17862 12424 17868 12436
rect 16853 12387 16911 12393
rect 16960 12396 17868 12424
rect 13538 12316 13544 12368
rect 13596 12316 13602 12368
rect 14277 12359 14335 12365
rect 14277 12325 14289 12359
rect 14323 12325 14335 12359
rect 16117 12359 16175 12365
rect 16117 12356 16129 12359
rect 14277 12319 14335 12325
rect 14936 12328 16129 12356
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 8754 12288 8760 12300
rect 7892 12260 8760 12288
rect 7892 12248 7898 12260
rect 8754 12248 8760 12260
rect 8812 12288 8818 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 8812 12260 9413 12288
rect 8812 12248 8818 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 11698 12248 11704 12300
rect 11756 12248 11762 12300
rect 12710 12288 12716 12300
rect 12636 12260 12716 12288
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 10318 12220 10324 12232
rect 9723 12192 10324 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11716 12220 11744 12248
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11716 12192 11989 12220
rect 11977 12189 11989 12192
rect 12023 12220 12035 12223
rect 12158 12220 12164 12232
rect 12023 12192 12164 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 12636 12229 12664 12260
rect 12710 12248 12716 12260
rect 12768 12288 12774 12300
rect 14292 12288 14320 12319
rect 14936 12297 14964 12328
rect 16117 12325 16129 12328
rect 16163 12325 16175 12359
rect 16117 12319 16175 12325
rect 16758 12316 16764 12368
rect 16816 12356 16822 12368
rect 16960 12356 16988 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18049 12427 18107 12433
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 20901 12427 20959 12433
rect 18095 12396 19840 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18064 12356 18092 12387
rect 16816 12328 16988 12356
rect 17052 12328 18092 12356
rect 16816 12316 16822 12328
rect 12768 12260 14320 12288
rect 14921 12291 14979 12297
rect 12768 12248 12774 12260
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 15562 12288 15568 12300
rect 14921 12251 14979 12257
rect 15396 12260 15568 12288
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 15396 12229 15424 12260
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 16666 12288 16672 12300
rect 15703 12260 16672 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 17052 12297 17080 12328
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18288 12328 19012 12356
rect 18288 12316 18294 12328
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 14402 12223 14460 12229
rect 14402 12220 14414 12223
rect 13372 12192 14414 12220
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11701 12155 11759 12161
rect 11701 12152 11713 12155
rect 11204 12124 11713 12152
rect 11204 12112 11210 12124
rect 11701 12121 11713 12124
rect 11747 12152 11759 12155
rect 12342 12152 12348 12164
rect 11747 12124 12348 12152
rect 11747 12121 11759 12124
rect 11701 12115 11759 12121
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 12805 12155 12863 12161
rect 12805 12121 12817 12155
rect 12851 12152 12863 12155
rect 12894 12152 12900 12164
rect 12851 12124 12900 12152
rect 12851 12121 12863 12124
rect 12805 12115 12863 12121
rect 12894 12112 12900 12124
rect 12952 12112 12958 12164
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 13372 12161 13400 12192
rect 14402 12189 14414 12192
rect 14448 12189 14460 12223
rect 14402 12183 14460 12189
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15746 12220 15752 12232
rect 15519 12192 15752 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 15988 12192 16405 12220
rect 15988 12180 15994 12192
rect 16393 12189 16405 12192
rect 16439 12220 16451 12223
rect 17052 12220 17080 12251
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 17494 12288 17500 12300
rect 17184 12260 17500 12288
rect 17184 12248 17190 12260
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12288 17923 12291
rect 17954 12288 17960 12300
rect 17911 12260 17960 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 17954 12248 17960 12260
rect 18012 12288 18018 12300
rect 18874 12288 18880 12300
rect 18012 12260 18880 12288
rect 18012 12248 18018 12260
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 18984 12288 19012 12328
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19705 12359 19763 12365
rect 19705 12356 19717 12359
rect 19392 12328 19717 12356
rect 19392 12316 19398 12328
rect 19705 12325 19717 12328
rect 19751 12325 19763 12359
rect 19812 12356 19840 12396
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 21174 12424 21180 12436
rect 20947 12396 21180 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 25866 12384 25872 12436
rect 25924 12424 25930 12436
rect 25961 12427 26019 12433
rect 25961 12424 25973 12427
rect 25924 12396 25973 12424
rect 25924 12384 25930 12396
rect 25961 12393 25973 12396
rect 26007 12393 26019 12427
rect 25961 12387 26019 12393
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 27798 12424 27804 12436
rect 27755 12396 27804 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 27798 12384 27804 12396
rect 27856 12384 27862 12436
rect 29086 12384 29092 12436
rect 29144 12424 29150 12436
rect 38010 12424 38016 12436
rect 29144 12396 38016 12424
rect 29144 12384 29150 12396
rect 22094 12356 22100 12368
rect 19812 12328 22100 12356
rect 19705 12319 19763 12325
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 31386 12316 31392 12368
rect 31444 12356 31450 12368
rect 31444 12328 31754 12356
rect 31444 12316 31450 12328
rect 20622 12288 20628 12300
rect 18984 12260 20628 12288
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 21913 12291 21971 12297
rect 21913 12288 21925 12291
rect 21560 12260 21925 12288
rect 21560 12232 21588 12260
rect 21913 12257 21925 12260
rect 21959 12257 21971 12291
rect 21913 12251 21971 12257
rect 24578 12248 24584 12300
rect 24636 12288 24642 12300
rect 25314 12288 25320 12300
rect 24636 12260 25320 12288
rect 24636 12248 24642 12260
rect 25314 12248 25320 12260
rect 25372 12288 25378 12300
rect 25409 12291 25467 12297
rect 25409 12288 25421 12291
rect 25372 12260 25421 12288
rect 25372 12248 25378 12260
rect 25409 12257 25421 12260
rect 25455 12257 25467 12291
rect 25409 12251 25467 12257
rect 31297 12291 31355 12297
rect 31297 12257 31309 12291
rect 31343 12288 31355 12291
rect 31478 12288 31484 12300
rect 31343 12260 31484 12288
rect 31343 12257 31355 12260
rect 31297 12251 31355 12257
rect 31478 12248 31484 12260
rect 31536 12248 31542 12300
rect 31726 12288 31754 12328
rect 32766 12288 32772 12300
rect 31726 12260 32772 12288
rect 32766 12248 32772 12260
rect 32824 12248 32830 12300
rect 32968 12297 32996 12396
rect 38010 12384 38016 12396
rect 38068 12384 38074 12436
rect 32953 12291 33011 12297
rect 32953 12257 32965 12291
rect 32999 12257 33011 12291
rect 32953 12251 33011 12257
rect 35713 12291 35771 12297
rect 35713 12257 35725 12291
rect 35759 12288 35771 12291
rect 35802 12288 35808 12300
rect 35759 12260 35808 12288
rect 35759 12257 35771 12260
rect 35713 12251 35771 12257
rect 35802 12248 35808 12260
rect 35860 12248 35866 12300
rect 16439 12192 17080 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 17218 12180 17224 12232
rect 17276 12180 17282 12232
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 18141 12223 18199 12229
rect 17359 12192 17908 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 13228 12124 13369 12152
rect 13228 12112 13234 12124
rect 13357 12121 13369 12124
rect 13403 12121 13415 12155
rect 13357 12115 13415 12121
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 13587 12124 15884 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 11974 12044 11980 12096
rect 12032 12084 12038 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 12032 12056 12449 12084
rect 12032 12044 12038 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14240 12056 14473 12084
rect 14240 12044 14246 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 15654 12044 15660 12096
rect 15712 12044 15718 12096
rect 15856 12084 15884 12124
rect 16114 12112 16120 12164
rect 16172 12112 16178 12164
rect 17402 12152 17408 12164
rect 16224 12124 17408 12152
rect 16224 12084 16252 12124
rect 17402 12112 17408 12124
rect 17460 12112 17466 12164
rect 17880 12161 17908 12192
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 17865 12155 17923 12161
rect 17865 12121 17877 12155
rect 17911 12121 17923 12155
rect 17865 12115 17923 12121
rect 15856 12056 16252 12084
rect 16301 12087 16359 12093
rect 16301 12053 16313 12087
rect 16347 12084 16359 12087
rect 16666 12084 16672 12096
rect 16347 12056 16672 12084
rect 16347 12053 16359 12056
rect 16301 12047 16359 12053
rect 16666 12044 16672 12056
rect 16724 12084 16730 12096
rect 17678 12084 17684 12096
rect 16724 12056 17684 12084
rect 16724 12044 16730 12056
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17770 12044 17776 12096
rect 17828 12084 17834 12096
rect 18156 12084 18184 12183
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 18748 12192 19441 12220
rect 18748 12180 18754 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20254 12220 20260 12232
rect 19567 12192 20260 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20254 12180 20260 12192
rect 20312 12220 20318 12232
rect 20530 12220 20536 12232
rect 20312 12192 20536 12220
rect 20312 12180 20318 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21266 12180 21272 12232
rect 21324 12180 21330 12232
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12220 21419 12223
rect 21542 12220 21548 12232
rect 21407 12192 21548 12220
rect 21407 12189 21419 12192
rect 21361 12183 21419 12189
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12189 21879 12223
rect 21821 12183 21879 12189
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12152 19763 12155
rect 20162 12152 20168 12164
rect 19751 12124 20168 12152
rect 19751 12121 19763 12124
rect 19705 12115 19763 12121
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 17828 12056 18184 12084
rect 17828 12044 17834 12056
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 21836 12084 21864 12183
rect 22002 12180 22008 12232
rect 22060 12180 22066 12232
rect 27430 12180 27436 12232
rect 27488 12180 27494 12232
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 27709 12223 27767 12229
rect 27709 12220 27721 12223
rect 27672 12192 27721 12220
rect 27672 12180 27678 12192
rect 27709 12189 27721 12192
rect 27755 12189 27767 12223
rect 27709 12183 27767 12189
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 31570 12220 31576 12232
rect 31251 12192 31576 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 31570 12180 31576 12192
rect 31628 12220 31634 12232
rect 31628 12192 32812 12220
rect 31628 12180 31634 12192
rect 25685 12155 25743 12161
rect 25685 12121 25697 12155
rect 25731 12152 25743 12155
rect 25958 12152 25964 12164
rect 25731 12124 25964 12152
rect 25731 12121 25743 12124
rect 25685 12115 25743 12121
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 31113 12155 31171 12161
rect 27540 12124 31064 12152
rect 27540 12096 27568 12124
rect 19024 12056 21864 12084
rect 25501 12087 25559 12093
rect 19024 12044 19030 12056
rect 25501 12053 25513 12087
rect 25547 12084 25559 12087
rect 25590 12084 25596 12096
rect 25547 12056 25596 12084
rect 25547 12053 25559 12056
rect 25501 12047 25559 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 27522 12044 27528 12096
rect 27580 12044 27586 12096
rect 30558 12044 30564 12096
rect 30616 12084 30622 12096
rect 30745 12087 30803 12093
rect 30745 12084 30757 12087
rect 30616 12056 30757 12084
rect 30616 12044 30622 12056
rect 30745 12053 30757 12056
rect 30791 12053 30803 12087
rect 31036 12084 31064 12124
rect 31113 12121 31125 12155
rect 31159 12152 31171 12155
rect 31662 12152 31668 12164
rect 31159 12124 31668 12152
rect 31159 12121 31171 12124
rect 31113 12115 31171 12121
rect 31662 12112 31668 12124
rect 31720 12112 31726 12164
rect 32784 12096 32812 12192
rect 34606 12180 34612 12232
rect 34664 12220 34670 12232
rect 36909 12223 36967 12229
rect 36909 12220 36921 12223
rect 34664 12192 36921 12220
rect 34664 12180 34670 12192
rect 36909 12189 36921 12192
rect 36955 12189 36967 12223
rect 37918 12220 37924 12232
rect 36909 12183 36967 12189
rect 37108 12192 37924 12220
rect 32858 12112 32864 12164
rect 32916 12152 32922 12164
rect 35529 12155 35587 12161
rect 35529 12152 35541 12155
rect 32916 12124 35541 12152
rect 32916 12112 32922 12124
rect 35529 12121 35541 12124
rect 35575 12152 35587 12155
rect 37108 12152 37136 12192
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 35575 12124 37136 12152
rect 37176 12155 37234 12161
rect 35575 12121 35587 12124
rect 35529 12115 35587 12121
rect 37176 12121 37188 12155
rect 37222 12152 37234 12155
rect 37458 12152 37464 12164
rect 37222 12124 37464 12152
rect 37222 12121 37234 12124
rect 37176 12115 37234 12121
rect 37458 12112 37464 12124
rect 37516 12112 37522 12164
rect 32214 12084 32220 12096
rect 31036 12056 32220 12084
rect 30745 12047 30803 12053
rect 32214 12044 32220 12056
rect 32272 12044 32278 12096
rect 32306 12044 32312 12096
rect 32364 12044 32370 12096
rect 32674 12044 32680 12096
rect 32732 12044 32738 12096
rect 32766 12044 32772 12096
rect 32824 12044 32830 12096
rect 35069 12087 35127 12093
rect 35069 12053 35081 12087
rect 35115 12084 35127 12087
rect 35342 12084 35348 12096
rect 35115 12056 35348 12084
rect 35115 12053 35127 12056
rect 35069 12047 35127 12053
rect 35342 12044 35348 12056
rect 35400 12044 35406 12096
rect 35434 12044 35440 12096
rect 35492 12044 35498 12096
rect 37826 12044 37832 12096
rect 37884 12084 37890 12096
rect 38289 12087 38347 12093
rect 38289 12084 38301 12087
rect 37884 12056 38301 12084
rect 37884 12044 37890 12056
rect 38289 12053 38301 12056
rect 38335 12053 38347 12087
rect 38289 12047 38347 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 7834 11840 7840 11892
rect 7892 11840 7898 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11880 8999 11883
rect 9398 11880 9404 11892
rect 8987 11852 9404 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 15013 11883 15071 11889
rect 12308 11852 13032 11880
rect 12308 11840 12314 11852
rect 7852 11812 7880 11840
rect 7576 11784 7880 11812
rect 7576 11753 7604 11784
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 12342 11812 12348 11824
rect 10836 11784 11928 11812
rect 10836 11772 10842 11784
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7828 11747 7886 11753
rect 7828 11713 7840 11747
rect 7874 11744 7886 11747
rect 11054 11744 11060 11756
rect 7874 11716 11060 11744
rect 7874 11713 7886 11716
rect 7828 11707 7886 11713
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11900 11753 11928 11784
rect 12176 11784 12348 11812
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 12176 11753 12204 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 13004 11753 13032 11852
rect 15013 11849 15025 11883
rect 15059 11880 15071 11883
rect 15194 11880 15200 11892
rect 15059 11852 15200 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 21358 11880 21364 11892
rect 16540 11852 21364 11880
rect 16540 11840 16546 11852
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 16114 11812 16120 11824
rect 13320 11784 16120 11812
rect 13320 11772 13326 11784
rect 16114 11772 16120 11784
rect 16172 11812 16178 11824
rect 17126 11812 17132 11824
rect 16172 11784 17132 11812
rect 16172 11772 16178 11784
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 17681 11815 17739 11821
rect 17681 11781 17693 11815
rect 17727 11812 17739 11815
rect 17770 11812 17776 11824
rect 17727 11784 17776 11812
rect 17727 11781 17739 11784
rect 17681 11775 17739 11781
rect 17770 11772 17776 11784
rect 17828 11812 17834 11824
rect 17828 11784 19564 11812
rect 17828 11772 17834 11784
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12989 11747 13047 11753
rect 12299 11716 12940 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 10778 11636 10784 11688
rect 10836 11636 10842 11688
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11992 11676 12020 11704
rect 10919 11648 12020 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 12268 11608 12296 11707
rect 12710 11636 12716 11688
rect 12768 11636 12774 11688
rect 12912 11676 12940 11716
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 13998 11744 14004 11756
rect 13035 11716 14004 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15470 11744 15476 11756
rect 14967 11716 15476 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 15654 11744 15660 11756
rect 15528 11716 15660 11744
rect 15528 11704 15534 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 17310 11704 17316 11756
rect 17368 11704 17374 11756
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 18506 11704 18512 11756
rect 18564 11704 18570 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18616 11716 18705 11744
rect 15197 11679 15255 11685
rect 12912 11648 15148 11676
rect 11103 11580 12296 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 12894 11568 12900 11620
rect 12952 11608 12958 11620
rect 14553 11611 14611 11617
rect 14553 11608 14565 11611
rect 12952 11580 14565 11608
rect 12952 11568 12958 11580
rect 14553 11577 14565 11580
rect 14599 11577 14611 11611
rect 15120 11608 15148 11648
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15930 11676 15936 11688
rect 15243 11648 15936 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 18616 11676 18644 11716
rect 18693 11713 18705 11716
rect 18739 11744 18751 11747
rect 18739 11716 19196 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 16080 11648 18644 11676
rect 16080 11636 16086 11648
rect 15746 11608 15752 11620
rect 15120 11580 15752 11608
rect 14553 11571 14611 11577
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 18690 11568 18696 11620
rect 18748 11568 18754 11620
rect 19168 11608 19196 11716
rect 19334 11704 19340 11756
rect 19392 11704 19398 11756
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 19444 11620 19472 11707
rect 19536 11676 19564 11784
rect 19720 11753 19748 11852
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 24765 11883 24823 11889
rect 24765 11849 24777 11883
rect 24811 11849 24823 11883
rect 24765 11843 24823 11849
rect 23192 11815 23250 11821
rect 19687 11747 19748 11753
rect 19687 11713 19699 11747
rect 19733 11716 19748 11747
rect 19987 11784 20392 11812
rect 19987 11744 20015 11784
rect 19904 11716 20015 11744
rect 19733 11713 19745 11716
rect 19687 11707 19745 11713
rect 19904 11676 19932 11716
rect 20162 11704 20168 11756
rect 20220 11704 20226 11756
rect 20364 11753 20392 11784
rect 23192 11781 23204 11815
rect 23238 11812 23250 11815
rect 24780 11812 24808 11843
rect 25222 11840 25228 11892
rect 25280 11840 25286 11892
rect 32674 11840 32680 11892
rect 32732 11880 32738 11892
rect 33502 11880 33508 11892
rect 32732 11852 33508 11880
rect 32732 11840 32738 11852
rect 33502 11840 33508 11852
rect 33560 11880 33566 11892
rect 33689 11883 33747 11889
rect 33689 11880 33701 11883
rect 33560 11852 33701 11880
rect 33560 11840 33566 11852
rect 33689 11849 33701 11852
rect 33735 11849 33747 11883
rect 33689 11843 33747 11849
rect 34514 11840 34520 11892
rect 34572 11880 34578 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34572 11852 35173 11880
rect 34572 11840 34578 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 35161 11843 35219 11849
rect 37458 11840 37464 11892
rect 37516 11840 37522 11892
rect 37826 11840 37832 11892
rect 37884 11840 37890 11892
rect 37918 11840 37924 11892
rect 37976 11840 37982 11892
rect 23238 11784 24808 11812
rect 25133 11815 25191 11821
rect 23238 11781 23250 11784
rect 23192 11775 23250 11781
rect 25133 11781 25145 11815
rect 25179 11812 25191 11815
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 25179 11784 26157 11812
rect 25179 11781 25191 11784
rect 25133 11775 25191 11781
rect 26145 11781 26157 11784
rect 26191 11781 26203 11815
rect 26145 11775 26203 11781
rect 30392 11784 31754 11812
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 21726 11744 21732 11756
rect 20395 11716 21732 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 21726 11704 21732 11716
rect 21784 11704 21790 11756
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22612 11716 22937 11744
rect 22612 11704 22618 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 19536 11648 19932 11676
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 20036 11648 20637 11676
rect 20036 11636 20042 11648
rect 20625 11645 20637 11648
rect 20671 11676 20683 11679
rect 21634 11676 21640 11688
rect 20671 11648 21640 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 19168 11580 19334 11608
rect 10778 11500 10784 11552
rect 10836 11500 10842 11552
rect 11698 11500 11704 11552
rect 11756 11500 11762 11552
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12032 11512 12817 11540
rect 12032 11500 12038 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 18506 11540 18512 11552
rect 17368 11512 18512 11540
rect 17368 11500 17374 11512
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19150 11500 19156 11552
rect 19208 11500 19214 11552
rect 19306 11540 19334 11580
rect 19426 11568 19432 11620
rect 19484 11568 19490 11620
rect 19613 11611 19671 11617
rect 19613 11577 19625 11611
rect 19659 11608 19671 11611
rect 21266 11608 21272 11620
rect 19659 11580 21272 11608
rect 19659 11577 19671 11580
rect 19613 11571 19671 11577
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 24305 11611 24363 11617
rect 24305 11577 24317 11611
rect 24351 11608 24363 11611
rect 25148 11608 25176 11775
rect 30392 11756 30420 11784
rect 25866 11704 25872 11756
rect 25924 11744 25930 11756
rect 25961 11747 26019 11753
rect 25961 11744 25973 11747
rect 25924 11716 25973 11744
rect 25924 11704 25930 11716
rect 25961 11713 25973 11716
rect 26007 11713 26019 11747
rect 25961 11707 26019 11713
rect 26234 11704 26240 11756
rect 26292 11704 26298 11756
rect 30285 11747 30343 11753
rect 30285 11713 30297 11747
rect 30331 11744 30343 11747
rect 30374 11744 30380 11756
rect 30331 11716 30380 11744
rect 30331 11713 30343 11716
rect 30285 11707 30343 11713
rect 30374 11704 30380 11716
rect 30432 11704 30438 11756
rect 30558 11753 30564 11756
rect 30552 11744 30564 11753
rect 30519 11716 30564 11744
rect 30552 11707 30564 11716
rect 30558 11704 30564 11707
rect 30616 11704 30622 11756
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11676 25467 11679
rect 29086 11676 29092 11688
rect 25455 11648 29092 11676
rect 25455 11645 25467 11648
rect 25409 11639 25467 11645
rect 29086 11636 29092 11648
rect 29144 11636 29150 11688
rect 31726 11676 31754 11784
rect 32306 11772 32312 11824
rect 32364 11812 32370 11824
rect 32554 11815 32612 11821
rect 32554 11812 32566 11815
rect 32364 11784 32566 11812
rect 32364 11772 32370 11784
rect 32554 11781 32566 11784
rect 32600 11781 32612 11815
rect 32554 11775 32612 11781
rect 35253 11747 35311 11753
rect 35253 11713 35265 11747
rect 35299 11744 35311 11747
rect 35710 11744 35716 11756
rect 35299 11716 35716 11744
rect 35299 11713 35311 11716
rect 35253 11707 35311 11713
rect 35710 11704 35716 11716
rect 35768 11704 35774 11756
rect 35986 11704 35992 11756
rect 36044 11704 36050 11756
rect 36541 11747 36599 11753
rect 36541 11713 36553 11747
rect 36587 11744 36599 11747
rect 37844 11744 37872 11840
rect 36587 11716 37872 11744
rect 36587 11713 36599 11716
rect 36541 11707 36599 11713
rect 32309 11679 32367 11685
rect 32309 11676 32321 11679
rect 31726 11648 32321 11676
rect 32309 11645 32321 11648
rect 32355 11645 32367 11679
rect 32309 11639 32367 11645
rect 24351 11580 25176 11608
rect 24351 11577 24363 11580
rect 24305 11571 24363 11577
rect 25958 11568 25964 11620
rect 26016 11568 26022 11620
rect 19794 11540 19800 11552
rect 19306 11512 19800 11540
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 20496 11512 20545 11540
rect 20496 11500 20502 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 26234 11540 26240 11552
rect 20680 11512 26240 11540
rect 20680 11500 20686 11512
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 31662 11500 31668 11552
rect 31720 11500 31726 11552
rect 32324 11540 32352 11639
rect 35434 11636 35440 11688
rect 35492 11676 35498 11688
rect 35805 11679 35863 11685
rect 35805 11676 35817 11679
rect 35492 11648 35817 11676
rect 35492 11636 35498 11648
rect 35805 11645 35817 11648
rect 35851 11645 35863 11679
rect 35805 11639 35863 11645
rect 36262 11636 36268 11688
rect 36320 11636 36326 11688
rect 38010 11636 38016 11688
rect 38068 11636 38074 11688
rect 33042 11540 33048 11552
rect 32324 11512 33048 11540
rect 33042 11500 33048 11512
rect 33100 11500 33106 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 10318 11296 10324 11348
rect 10376 11296 10382 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 17954 11336 17960 11348
rect 12216 11308 17960 11336
rect 12216 11296 12222 11308
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 19886 11296 19892 11348
rect 19944 11336 19950 11348
rect 20438 11336 20444 11348
rect 19944 11308 20444 11336
rect 19944 11296 19950 11308
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 21910 11296 21916 11348
rect 21968 11296 21974 11348
rect 25682 11296 25688 11348
rect 25740 11296 25746 11348
rect 25866 11296 25872 11348
rect 25924 11296 25930 11348
rect 27614 11336 27620 11348
rect 26206 11308 27620 11336
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 16482 11268 16488 11280
rect 12400 11240 16488 11268
rect 12400 11228 12406 11240
rect 11698 11200 11704 11212
rect 10704 11172 11704 11200
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 10704 11141 10732 11172
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10468 11104 10517 11132
rect 10468 11092 10474 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 11882 11132 11888 11144
rect 11839 11104 11888 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 15764 11132 15792 11240
rect 16482 11228 16488 11240
rect 16540 11268 16546 11280
rect 16540 11240 17540 11268
rect 16540 11228 16546 11240
rect 17512 11209 17540 11240
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 21928 11268 21956 11296
rect 22278 11268 22284 11280
rect 18564 11240 21680 11268
rect 21928 11240 22284 11268
rect 18564 11228 18570 11240
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 16408 11172 17141 11200
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15764 11104 15853 11132
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 15933 11067 15991 11073
rect 14148 11036 15884 11064
rect 14148 11024 14154 11036
rect 11330 10956 11336 11008
rect 11388 10996 11394 11008
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11388 10968 11805 10996
rect 11388 10956 11394 10968
rect 11793 10965 11805 10968
rect 11839 10965 11851 10999
rect 15856 10996 15884 11036
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16298 11064 16304 11076
rect 15979 11036 16304 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 16408 10996 16436 11172
rect 17129 11169 17141 11172
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11200 17647 11203
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 17635 11172 18337 11200
rect 17635 11169 17647 11172
rect 17589 11163 17647 11169
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 16574 11092 16580 11144
rect 16632 11092 16638 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 17218 11132 17224 11144
rect 16715 11104 17224 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 17402 11092 17408 11144
rect 17460 11092 17466 11144
rect 17512 11132 17540 11163
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19024 11172 20024 11200
rect 19024 11160 19030 11172
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17512 11104 18245 11132
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 19518 11132 19524 11144
rect 18463 11104 19524 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 16592 11064 16620 11092
rect 19628 11064 19656 11095
rect 19794 11092 19800 11144
rect 19852 11092 19858 11144
rect 19886 11092 19892 11144
rect 19944 11092 19950 11144
rect 19996 11132 20024 11172
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 19996 11104 20361 11132
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 21508 11104 21557 11132
rect 21508 11092 21514 11104
rect 21545 11101 21557 11104
rect 21591 11101 21603 11135
rect 21652 11132 21680 11240
rect 22278 11228 22284 11240
rect 22336 11268 22342 11280
rect 22336 11240 22876 11268
rect 22336 11228 22342 11240
rect 21726 11160 21732 11212
rect 21784 11200 21790 11212
rect 22557 11203 22615 11209
rect 22557 11200 22569 11203
rect 21784 11172 22569 11200
rect 21784 11160 21790 11172
rect 22557 11169 22569 11172
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21652 11104 21833 11132
rect 21545 11095 21603 11101
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 22848 11141 22876 11240
rect 25774 11228 25780 11280
rect 25832 11268 25838 11280
rect 26206 11268 26234 11308
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 33134 11336 33140 11348
rect 31726 11308 33140 11336
rect 25832 11240 26234 11268
rect 25832 11228 25838 11240
rect 27890 11228 27896 11280
rect 27948 11268 27954 11280
rect 31726 11268 31754 11308
rect 33134 11296 33140 11308
rect 33192 11296 33198 11348
rect 35526 11296 35532 11348
rect 35584 11336 35590 11348
rect 36265 11339 36323 11345
rect 36265 11336 36277 11339
rect 35584 11308 36277 11336
rect 35584 11296 35590 11308
rect 36265 11305 36277 11308
rect 36311 11305 36323 11339
rect 36265 11299 36323 11305
rect 27948 11240 30512 11268
rect 27948 11228 27954 11240
rect 27614 11160 27620 11212
rect 27672 11200 27678 11212
rect 28905 11203 28963 11209
rect 28905 11200 28917 11203
rect 27672 11172 28917 11200
rect 27672 11160 27678 11172
rect 28905 11169 28917 11172
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 29086 11160 29092 11212
rect 29144 11160 29150 11212
rect 29362 11160 29368 11212
rect 29420 11200 29426 11212
rect 30484 11209 30512 11240
rect 30944 11240 31754 11268
rect 32493 11271 32551 11277
rect 29825 11203 29883 11209
rect 29825 11200 29837 11203
rect 29420 11172 29837 11200
rect 29420 11160 29426 11172
rect 29825 11169 29837 11172
rect 29871 11169 29883 11203
rect 29825 11163 29883 11169
rect 30469 11203 30527 11209
rect 30469 11169 30481 11203
rect 30515 11169 30527 11203
rect 30469 11163 30527 11169
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22244 11104 22753 11132
rect 22244 11092 22250 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 25424 11104 25636 11132
rect 21082 11064 21088 11076
rect 16592 11036 21088 11064
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 24854 11064 24860 11076
rect 21192 11036 24860 11064
rect 15856 10968 16436 10996
rect 16577 10999 16635 11005
rect 11793 10959 11851 10965
rect 16577 10965 16589 10999
rect 16623 10996 16635 10999
rect 17678 10996 17684 11008
rect 16623 10968 17684 10996
rect 16623 10965 16635 10968
rect 16577 10959 16635 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 21192 10996 21220 11036
rect 24854 11024 24860 11036
rect 24912 11064 24918 11076
rect 25424 11064 25452 11104
rect 24912 11036 25452 11064
rect 24912 11024 24918 11036
rect 25498 11024 25504 11076
rect 25556 11024 25562 11076
rect 25608 11064 25636 11104
rect 26510 11092 26516 11144
rect 26568 11132 26574 11144
rect 27706 11132 27712 11144
rect 26568 11104 27712 11132
rect 26568 11092 26574 11104
rect 27706 11092 27712 11104
rect 27764 11092 27770 11144
rect 29638 11092 29644 11144
rect 29696 11132 29702 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29696 11104 29745 11132
rect 29696 11092 29702 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 30653 11135 30711 11141
rect 30653 11101 30665 11135
rect 30699 11132 30711 11135
rect 30944 11132 30972 11240
rect 32493 11237 32505 11271
rect 32539 11268 32551 11271
rect 33410 11268 33416 11280
rect 32539 11240 33416 11268
rect 32539 11237 32551 11240
rect 32493 11231 32551 11237
rect 33410 11228 33416 11240
rect 33468 11228 33474 11280
rect 31662 11160 31668 11212
rect 31720 11200 31726 11212
rect 32953 11203 33011 11209
rect 32953 11200 32965 11203
rect 31720 11172 32965 11200
rect 31720 11160 31726 11172
rect 32953 11169 32965 11172
rect 32999 11169 33011 11203
rect 32953 11163 33011 11169
rect 34606 11160 34612 11212
rect 34664 11200 34670 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34664 11172 34897 11200
rect 34664 11160 34670 11172
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 34885 11163 34943 11169
rect 30699 11104 30972 11132
rect 31021 11135 31079 11141
rect 30699 11101 30711 11104
rect 30653 11095 30711 11101
rect 31021 11101 31033 11135
rect 31067 11101 31079 11135
rect 31021 11095 31079 11101
rect 31573 11135 31631 11141
rect 31573 11101 31585 11135
rect 31619 11101 31631 11135
rect 31573 11095 31631 11101
rect 25701 11067 25759 11073
rect 25701 11064 25713 11067
rect 25608 11036 25713 11064
rect 25701 11033 25713 11036
rect 25747 11033 25759 11067
rect 25701 11027 25759 11033
rect 26780 11067 26838 11073
rect 26780 11033 26792 11067
rect 26826 11064 26838 11067
rect 27154 11064 27160 11076
rect 26826 11036 27160 11064
rect 26826 11033 26838 11036
rect 26780 11027 26838 11033
rect 27154 11024 27160 11036
rect 27212 11024 27218 11076
rect 28813 11067 28871 11073
rect 28813 11033 28825 11067
rect 28859 11064 28871 11067
rect 29914 11064 29920 11076
rect 28859 11036 29920 11064
rect 28859 11033 28871 11036
rect 28813 11027 28871 11033
rect 29914 11024 29920 11036
rect 29972 11064 29978 11076
rect 31036 11064 31064 11095
rect 29972 11036 31064 11064
rect 29972 11024 29978 11036
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 31588 11064 31616 11095
rect 32214 11092 32220 11144
rect 32272 11092 32278 11144
rect 33134 11092 33140 11144
rect 33192 11092 33198 11144
rect 33413 11135 33471 11141
rect 33413 11101 33425 11135
rect 33459 11101 33471 11135
rect 33413 11095 33471 11101
rect 33428 11064 33456 11095
rect 33502 11092 33508 11144
rect 33560 11092 33566 11144
rect 34900 11132 34928 11163
rect 36817 11135 36875 11141
rect 36817 11132 36829 11135
rect 34900 11104 36829 11132
rect 36817 11101 36829 11104
rect 36863 11101 36875 11135
rect 36817 11095 36875 11101
rect 35152 11067 35210 11073
rect 31352 11036 35112 11064
rect 31352 11024 31358 11036
rect 17920 10968 21220 10996
rect 17920 10956 17926 10968
rect 22094 10956 22100 11008
rect 22152 10956 22158 11008
rect 22370 10956 22376 11008
rect 22428 10996 22434 11008
rect 22557 10999 22615 11005
rect 22557 10996 22569 10999
rect 22428 10968 22569 10996
rect 22428 10956 22434 10968
rect 22557 10965 22569 10968
rect 22603 10965 22615 10999
rect 22557 10959 22615 10965
rect 28442 10956 28448 11008
rect 28500 10956 28506 11008
rect 31478 10956 31484 11008
rect 31536 10996 31542 11008
rect 34514 10996 34520 11008
rect 31536 10968 34520 10996
rect 31536 10956 31542 10968
rect 34514 10956 34520 10968
rect 34572 10956 34578 11008
rect 35084 10996 35112 11036
rect 35152 11033 35164 11067
rect 35198 11064 35210 11067
rect 35342 11064 35348 11076
rect 35198 11036 35348 11064
rect 35198 11033 35210 11036
rect 35152 11027 35210 11033
rect 35342 11024 35348 11036
rect 35400 11024 35406 11076
rect 36262 11064 36268 11076
rect 35452 11036 36268 11064
rect 35452 10996 35480 11036
rect 36262 11024 36268 11036
rect 36320 11024 36326 11076
rect 37084 11067 37142 11073
rect 37084 11033 37096 11067
rect 37130 11064 37142 11067
rect 37458 11064 37464 11076
rect 37130 11036 37464 11064
rect 37130 11033 37142 11036
rect 37084 11027 37142 11033
rect 37458 11024 37464 11036
rect 37516 11024 37522 11076
rect 35084 10968 35480 10996
rect 38194 10956 38200 11008
rect 38252 10956 38258 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 10134 10752 10140 10804
rect 10192 10752 10198 10804
rect 17221 10795 17279 10801
rect 17221 10761 17233 10795
rect 17267 10792 17279 10795
rect 17310 10792 17316 10804
rect 17267 10764 17316 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17678 10752 17684 10804
rect 17736 10752 17742 10804
rect 21177 10795 21235 10801
rect 21177 10761 21189 10795
rect 21223 10792 21235 10795
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21223 10764 22017 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 26878 10792 26884 10804
rect 22005 10755 22063 10761
rect 22112 10764 26884 10792
rect 14734 10724 14740 10736
rect 13648 10696 14740 10724
rect 13648 10668 13676 10696
rect 14734 10684 14740 10696
rect 14792 10724 14798 10736
rect 15105 10727 15163 10733
rect 15105 10724 15117 10727
rect 14792 10696 15117 10724
rect 14792 10684 14798 10696
rect 15105 10693 15117 10696
rect 15151 10693 15163 10727
rect 15105 10687 15163 10693
rect 17589 10727 17647 10733
rect 17589 10693 17601 10727
rect 17635 10724 17647 10727
rect 17770 10724 17776 10736
rect 17635 10696 17776 10724
rect 17635 10693 17647 10696
rect 17589 10687 17647 10693
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18138 10684 18144 10736
rect 18196 10724 18202 10736
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 18196 10696 18889 10724
rect 18196 10684 18202 10696
rect 18877 10693 18889 10696
rect 18923 10724 18935 10727
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 18923 10696 21097 10724
rect 18923 10693 18935 10696
rect 18877 10687 18935 10693
rect 21085 10693 21097 10696
rect 21131 10724 21143 10727
rect 22112 10724 22140 10764
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 27154 10752 27160 10804
rect 27212 10752 27218 10804
rect 27525 10795 27583 10801
rect 27525 10761 27537 10795
rect 27571 10792 27583 10795
rect 27890 10792 27896 10804
rect 27571 10764 27896 10792
rect 27571 10761 27583 10764
rect 27525 10755 27583 10761
rect 27890 10752 27896 10764
rect 27948 10752 27954 10804
rect 29733 10795 29791 10801
rect 29733 10761 29745 10795
rect 29779 10792 29791 10795
rect 29914 10792 29920 10804
rect 29779 10764 29920 10792
rect 29779 10761 29791 10764
rect 29733 10755 29791 10761
rect 29914 10752 29920 10764
rect 29972 10752 29978 10804
rect 37458 10752 37464 10804
rect 37516 10752 37522 10804
rect 21131 10696 22140 10724
rect 21131 10693 21143 10696
rect 21085 10687 21143 10693
rect 22278 10684 22284 10736
rect 22336 10684 22342 10736
rect 22370 10684 22376 10736
rect 22428 10684 22434 10736
rect 26510 10724 26516 10736
rect 24412 10696 26516 10724
rect 8754 10616 8760 10668
rect 8812 10616 8818 10668
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14182 10656 14188 10668
rect 13863 10628 14188 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 22186 10616 22192 10668
rect 22244 10616 22250 10668
rect 24412 10665 24440 10696
rect 26510 10684 26516 10696
rect 26568 10684 26574 10736
rect 27614 10684 27620 10736
rect 27672 10684 27678 10736
rect 27706 10684 27712 10736
rect 27764 10684 27770 10736
rect 28442 10684 28448 10736
rect 28500 10724 28506 10736
rect 28598 10727 28656 10733
rect 28598 10724 28610 10727
rect 28500 10696 28610 10724
rect 28500 10684 28506 10696
rect 28598 10693 28610 10696
rect 28644 10693 28656 10727
rect 37642 10724 37648 10736
rect 28598 10687 28656 10693
rect 34256 10696 37648 10724
rect 24670 10665 24676 10668
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24664 10619 24676 10665
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 10318 10588 10324 10600
rect 9079 10560 10324 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 15654 10548 15660 10600
rect 15712 10548 15718 10600
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 17911 10560 18429 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 21358 10548 21364 10600
rect 21416 10548 21422 10600
rect 22094 10548 22100 10600
rect 22152 10588 22158 10600
rect 22572 10588 22600 10619
rect 24670 10616 24676 10619
rect 24728 10616 24734 10668
rect 26142 10616 26148 10668
rect 26200 10656 26206 10668
rect 27724 10656 27752 10684
rect 28353 10659 28411 10665
rect 28353 10656 28365 10659
rect 26200 10616 26234 10656
rect 27724 10628 28365 10656
rect 28353 10625 28365 10628
rect 28399 10625 28411 10659
rect 28353 10619 28411 10625
rect 34146 10616 34152 10668
rect 34204 10616 34210 10668
rect 22152 10560 22600 10588
rect 22152 10548 22158 10560
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18601 10523 18659 10529
rect 18601 10520 18613 10523
rect 17828 10492 18613 10520
rect 17828 10480 17834 10492
rect 18601 10489 18613 10492
rect 18647 10520 18659 10523
rect 22646 10520 22652 10532
rect 18647 10492 22652 10520
rect 18647 10489 18659 10492
rect 18601 10483 18659 10489
rect 22646 10480 22652 10492
rect 22704 10480 22710 10532
rect 13446 10412 13452 10464
rect 13504 10412 13510 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13596 10424 13645 10452
rect 13596 10412 13602 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 20898 10452 20904 10464
rect 20763 10424 20904 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 25498 10452 25504 10464
rect 25188 10424 25504 10452
rect 25188 10412 25194 10424
rect 25498 10412 25504 10424
rect 25556 10452 25562 10464
rect 25777 10455 25835 10461
rect 25777 10452 25789 10455
rect 25556 10424 25789 10452
rect 25556 10412 25562 10424
rect 25777 10421 25789 10424
rect 25823 10421 25835 10455
rect 26206 10452 26234 10616
rect 27798 10548 27804 10600
rect 27856 10548 27862 10600
rect 33962 10588 33968 10600
rect 31726 10560 33968 10588
rect 31726 10452 31754 10560
rect 33962 10548 33968 10560
rect 34020 10588 34026 10600
rect 34256 10597 34284 10696
rect 37642 10684 37648 10696
rect 37700 10724 37706 10736
rect 37921 10727 37979 10733
rect 37921 10724 37933 10727
rect 37700 10696 37933 10724
rect 37700 10684 37706 10696
rect 37921 10693 37933 10696
rect 37967 10693 37979 10727
rect 37921 10687 37979 10693
rect 37366 10616 37372 10668
rect 37424 10656 37430 10668
rect 37829 10659 37887 10665
rect 37829 10656 37841 10659
rect 37424 10628 37841 10656
rect 37424 10616 37430 10628
rect 37829 10625 37841 10628
rect 37875 10656 37887 10659
rect 38194 10656 38200 10668
rect 37875 10628 38200 10656
rect 37875 10625 37887 10628
rect 37829 10619 37887 10625
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 34241 10591 34299 10597
rect 34241 10588 34253 10591
rect 34020 10560 34253 10588
rect 34020 10548 34026 10560
rect 34241 10557 34253 10560
rect 34287 10557 34299 10591
rect 34241 10551 34299 10557
rect 34425 10591 34483 10597
rect 34425 10557 34437 10591
rect 34471 10588 34483 10591
rect 34514 10588 34520 10600
rect 34471 10560 34520 10588
rect 34471 10557 34483 10560
rect 34425 10551 34483 10557
rect 34514 10548 34520 10560
rect 34572 10588 34578 10600
rect 35802 10588 35808 10600
rect 34572 10560 35808 10588
rect 34572 10548 34578 10560
rect 35802 10548 35808 10560
rect 35860 10548 35866 10600
rect 38010 10548 38016 10600
rect 38068 10548 38074 10600
rect 26206 10424 31754 10452
rect 25777 10415 25835 10421
rect 33778 10412 33784 10464
rect 33836 10412 33842 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10318 10208 10324 10260
rect 10376 10208 10382 10260
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 11149 10251 11207 10257
rect 11149 10248 11161 10251
rect 10928 10220 11161 10248
rect 10928 10208 10934 10220
rect 11149 10217 11161 10220
rect 11195 10217 11207 10251
rect 11149 10211 11207 10217
rect 17402 10208 17408 10260
rect 17460 10248 17466 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 17460 10220 17509 10248
rect 17460 10208 17466 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 21821 10251 21879 10257
rect 17736 10220 19564 10248
rect 17736 10208 17742 10220
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 10888 10112 10916 10208
rect 14182 10140 14188 10192
rect 14240 10180 14246 10192
rect 14829 10183 14887 10189
rect 14829 10180 14841 10183
rect 14240 10152 14841 10180
rect 14240 10140 14246 10152
rect 14829 10149 14841 10152
rect 14875 10149 14887 10183
rect 19426 10180 19432 10192
rect 14829 10143 14887 10149
rect 15488 10152 19432 10180
rect 10735 10084 10916 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 12066 10112 12072 10124
rect 11112 10084 12072 10112
rect 11112 10072 11118 10084
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 15488 10121 15516 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 19536 10180 19564 10220
rect 21821 10217 21833 10251
rect 21867 10248 21879 10251
rect 22186 10248 22192 10260
rect 21867 10220 22192 10248
rect 21867 10217 21879 10220
rect 21821 10211 21879 10217
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 24765 10251 24823 10257
rect 24765 10248 24777 10251
rect 24728 10220 24777 10248
rect 24728 10208 24734 10220
rect 24765 10217 24777 10220
rect 24811 10217 24823 10251
rect 24765 10211 24823 10217
rect 31757 10251 31815 10257
rect 31757 10217 31769 10251
rect 31803 10248 31815 10251
rect 32214 10248 32220 10260
rect 31803 10220 32220 10248
rect 31803 10217 31815 10220
rect 31757 10211 31815 10217
rect 32214 10208 32220 10220
rect 32272 10208 32278 10260
rect 19536 10152 21956 10180
rect 15473 10115 15531 10121
rect 15473 10081 15485 10115
rect 15519 10081 15531 10115
rect 15473 10075 15531 10081
rect 16040 10084 16574 10112
rect 16040 10056 16068 10084
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11790 10044 11796 10056
rect 11655 10016 11796 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 11900 10016 12357 10044
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11900 9976 11928 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14826 10044 14832 10056
rect 13771 10016 14832 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10044 15255 10047
rect 15286 10044 15292 10056
rect 15243 10016 15292 10044
rect 15243 10013 15255 10016
rect 15197 10007 15255 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 11296 9948 11928 9976
rect 15304 9976 15332 10004
rect 16117 9979 16175 9985
rect 16117 9976 16129 9979
rect 15304 9948 16129 9976
rect 11296 9936 11302 9948
rect 16117 9945 16129 9948
rect 16163 9945 16175 9979
rect 16117 9939 16175 9945
rect 11514 9868 11520 9920
rect 11572 9868 11578 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 15252 9880 15301 9908
rect 15252 9868 15258 9880
rect 15289 9877 15301 9880
rect 15335 9908 15347 9911
rect 16224 9908 16252 10007
rect 16546 9976 16574 10084
rect 17678 10072 17684 10124
rect 17736 10072 17742 10124
rect 17770 10072 17776 10124
rect 17828 10072 17834 10124
rect 18138 10072 18144 10124
rect 18196 10072 18202 10124
rect 20070 10112 20076 10124
rect 19352 10084 20076 10112
rect 19352 9976 19380 10084
rect 20070 10072 20076 10084
rect 20128 10112 20134 10124
rect 20349 10115 20407 10121
rect 20128 10084 20300 10112
rect 20128 10072 20134 10084
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20272 10044 20300 10084
rect 20349 10081 20361 10115
rect 20395 10112 20407 10115
rect 20714 10112 20720 10124
rect 20395 10084 20720 10112
rect 20395 10081 20407 10084
rect 20349 10075 20407 10081
rect 20714 10072 20720 10084
rect 20772 10112 20778 10124
rect 20772 10084 21128 10112
rect 20772 10072 20778 10084
rect 20441 10047 20499 10053
rect 20441 10044 20453 10047
rect 20272 10016 20453 10044
rect 20165 10007 20223 10013
rect 20441 10013 20453 10016
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 16546 9948 19380 9976
rect 20180 9976 20208 10007
rect 20898 10004 20904 10056
rect 20956 10004 20962 10056
rect 21100 10053 21128 10084
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10013 21143 10047
rect 21085 10007 21143 10013
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21928 10053 21956 10152
rect 34146 10140 34152 10192
rect 34204 10180 34210 10192
rect 34333 10183 34391 10189
rect 34333 10180 34345 10183
rect 34204 10152 34345 10180
rect 34204 10140 34210 10152
rect 34333 10149 34345 10152
rect 34379 10149 34391 10183
rect 34333 10143 34391 10149
rect 25222 10072 25228 10124
rect 25280 10072 25286 10124
rect 25409 10115 25467 10121
rect 25409 10081 25421 10115
rect 25455 10112 25467 10115
rect 27798 10112 27804 10124
rect 25455 10084 27804 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 27798 10072 27804 10084
rect 27856 10072 27862 10124
rect 34348 10112 34376 10143
rect 34422 10140 34428 10192
rect 34480 10180 34486 10192
rect 35161 10183 35219 10189
rect 35161 10180 35173 10183
rect 34480 10152 35173 10180
rect 34480 10140 34486 10152
rect 35161 10149 35173 10152
rect 35207 10149 35219 10183
rect 35161 10143 35219 10149
rect 35805 10115 35863 10121
rect 35805 10112 35817 10115
rect 34348 10084 35817 10112
rect 35805 10081 35817 10084
rect 35851 10081 35863 10115
rect 35805 10075 35863 10081
rect 36262 10072 36268 10124
rect 36320 10072 36326 10124
rect 37366 10112 37372 10124
rect 36556 10084 37372 10112
rect 21729 10047 21787 10053
rect 21729 10044 21741 10047
rect 21508 10016 21741 10044
rect 21508 10004 21514 10016
rect 21729 10013 21741 10016
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 25130 10004 25136 10056
rect 25188 10004 25194 10056
rect 32030 10004 32036 10056
rect 32088 10004 32094 10056
rect 32122 10004 32128 10056
rect 32180 10004 32186 10056
rect 32217 10047 32275 10053
rect 32217 10013 32229 10047
rect 32263 10013 32275 10047
rect 32217 10007 32275 10013
rect 32401 10047 32459 10053
rect 32401 10013 32413 10047
rect 32447 10013 32459 10047
rect 32401 10007 32459 10013
rect 32953 10047 33011 10053
rect 32953 10013 32965 10047
rect 32999 10044 33011 10047
rect 33042 10044 33048 10056
rect 32999 10016 33048 10044
rect 32999 10013 33011 10016
rect 32953 10007 33011 10013
rect 20916 9976 20944 10004
rect 20180 9948 20944 9976
rect 15335 9880 16252 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 19978 9868 19984 9920
rect 20036 9868 20042 9920
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20956 9880 21005 9908
rect 20956 9868 20962 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 32232 9908 32260 10007
rect 32416 9976 32444 10007
rect 33042 10004 33048 10016
rect 33100 10004 33106 10056
rect 33220 10047 33278 10053
rect 33220 10013 33232 10047
rect 33266 10044 33278 10047
rect 33778 10044 33784 10056
rect 33266 10016 33784 10044
rect 33266 10013 33278 10016
rect 33220 10007 33278 10013
rect 33778 10004 33784 10016
rect 33836 10004 33842 10056
rect 35253 10047 35311 10053
rect 35253 10013 35265 10047
rect 35299 10044 35311 10047
rect 35434 10044 35440 10056
rect 35299 10016 35440 10044
rect 35299 10013 35311 10016
rect 35253 10007 35311 10013
rect 35434 10004 35440 10016
rect 35492 10004 35498 10056
rect 35986 10004 35992 10056
rect 36044 10044 36050 10056
rect 36354 10044 36360 10056
rect 36044 10016 36360 10044
rect 36044 10004 36050 10016
rect 36354 10004 36360 10016
rect 36412 10004 36418 10056
rect 36556 10053 36584 10084
rect 37366 10072 37372 10084
rect 37424 10072 37430 10124
rect 38105 10115 38163 10121
rect 38105 10081 38117 10115
rect 38151 10112 38163 10115
rect 39022 10112 39028 10124
rect 38151 10084 39028 10112
rect 38151 10081 38163 10084
rect 38105 10075 38163 10081
rect 39022 10072 39028 10084
rect 39080 10072 39086 10124
rect 36541 10047 36599 10053
rect 36541 10013 36553 10047
rect 36587 10013 36599 10047
rect 36541 10007 36599 10013
rect 37826 10004 37832 10056
rect 37884 10004 37890 10056
rect 33870 9976 33876 9988
rect 32416 9948 33876 9976
rect 33870 9936 33876 9948
rect 33928 9936 33934 9988
rect 32950 9908 32956 9920
rect 32232 9880 32956 9908
rect 20993 9871 21051 9877
rect 32950 9868 32956 9880
rect 33008 9868 33014 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 10870 9664 10876 9716
rect 10928 9664 10934 9716
rect 13357 9707 13415 9713
rect 13357 9673 13369 9707
rect 13403 9704 13415 9707
rect 13446 9704 13452 9716
rect 13403 9676 13452 9704
rect 13403 9673 13415 9676
rect 13357 9667 13415 9673
rect 10410 9596 10416 9648
rect 10468 9596 10474 9648
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11388 9608 11989 9636
rect 11388 9596 11394 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 13372 9636 13400 9667
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 15286 9664 15292 9716
rect 15344 9664 15350 9716
rect 20714 9664 20720 9716
rect 20772 9664 20778 9716
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 26510 9704 26516 9716
rect 22612 9676 26516 9704
rect 22612 9664 22618 9676
rect 26510 9664 26516 9676
rect 26568 9664 26574 9716
rect 27798 9664 27804 9716
rect 27856 9704 27862 9716
rect 28442 9704 28448 9716
rect 27856 9676 28448 9704
rect 27856 9664 27862 9676
rect 28442 9664 28448 9676
rect 28500 9704 28506 9716
rect 28500 9676 29776 9704
rect 28500 9664 28506 9676
rect 11977 9599 12035 9605
rect 12544 9608 13400 9636
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10560 9540 10701 9568
rect 10560 9528 10566 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10704 9432 10732 9531
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11238 9568 11244 9580
rect 11195 9540 11244 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11572 9540 11713 9568
rect 11572 9528 11578 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11716 9500 11744 9531
rect 11790 9528 11796 9580
rect 11848 9528 11854 9580
rect 12544 9500 12572 9608
rect 13998 9596 14004 9648
rect 14056 9596 14062 9648
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15381 9639 15439 9645
rect 15381 9636 15393 9639
rect 15252 9608 15393 9636
rect 15252 9596 15258 9608
rect 15381 9605 15393 9608
rect 15427 9636 15439 9639
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 15427 9608 16574 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 12943 9540 13829 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 14016 9568 14044 9596
rect 15470 9568 15476 9580
rect 14016 9540 15476 9568
rect 13817 9531 13875 9537
rect 15470 9528 15476 9540
rect 15528 9568 15534 9580
rect 16022 9568 16028 9580
rect 15528 9540 16028 9568
rect 15528 9528 15534 9540
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 16546 9568 16574 9608
rect 17052 9608 19073 9636
rect 17052 9577 17080 9608
rect 19061 9605 19073 9608
rect 19107 9636 19119 9639
rect 21177 9639 21235 9645
rect 21177 9636 21189 9639
rect 19107 9608 21189 9636
rect 19107 9605 19119 9608
rect 19061 9599 19119 9605
rect 21177 9605 21189 9608
rect 21223 9636 21235 9639
rect 22462 9636 22468 9648
rect 21223 9608 22468 9636
rect 21223 9605 21235 9608
rect 21177 9599 21235 9605
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 24857 9639 24915 9645
rect 24857 9605 24869 9639
rect 24903 9636 24915 9639
rect 25222 9636 25228 9648
rect 24903 9608 25228 9636
rect 24903 9605 24915 9608
rect 24857 9599 24915 9605
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 25590 9596 25596 9648
rect 25648 9596 25654 9648
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16546 9540 17049 9568
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 19153 9571 19211 9577
rect 19153 9568 19165 9571
rect 17644 9540 19165 9568
rect 17644 9528 17650 9540
rect 19153 9537 19165 9540
rect 19199 9568 19211 9571
rect 21082 9568 21088 9580
rect 19199 9540 21088 9568
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 22824 9571 22882 9577
rect 22824 9537 22836 9571
rect 22870 9568 22882 9571
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 22870 9540 24440 9568
rect 22870 9537 22882 9540
rect 22824 9531 22882 9537
rect 11716 9472 12572 9500
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 17770 9500 17776 9512
rect 15611 9472 17776 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 11701 9435 11759 9441
rect 11701 9432 11713 9435
rect 10704 9404 11713 9432
rect 11701 9401 11713 9404
rect 11747 9401 11759 9435
rect 13004 9432 13032 9463
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 21361 9503 21419 9509
rect 21361 9469 21373 9503
rect 21407 9500 21419 9503
rect 21450 9500 21456 9512
rect 21407 9472 21456 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 13538 9432 13544 9444
rect 13004 9404 13544 9432
rect 11701 9395 11759 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 18984 9432 19012 9463
rect 21450 9460 21456 9472
rect 21508 9460 21514 9512
rect 20530 9432 20536 9444
rect 18984 9404 20536 9432
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 24412 9441 24440 9540
rect 24688 9540 24777 9568
rect 24397 9435 24455 9441
rect 24397 9401 24409 9435
rect 24443 9401 24455 9435
rect 24397 9395 24455 9401
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11146 9364 11152 9376
rect 11103 9336 11152 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 12713 9367 12771 9373
rect 12713 9333 12725 9367
rect 12759 9364 12771 9367
rect 12802 9364 12808 9376
rect 12759 9336 12808 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14608 9336 14933 9364
rect 14608 9324 14614 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16540 9336 16957 9364
rect 16540 9324 16546 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 19521 9367 19579 9373
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 19794 9364 19800 9376
rect 19567 9336 19800 9364
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 23937 9367 23995 9373
rect 23937 9333 23949 9367
rect 23983 9364 23995 9367
rect 24688 9364 24716 9540
rect 24765 9537 24777 9540
rect 24811 9568 24823 9571
rect 25869 9571 25927 9577
rect 25869 9568 25881 9571
rect 24811 9540 25881 9568
rect 24811 9537 24823 9540
rect 24765 9531 24823 9537
rect 25869 9537 25881 9540
rect 25915 9537 25927 9571
rect 26528 9568 26556 9664
rect 29196 9608 29500 9636
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26528 9540 27169 9568
rect 25869 9531 25927 9537
rect 27157 9537 27169 9540
rect 27203 9568 27215 9571
rect 27246 9568 27252 9580
rect 27203 9540 27252 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 27246 9528 27252 9540
rect 27304 9528 27310 9580
rect 27430 9577 27436 9580
rect 27424 9531 27436 9577
rect 27430 9528 27436 9531
rect 27488 9528 27494 9580
rect 28994 9528 29000 9580
rect 29052 9528 29058 9580
rect 29196 9577 29224 9608
rect 29181 9571 29239 9577
rect 29181 9537 29193 9571
rect 29227 9537 29239 9571
rect 29181 9531 29239 9537
rect 29270 9528 29276 9580
rect 29328 9528 29334 9580
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 25038 9460 25044 9512
rect 25096 9460 25102 9512
rect 25314 9460 25320 9512
rect 25372 9500 25378 9512
rect 25593 9503 25651 9509
rect 25593 9500 25605 9503
rect 25372 9472 25605 9500
rect 25372 9460 25378 9472
rect 25593 9469 25605 9472
rect 25639 9469 25651 9503
rect 29380 9500 29408 9531
rect 25593 9463 25651 9469
rect 28552 9472 29408 9500
rect 28552 9376 28580 9472
rect 23983 9336 24716 9364
rect 25777 9367 25835 9373
rect 23983 9333 23995 9336
rect 23937 9327 23995 9333
rect 25777 9333 25789 9367
rect 25823 9364 25835 9367
rect 26234 9364 26240 9376
rect 25823 9336 26240 9364
rect 25823 9333 25835 9336
rect 25777 9327 25835 9333
rect 26234 9324 26240 9336
rect 26292 9364 26298 9376
rect 26878 9364 26884 9376
rect 26292 9336 26884 9364
rect 26292 9324 26298 9336
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 28534 9324 28540 9376
rect 28592 9324 28598 9376
rect 29472 9364 29500 9608
rect 29638 9596 29644 9648
rect 29696 9596 29702 9648
rect 29748 9636 29776 9676
rect 32030 9664 32036 9716
rect 32088 9704 32094 9716
rect 32677 9707 32735 9713
rect 32677 9704 32689 9707
rect 32088 9676 32689 9704
rect 32088 9664 32094 9676
rect 32677 9673 32689 9676
rect 32723 9673 32735 9707
rect 32677 9667 32735 9673
rect 34977 9707 35035 9713
rect 34977 9673 34989 9707
rect 35023 9673 35035 9707
rect 34977 9667 35035 9673
rect 30101 9639 30159 9645
rect 30101 9636 30113 9639
rect 29748 9608 30113 9636
rect 30101 9605 30113 9608
rect 30147 9636 30159 9639
rect 31478 9636 31484 9648
rect 30147 9608 31484 9636
rect 30147 9605 30159 9608
rect 30101 9599 30159 9605
rect 31478 9596 31484 9608
rect 31536 9596 31542 9648
rect 33134 9596 33140 9648
rect 33192 9636 33198 9648
rect 34992 9636 35020 9667
rect 36354 9636 36360 9648
rect 33192 9608 36360 9636
rect 33192 9596 33198 9608
rect 36354 9596 36360 9608
rect 36412 9596 36418 9648
rect 38105 9639 38163 9645
rect 38105 9605 38117 9639
rect 38151 9636 38163 9639
rect 39022 9636 39028 9648
rect 38151 9608 39028 9636
rect 38151 9605 38163 9608
rect 38105 9599 38163 9605
rect 39022 9596 39028 9608
rect 39080 9596 39086 9648
rect 30190 9528 30196 9580
rect 30248 9568 30254 9580
rect 30561 9571 30619 9577
rect 30561 9568 30573 9571
rect 30248 9540 30573 9568
rect 30248 9528 30254 9540
rect 30561 9537 30573 9540
rect 30607 9537 30619 9571
rect 30561 9531 30619 9537
rect 30653 9571 30711 9577
rect 30653 9537 30665 9571
rect 30699 9568 30711 9571
rect 33152 9568 33180 9596
rect 30699 9540 33180 9568
rect 34333 9571 34391 9577
rect 30699 9537 30711 9540
rect 30653 9531 30711 9537
rect 34333 9537 34345 9571
rect 34379 9537 34391 9571
rect 34333 9531 34391 9537
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 30340 9472 31754 9500
rect 30340 9460 30346 9472
rect 31726 9432 31754 9472
rect 32766 9460 32772 9512
rect 32824 9460 32830 9512
rect 32858 9460 32864 9512
rect 32916 9460 32922 9512
rect 32950 9460 32956 9512
rect 33008 9500 33014 9512
rect 34348 9500 34376 9531
rect 34514 9528 34520 9580
rect 34572 9528 34578 9580
rect 37829 9571 37887 9577
rect 37829 9537 37841 9571
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 34698 9500 34704 9512
rect 33008 9472 34704 9500
rect 33008 9460 33014 9472
rect 34698 9460 34704 9472
rect 34756 9460 34762 9512
rect 37844 9432 37872 9531
rect 31726 9404 37872 9432
rect 30558 9364 30564 9376
rect 29472 9336 30564 9364
rect 30558 9324 30564 9336
rect 30616 9324 30622 9376
rect 31202 9324 31208 9376
rect 31260 9364 31266 9376
rect 32309 9367 32367 9373
rect 32309 9364 32321 9367
rect 31260 9336 32321 9364
rect 31260 9324 31266 9336
rect 32309 9333 32321 9336
rect 32355 9333 32367 9367
rect 32309 9327 32367 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 16206 9160 16212 9172
rect 10836 9132 16212 9160
rect 10836 9120 10842 9132
rect 16206 9120 16212 9132
rect 16264 9160 16270 9172
rect 17770 9160 17776 9172
rect 16264 9132 17776 9160
rect 16264 9120 16270 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19392 9132 20944 9160
rect 19392 9120 19398 9132
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 17586 9092 17592 9104
rect 15712 9064 17592 9092
rect 15712 9052 15718 9064
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 20806 9052 20812 9104
rect 20864 9052 20870 9104
rect 20916 9092 20944 9132
rect 25314 9120 25320 9172
rect 25372 9120 25378 9172
rect 30009 9163 30067 9169
rect 30009 9129 30021 9163
rect 30055 9160 30067 9163
rect 30650 9160 30656 9172
rect 30055 9132 30656 9160
rect 30055 9129 30067 9132
rect 30009 9123 30067 9129
rect 30650 9120 30656 9132
rect 30708 9160 30714 9172
rect 32858 9160 32864 9172
rect 30708 9132 32864 9160
rect 30708 9120 30714 9132
rect 32858 9120 32864 9132
rect 32916 9120 32922 9172
rect 36262 9120 36268 9172
rect 36320 9120 36326 9172
rect 30558 9092 30564 9104
rect 20916 9064 30564 9092
rect 30558 9052 30564 9064
rect 30616 9052 30622 9104
rect 32030 9052 32036 9104
rect 32088 9092 32094 9104
rect 32309 9095 32367 9101
rect 32309 9092 32321 9095
rect 32088 9064 32321 9092
rect 32088 9052 32094 9064
rect 32309 9061 32321 9064
rect 32355 9061 32367 9095
rect 32309 9055 32367 9061
rect 35618 9052 35624 9104
rect 35676 9052 35682 9104
rect 36280 9092 36308 9120
rect 36280 9064 36768 9092
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 17034 9024 17040 9036
rect 16439 8996 17040 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 17034 8984 17040 8996
rect 17092 8984 17098 9036
rect 14550 8916 14556 8968
rect 14608 8916 14614 8968
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 14792 8928 15393 8956
rect 14792 8916 14798 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 16482 8956 16488 8968
rect 15795 8928 16488 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 14366 8848 14372 8900
rect 14424 8848 14430 8900
rect 15580 8888 15608 8919
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 17604 8965 17632 9052
rect 19981 9027 20039 9033
rect 18892 8996 19840 9024
rect 18892 8965 18920 8996
rect 19812 8968 19840 8996
rect 19981 8993 19993 9027
rect 20027 9024 20039 9027
rect 20070 9024 20076 9036
rect 20027 8996 20076 9024
rect 20027 8993 20039 8996
rect 19981 8987 20039 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 21082 8984 21088 9036
rect 21140 9024 21146 9036
rect 21177 9027 21235 9033
rect 21177 9024 21189 9027
rect 21140 8996 21189 9024
rect 21140 8984 21146 8996
rect 21177 8993 21189 8996
rect 21223 8993 21235 9027
rect 21177 8987 21235 8993
rect 21361 9027 21419 9033
rect 21361 8993 21373 9027
rect 21407 9024 21419 9027
rect 22002 9024 22008 9036
rect 21407 8996 22008 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 27246 8984 27252 9036
rect 27304 8984 27310 9036
rect 28092 8996 30604 9024
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 16022 8888 16028 8900
rect 15580 8860 16028 8888
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 16577 8891 16635 8897
rect 16577 8857 16589 8891
rect 16623 8888 16635 8891
rect 17497 8891 17555 8897
rect 17497 8888 17509 8891
rect 16623 8860 17509 8888
rect 16623 8857 16635 8860
rect 16577 8851 16635 8857
rect 17497 8857 17509 8860
rect 17543 8857 17555 8891
rect 17497 8851 17555 8857
rect 18325 8891 18383 8897
rect 18325 8857 18337 8891
rect 18371 8888 18383 8891
rect 18414 8888 18420 8900
rect 18371 8860 18420 8888
rect 18371 8857 18383 8860
rect 18325 8851 18383 8857
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 18708 8888 18736 8919
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19208 8928 19441 8956
rect 19208 8916 19214 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19794 8916 19800 8968
rect 19852 8916 19858 8968
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 24946 8916 24952 8968
rect 25004 8916 25010 8968
rect 25130 8916 25136 8968
rect 25188 8916 25194 8968
rect 26694 8916 26700 8968
rect 26752 8956 26758 8968
rect 28092 8965 28120 8996
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 26752 8928 28089 8956
rect 26752 8916 26758 8928
rect 28077 8925 28089 8928
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 30190 8916 30196 8968
rect 30248 8916 30254 8968
rect 30466 8916 30472 8968
rect 30524 8916 30530 8968
rect 30576 8956 30604 8996
rect 33042 8984 33048 9036
rect 33100 8984 33106 9036
rect 36262 8984 36268 9036
rect 36320 8984 36326 9036
rect 36740 9033 36768 9064
rect 36725 9027 36783 9033
rect 36725 8993 36737 9027
rect 36771 8993 36783 9027
rect 36725 8987 36783 8993
rect 30576 8928 30880 8956
rect 19168 8888 19196 8916
rect 18708 8860 19196 8888
rect 19521 8891 19579 8897
rect 19521 8857 19533 8891
rect 19567 8857 19579 8891
rect 19521 8851 19579 8857
rect 21269 8891 21327 8897
rect 21269 8857 21281 8891
rect 21315 8888 21327 8891
rect 22462 8888 22468 8900
rect 21315 8860 22468 8888
rect 21315 8857 21327 8860
rect 21269 8851 21327 8857
rect 16945 8823 17003 8829
rect 16945 8789 16957 8823
rect 16991 8820 17003 8823
rect 17126 8820 17132 8832
rect 16991 8792 17132 8820
rect 16991 8789 17003 8792
rect 16945 8783 17003 8789
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19536 8820 19564 8851
rect 22462 8848 22468 8860
rect 22520 8848 22526 8900
rect 24302 8848 24308 8900
rect 24360 8888 24366 8900
rect 25869 8891 25927 8897
rect 25869 8888 25881 8891
rect 24360 8860 25881 8888
rect 24360 8848 24366 8860
rect 25869 8857 25881 8860
rect 25915 8888 25927 8891
rect 26418 8888 26424 8900
rect 25915 8860 26424 8888
rect 25915 8857 25927 8860
rect 25869 8851 25927 8857
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 29362 8888 29368 8900
rect 26804 8860 29368 8888
rect 19024 8792 19564 8820
rect 19024 8780 19030 8792
rect 25406 8780 25412 8832
rect 25464 8820 25470 8832
rect 26804 8820 26832 8860
rect 29362 8848 29368 8860
rect 29420 8888 29426 8900
rect 30285 8891 30343 8897
rect 30285 8888 30297 8891
rect 29420 8860 30297 8888
rect 29420 8848 29426 8860
rect 30285 8857 30297 8860
rect 30331 8888 30343 8891
rect 30742 8888 30748 8900
rect 30331 8860 30748 8888
rect 30331 8857 30343 8860
rect 30285 8851 30343 8857
rect 30742 8848 30748 8860
rect 30800 8848 30806 8900
rect 30852 8888 30880 8928
rect 30926 8916 30932 8968
rect 30984 8916 30990 8968
rect 33778 8956 33784 8968
rect 31036 8928 33784 8956
rect 31036 8888 31064 8928
rect 33778 8916 33784 8928
rect 33836 8956 33842 8968
rect 33873 8959 33931 8965
rect 33873 8956 33885 8959
rect 33836 8928 33885 8956
rect 33836 8916 33842 8928
rect 33873 8925 33885 8928
rect 33919 8925 33931 8959
rect 33873 8919 33931 8925
rect 35526 8916 35532 8968
rect 35584 8916 35590 8968
rect 36354 8916 36360 8968
rect 36412 8916 36418 8968
rect 37001 8959 37059 8965
rect 37001 8925 37013 8959
rect 37047 8925 37059 8959
rect 37001 8919 37059 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 31202 8897 31208 8900
rect 31196 8888 31208 8897
rect 30852 8860 31064 8888
rect 31163 8860 31208 8888
rect 31196 8851 31208 8860
rect 31202 8848 31208 8851
rect 31260 8848 31266 8900
rect 37016 8888 37044 8919
rect 37734 8888 37740 8900
rect 37016 8860 37740 8888
rect 37734 8848 37740 8860
rect 37792 8848 37798 8900
rect 25464 8792 26832 8820
rect 25464 8780 25470 8792
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 28810 8820 28816 8832
rect 26936 8792 28816 8820
rect 26936 8780 26942 8792
rect 28810 8780 28816 8792
rect 28868 8780 28874 8832
rect 30760 8820 30788 8848
rect 32950 8820 32956 8832
rect 30760 8792 32956 8820
rect 32950 8780 32956 8792
rect 33008 8780 33014 8832
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 37844 8820 37872 8919
rect 38102 8848 38108 8900
rect 38160 8848 38166 8900
rect 34848 8792 37872 8820
rect 34848 8780 34854 8792
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11296 8588 12081 8616
rect 11296 8576 11302 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 20898 8616 20904 8628
rect 14700 8588 20904 8616
rect 14700 8576 14706 8588
rect 12621 8551 12679 8557
rect 12621 8517 12633 8551
rect 12667 8548 12679 8551
rect 13078 8548 13084 8560
rect 12667 8520 13084 8548
rect 12667 8517 12679 8520
rect 12621 8511 12679 8517
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 19812 8557 19840 8588
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 25188 8588 25697 8616
rect 25188 8576 25194 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 27525 8619 27583 8625
rect 27525 8616 27537 8619
rect 27488 8588 27537 8616
rect 27488 8576 27494 8588
rect 27525 8585 27537 8588
rect 27571 8585 27583 8619
rect 27525 8579 27583 8585
rect 27893 8619 27951 8625
rect 27893 8585 27905 8619
rect 27939 8616 27951 8619
rect 28534 8616 28540 8628
rect 27939 8588 28540 8616
rect 27939 8585 27951 8588
rect 27893 8579 27951 8585
rect 28534 8576 28540 8588
rect 28592 8576 28598 8628
rect 29822 8576 29828 8628
rect 29880 8616 29886 8628
rect 34790 8616 34796 8628
rect 29880 8588 34796 8616
rect 29880 8576 29886 8588
rect 34790 8576 34796 8588
rect 34848 8576 34854 8628
rect 36262 8576 36268 8628
rect 36320 8616 36326 8628
rect 36357 8619 36415 8625
rect 36357 8616 36369 8619
rect 36320 8588 36369 8616
rect 36320 8576 36326 8588
rect 36357 8585 36369 8588
rect 36403 8585 36415 8619
rect 36357 8579 36415 8585
rect 37734 8576 37740 8628
rect 37792 8616 37798 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 37792 8588 37841 8616
rect 37792 8576 37798 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 19797 8551 19855 8557
rect 15948 8520 17172 8548
rect 11790 8440 11796 8492
rect 11848 8440 11854 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12575 8452 12756 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 11900 8412 11928 8443
rect 12728 8412 12756 8452
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 15948 8489 15976 8520
rect 17144 8492 17172 8520
rect 19797 8517 19809 8551
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 19978 8508 19984 8560
rect 20036 8508 20042 8560
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 20625 8551 20683 8557
rect 20625 8548 20637 8551
rect 20128 8520 20637 8548
rect 20128 8508 20134 8520
rect 20625 8517 20637 8520
rect 20671 8517 20683 8551
rect 20625 8511 20683 8517
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 30190 8548 30196 8560
rect 23440 8520 30196 8548
rect 23440 8508 23446 8520
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 16224 8412 16252 8443
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16356 8452 16865 8480
rect 16356 8440 16362 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18414 8480 18420 8492
rect 18371 8452 18420 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 24572 8483 24630 8489
rect 24572 8449 24584 8483
rect 24618 8480 24630 8483
rect 24854 8480 24860 8492
rect 24618 8452 24860 8480
rect 24618 8449 24630 8452
rect 24572 8443 24630 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 25038 8440 25044 8492
rect 25096 8480 25102 8492
rect 25096 8452 26234 8480
rect 25096 8440 25102 8452
rect 16960 8412 16988 8440
rect 11900 8384 12572 8412
rect 12728 8384 13768 8412
rect 16224 8384 16988 8412
rect 12544 8353 12572 8384
rect 13740 8356 13768 8384
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18288 8384 18521 8412
rect 18288 8372 18294 8384
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8412 19671 8415
rect 21266 8412 21272 8424
rect 19659 8384 21272 8412
rect 19659 8381 19671 8384
rect 19613 8375 19671 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 24302 8412 24308 8424
rect 22112 8384 24308 8412
rect 12529 8347 12587 8353
rect 12529 8313 12541 8347
rect 12575 8313 12587 8347
rect 12529 8307 12587 8313
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 13780 8316 14013 8344
rect 13780 8304 13786 8316
rect 14001 8313 14013 8316
rect 14047 8313 14059 8347
rect 14001 8307 14059 8313
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 16540 8316 17325 8344
rect 16540 8304 16546 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 20441 8347 20499 8353
rect 20441 8313 20453 8347
rect 20487 8344 20499 8347
rect 20714 8344 20720 8356
rect 20487 8316 20720 8344
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 15712 8248 15761 8276
rect 15712 8236 15718 8248
rect 15749 8245 15761 8248
rect 15795 8245 15807 8279
rect 15749 8239 15807 8245
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 22112 8276 22140 8384
rect 24302 8372 24308 8384
rect 24360 8372 24366 8424
rect 26206 8412 26234 8452
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 29196 8489 29224 8520
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 31294 8508 31300 8560
rect 31352 8508 31358 8560
rect 33778 8508 33784 8560
rect 33836 8508 33842 8560
rect 36814 8548 36820 8560
rect 34992 8520 36820 8548
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 27672 8452 27997 8480
rect 27672 8440 27678 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 29181 8483 29239 8489
rect 29181 8449 29193 8483
rect 29227 8449 29239 8483
rect 29181 8443 29239 8449
rect 29273 8483 29331 8489
rect 29273 8449 29285 8483
rect 29319 8480 29331 8483
rect 29362 8480 29368 8492
rect 29319 8452 29368 8480
rect 29319 8449 29331 8452
rect 29273 8443 29331 8449
rect 29362 8440 29368 8452
rect 29420 8440 29426 8492
rect 30466 8440 30472 8492
rect 30524 8440 30530 8492
rect 30742 8440 30748 8492
rect 30800 8440 30806 8492
rect 32950 8440 32956 8492
rect 33008 8480 33014 8492
rect 34992 8489 35020 8520
rect 36814 8508 36820 8520
rect 36872 8508 36878 8560
rect 35250 8489 35256 8492
rect 33045 8483 33103 8489
rect 33045 8480 33057 8483
rect 33008 8452 33057 8480
rect 33008 8440 33014 8452
rect 33045 8449 33057 8452
rect 33091 8480 33103 8483
rect 34977 8483 35035 8489
rect 34977 8480 34989 8483
rect 33091 8452 34989 8480
rect 33091 8449 33103 8452
rect 33045 8443 33103 8449
rect 34977 8449 34989 8452
rect 35023 8449 35035 8483
rect 34977 8443 35035 8449
rect 35244 8443 35256 8489
rect 35250 8440 35256 8443
rect 35308 8440 35314 8492
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 26206 8384 28089 8412
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 28258 8372 28264 8424
rect 28316 8412 28322 8424
rect 30484 8412 30512 8440
rect 34238 8412 34244 8424
rect 28316 8384 34244 8412
rect 28316 8372 28322 8384
rect 34238 8372 34244 8384
rect 34296 8372 34302 8424
rect 35986 8372 35992 8424
rect 36044 8412 36050 8424
rect 37921 8415 37979 8421
rect 37921 8412 37933 8415
rect 36044 8384 37933 8412
rect 36044 8372 36050 8384
rect 37921 8381 37933 8384
rect 37967 8381 37979 8415
rect 37921 8375 37979 8381
rect 38010 8372 38016 8424
rect 38068 8372 38074 8424
rect 29454 8304 29460 8356
rect 29512 8344 29518 8356
rect 32122 8344 32128 8356
rect 29512 8316 32128 8344
rect 29512 8304 29518 8316
rect 32122 8304 32128 8316
rect 32180 8304 32186 8356
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 37461 8347 37519 8353
rect 37461 8344 37473 8347
rect 37240 8316 37473 8344
rect 37240 8304 37246 8316
rect 37461 8313 37473 8316
rect 37507 8313 37519 8347
rect 37461 8307 37519 8313
rect 21600 8248 22140 8276
rect 21600 8236 21606 8248
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 28997 8279 29055 8285
rect 28997 8276 29009 8279
rect 27856 8248 29009 8276
rect 27856 8236 27862 8248
rect 28997 8245 29009 8248
rect 29043 8276 29055 8279
rect 33042 8276 33048 8288
rect 29043 8248 33048 8276
rect 29043 8245 29055 8248
rect 28997 8239 29055 8245
rect 33042 8236 33048 8248
rect 33100 8236 33106 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 15528 8044 15577 8072
rect 15528 8032 15534 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 16080 8044 16221 8072
rect 16080 8032 16086 8044
rect 16209 8041 16221 8044
rect 16255 8041 16267 8075
rect 16209 8035 16267 8041
rect 16546 8044 22508 8072
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 14148 7976 14473 8004
rect 14148 7964 14154 7976
rect 14461 7973 14473 7976
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 11054 7936 11060 7948
rect 10643 7908 11060 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7936 12311 7939
rect 16546 7936 16574 8044
rect 22480 8004 22508 8044
rect 22922 8032 22928 8084
rect 22980 8032 22986 8084
rect 24854 8032 24860 8084
rect 24912 8032 24918 8084
rect 28629 8075 28687 8081
rect 28629 8041 28641 8075
rect 28675 8072 28687 8075
rect 28994 8072 29000 8084
rect 28675 8044 29000 8072
rect 28675 8041 28687 8044
rect 28629 8035 28687 8041
rect 28994 8032 29000 8044
rect 29052 8032 29058 8084
rect 31202 8072 31208 8084
rect 30300 8044 31208 8072
rect 23198 8004 23204 8016
rect 22480 7976 23204 8004
rect 23198 7964 23204 7976
rect 23256 7964 23262 8016
rect 25222 7964 25228 8016
rect 25280 7964 25286 8016
rect 20990 7936 20996 7948
rect 12299 7908 16574 7936
rect 20548 7908 20996 7936
rect 12299 7905 12311 7908
rect 12253 7899 12311 7905
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 11146 7868 11152 7880
rect 10919 7840 11152 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11146 7828 11152 7840
rect 11204 7868 11210 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 11204 7840 12725 7868
rect 11204 7828 11210 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 14240 7840 14289 7868
rect 14240 7828 14246 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14424 7840 14933 7868
rect 14424 7828 14430 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 15528 7840 16313 7868
rect 15528 7828 15534 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18506 7868 18512 7880
rect 18279 7840 18512 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18064 7800 18092 7831
rect 18506 7828 18512 7840
rect 18564 7868 18570 7880
rect 20548 7877 20576 7908
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 25240 7936 25268 7964
rect 25317 7939 25375 7945
rect 25317 7936 25329 7939
rect 25240 7908 25329 7936
rect 25317 7905 25329 7908
rect 25363 7905 25375 7939
rect 25317 7899 25375 7905
rect 25498 7896 25504 7948
rect 25556 7896 25562 7948
rect 29086 7896 29092 7948
rect 29144 7936 29150 7948
rect 30300 7945 30328 8044
rect 31202 8032 31208 8044
rect 31260 8032 31266 8084
rect 32398 8032 32404 8084
rect 32456 8072 32462 8084
rect 32456 8044 33824 8072
rect 32456 8032 32462 8044
rect 32217 8007 32275 8013
rect 32217 7973 32229 8007
rect 32263 7973 32275 8007
rect 32217 7967 32275 7973
rect 29733 7939 29791 7945
rect 29733 7936 29745 7939
rect 29144 7908 29745 7936
rect 29144 7896 29150 7908
rect 29733 7905 29745 7908
rect 29779 7905 29791 7939
rect 29733 7899 29791 7905
rect 30285 7939 30343 7945
rect 30285 7905 30297 7939
rect 30331 7905 30343 7939
rect 32232 7936 32260 7967
rect 33042 7964 33048 8016
rect 33100 8004 33106 8016
rect 33100 7976 33272 8004
rect 33100 7964 33106 7976
rect 33244 7945 33272 7976
rect 33229 7939 33287 7945
rect 32232 7908 33088 7936
rect 30285 7899 30343 7905
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 18564 7840 20085 7868
rect 18564 7828 18570 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20714 7828 20720 7880
rect 20772 7828 20778 7880
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 21082 7868 21088 7880
rect 20855 7840 21088 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21082 7828 21088 7840
rect 21140 7828 21146 7880
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25225 7871 25283 7877
rect 25225 7868 25237 7871
rect 25188 7840 25237 7868
rect 25188 7828 25194 7840
rect 25225 7837 25237 7840
rect 25271 7837 25283 7871
rect 25225 7831 25283 7837
rect 26418 7828 26424 7880
rect 26476 7828 26482 7880
rect 28258 7828 28264 7880
rect 28316 7828 28322 7880
rect 30190 7828 30196 7880
rect 30248 7828 30254 7880
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7868 30895 7871
rect 30926 7868 30932 7880
rect 30883 7840 30932 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 30926 7828 30932 7840
rect 30984 7868 30990 7880
rect 32950 7868 32956 7880
rect 30984 7840 32956 7868
rect 30984 7828 30990 7840
rect 32950 7828 32956 7840
rect 33008 7828 33014 7880
rect 33060 7877 33088 7908
rect 33229 7905 33241 7939
rect 33275 7905 33287 7939
rect 33796 7936 33824 8044
rect 33870 8032 33876 8084
rect 33928 8032 33934 8084
rect 35253 8075 35311 8081
rect 35253 8041 35265 8075
rect 35299 8072 35311 8075
rect 35342 8072 35348 8084
rect 35299 8044 35348 8072
rect 35299 8041 35311 8044
rect 35253 8035 35311 8041
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 37826 8032 37832 8084
rect 37884 8072 37890 8084
rect 38289 8075 38347 8081
rect 38289 8072 38301 8075
rect 37884 8044 38301 8072
rect 37884 8032 37890 8044
rect 38289 8041 38301 8044
rect 38335 8041 38347 8075
rect 38289 8035 38347 8041
rect 35986 8004 35992 8016
rect 35728 7976 35992 8004
rect 35728 7945 35756 7976
rect 35986 7964 35992 7976
rect 36044 7964 36050 8016
rect 35713 7939 35771 7945
rect 35713 7936 35725 7939
rect 33796 7908 35725 7936
rect 33229 7899 33287 7905
rect 35713 7905 35725 7908
rect 35759 7905 35771 7939
rect 35713 7899 35771 7905
rect 35802 7896 35808 7948
rect 35860 7896 35866 7948
rect 33045 7871 33103 7877
rect 33045 7837 33057 7871
rect 33091 7868 33103 7871
rect 34057 7871 34115 7877
rect 34057 7868 34069 7871
rect 33091 7840 34069 7868
rect 33091 7837 33103 7840
rect 33045 7831 33103 7837
rect 34057 7837 34069 7840
rect 34103 7837 34115 7871
rect 34057 7831 34115 7837
rect 34238 7828 34244 7880
rect 34296 7828 34302 7880
rect 35621 7871 35679 7877
rect 35621 7837 35633 7871
rect 35667 7868 35679 7871
rect 36262 7868 36268 7880
rect 35667 7840 36268 7868
rect 35667 7837 35679 7840
rect 35621 7831 35679 7837
rect 36262 7828 36268 7840
rect 36320 7828 36326 7880
rect 36814 7828 36820 7880
rect 36872 7868 36878 7880
rect 37182 7877 37188 7880
rect 36909 7871 36967 7877
rect 36909 7868 36921 7871
rect 36872 7840 36921 7868
rect 36872 7828 36878 7840
rect 36909 7837 36921 7840
rect 36955 7837 36967 7871
rect 37176 7868 37188 7877
rect 37143 7840 37188 7868
rect 36909 7831 36967 7837
rect 37176 7831 37188 7840
rect 37182 7828 37188 7831
rect 37240 7828 37246 7880
rect 18966 7800 18972 7812
rect 18012 7772 18972 7800
rect 18012 7760 18018 7772
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 21812 7803 21870 7809
rect 21812 7769 21824 7803
rect 21858 7800 21870 7803
rect 22002 7800 22008 7812
rect 21858 7772 22008 7800
rect 21858 7769 21870 7772
rect 21812 7763 21870 7769
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 26688 7803 26746 7809
rect 26688 7769 26700 7803
rect 26734 7800 26746 7803
rect 27154 7800 27160 7812
rect 26734 7772 27160 7800
rect 26734 7769 26746 7772
rect 26688 7763 26746 7769
rect 27154 7760 27160 7772
rect 27212 7760 27218 7812
rect 28445 7803 28503 7809
rect 28445 7769 28457 7803
rect 28491 7769 28503 7803
rect 28445 7763 28503 7769
rect 31104 7803 31162 7809
rect 31104 7769 31116 7803
rect 31150 7800 31162 7803
rect 31150 7772 32720 7800
rect 31150 7769 31162 7772
rect 31104 7763 31162 7769
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 19426 7732 19432 7744
rect 18187 7704 19432 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 27522 7692 27528 7744
rect 27580 7732 27586 7744
rect 27801 7735 27859 7741
rect 27801 7732 27813 7735
rect 27580 7704 27813 7732
rect 27580 7692 27586 7704
rect 27801 7701 27813 7704
rect 27847 7732 27859 7735
rect 28460 7732 28488 7763
rect 32692 7741 32720 7772
rect 32766 7760 32772 7812
rect 32824 7800 32830 7812
rect 33137 7803 33195 7809
rect 33137 7800 33149 7803
rect 32824 7772 33149 7800
rect 32824 7760 32830 7772
rect 33137 7769 33149 7772
rect 33183 7769 33195 7803
rect 33137 7763 33195 7769
rect 27847 7704 28488 7732
rect 32677 7735 32735 7741
rect 27847 7701 27859 7704
rect 27801 7695 27859 7701
rect 32677 7701 32689 7735
rect 32723 7701 32735 7735
rect 32677 7695 32735 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 11790 7488 11796 7540
rect 11848 7488 11854 7540
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 12207 7500 13308 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 12802 7460 12808 7472
rect 11992 7432 12808 7460
rect 11992 7401 12020 7432
rect 12802 7420 12808 7432
rect 12860 7420 12866 7472
rect 13280 7460 13308 7500
rect 21082 7488 21088 7540
rect 21140 7488 21146 7540
rect 22002 7488 22008 7540
rect 22060 7488 22066 7540
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 24147 7531 24205 7537
rect 24147 7528 24159 7531
rect 23808 7500 24159 7528
rect 23808 7488 23814 7500
rect 24147 7497 24159 7500
rect 24193 7528 24205 7531
rect 24762 7528 24768 7540
rect 24193 7500 24768 7528
rect 24193 7497 24205 7500
rect 24147 7491 24205 7497
rect 24762 7488 24768 7500
rect 24820 7528 24826 7540
rect 26234 7528 26240 7540
rect 24820 7500 26240 7528
rect 24820 7488 24826 7500
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 27154 7488 27160 7540
rect 27212 7488 27218 7540
rect 27522 7488 27528 7540
rect 27580 7488 27586 7540
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 28960 7500 37872 7528
rect 28960 7488 28966 7500
rect 13280 7432 13768 7460
rect 13740 7404 13768 7432
rect 18414 7420 18420 7472
rect 18472 7460 18478 7472
rect 18472 7432 18920 7460
rect 18472 7420 18478 7432
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12299 7364 13124 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 13096 7336 13124 7364
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 14090 7352 14096 7404
rect 14148 7352 14154 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14734 7392 14740 7404
rect 14507 7364 14740 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15654 7392 15660 7404
rect 15615 7364 15660 7392
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16482 7392 16488 7404
rect 15795 7364 16488 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 18892 7401 18920 7432
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19024 7432 20300 7460
rect 19024 7420 19030 7432
rect 20272 7401 20300 7432
rect 23934 7420 23940 7472
rect 23992 7420 23998 7472
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 27617 7463 27675 7469
rect 27617 7460 27629 7463
rect 27488 7432 27629 7460
rect 27488 7420 27494 7432
rect 27617 7429 27629 7432
rect 27663 7429 27675 7463
rect 27617 7423 27675 7429
rect 32944 7463 33002 7469
rect 32944 7429 32956 7463
rect 32990 7460 33002 7463
rect 33134 7460 33140 7472
rect 32990 7432 33140 7460
rect 32990 7429 33002 7432
rect 32944 7423 33002 7429
rect 33134 7420 33140 7432
rect 33192 7420 33198 7472
rect 35345 7463 35403 7469
rect 35345 7429 35357 7463
rect 35391 7460 35403 7463
rect 35710 7460 35716 7472
rect 35391 7432 35716 7460
rect 35391 7429 35403 7432
rect 35345 7423 35403 7429
rect 35710 7420 35716 7432
rect 35768 7420 35774 7472
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7361 20315 7395
rect 20806 7392 20812 7404
rect 20257 7355 20315 7361
rect 20456 7364 20812 7392
rect 13078 7284 13084 7336
rect 13136 7324 13142 7336
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 13136 7296 13369 7324
rect 13136 7284 13142 7296
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 14642 7284 14648 7336
rect 14700 7284 14706 7336
rect 18322 7284 18328 7336
rect 18380 7324 18386 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18380 7296 18429 7324
rect 18380 7284 18386 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18524 7324 18552 7352
rect 20180 7324 20208 7355
rect 20456 7333 20484 7364
rect 20806 7352 20812 7364
rect 20864 7392 20870 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20864 7364 21005 7392
rect 20864 7352 20870 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 20993 7355 21051 7361
rect 21100 7364 22017 7392
rect 18524 7296 20208 7324
rect 20441 7327 20499 7333
rect 18417 7287 18475 7293
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20898 7324 20904 7336
rect 20579 7296 20904 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 19242 7216 19248 7268
rect 19300 7216 19306 7268
rect 21100 7256 21128 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 22152 7364 22201 7392
rect 22152 7352 22158 7364
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 32677 7395 32735 7401
rect 32677 7361 32689 7395
rect 32723 7392 32735 7395
rect 32766 7392 32772 7404
rect 32723 7364 32772 7392
rect 32723 7361 32735 7364
rect 32677 7355 32735 7361
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 34698 7352 34704 7404
rect 34756 7352 34762 7404
rect 34790 7352 34796 7404
rect 34848 7392 34854 7404
rect 34885 7395 34943 7401
rect 34885 7392 34897 7395
rect 34848 7364 34897 7392
rect 34848 7352 34854 7364
rect 34885 7361 34897 7364
rect 34931 7361 34943 7395
rect 34885 7355 34943 7361
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7361 35035 7395
rect 34977 7355 35035 7361
rect 35069 7395 35127 7401
rect 35069 7361 35081 7395
rect 35115 7392 35127 7395
rect 37734 7392 37740 7404
rect 35115 7364 37740 7392
rect 35115 7361 35127 7364
rect 35069 7355 35127 7361
rect 25498 7284 25504 7336
rect 25556 7324 25562 7336
rect 25866 7324 25872 7336
rect 25556 7296 25872 7324
rect 25556 7284 25562 7296
rect 25866 7284 25872 7296
rect 25924 7324 25930 7336
rect 27798 7324 27804 7336
rect 25924 7296 27804 7324
rect 25924 7284 25930 7296
rect 27798 7284 27804 7296
rect 27856 7284 27862 7336
rect 34606 7284 34612 7336
rect 34664 7324 34670 7336
rect 34992 7324 35020 7355
rect 37734 7352 37740 7364
rect 37792 7352 37798 7404
rect 37844 7401 37872 7500
rect 37829 7395 37887 7401
rect 37829 7361 37841 7395
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 34664 7296 35020 7324
rect 34664 7284 34670 7296
rect 38102 7284 38108 7336
rect 38160 7284 38166 7336
rect 20364 7228 21128 7256
rect 20364 7200 20392 7228
rect 15562 7148 15568 7200
rect 15620 7148 15626 7200
rect 19981 7191 20039 7197
rect 19981 7157 19993 7191
rect 20027 7188 20039 7191
rect 20346 7188 20352 7200
rect 20027 7160 20352 7188
rect 20027 7157 20039 7160
rect 19981 7151 20039 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 24118 7148 24124 7200
rect 24176 7148 24182 7200
rect 24302 7148 24308 7200
rect 24360 7148 24366 7200
rect 34054 7148 34060 7200
rect 34112 7148 34118 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 14277 6987 14335 6993
rect 14277 6984 14289 6987
rect 12952 6956 14289 6984
rect 12952 6944 12958 6956
rect 14277 6953 14289 6956
rect 14323 6953 14335 6987
rect 14277 6947 14335 6953
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18506 6984 18512 6996
rect 18288 6956 18512 6984
rect 18288 6944 18294 6956
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 20346 6944 20352 6996
rect 20404 6984 20410 6996
rect 21453 6987 21511 6993
rect 21453 6984 21465 6987
rect 20404 6956 21465 6984
rect 20404 6944 20410 6956
rect 21453 6953 21465 6956
rect 21499 6953 21511 6987
rect 21453 6947 21511 6953
rect 23661 6987 23719 6993
rect 23661 6953 23673 6987
rect 23707 6984 23719 6987
rect 23934 6984 23940 6996
rect 23707 6956 23940 6984
rect 23707 6953 23719 6956
rect 23661 6947 23719 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 26326 6944 26332 6996
rect 26384 6984 26390 6996
rect 26421 6987 26479 6993
rect 26421 6984 26433 6987
rect 26384 6956 26433 6984
rect 26384 6944 26390 6956
rect 26421 6953 26433 6956
rect 26467 6953 26479 6987
rect 26421 6947 26479 6953
rect 33134 6944 33140 6996
rect 33192 6944 33198 6996
rect 37734 6944 37740 6996
rect 37792 6984 37798 6996
rect 38105 6987 38163 6993
rect 38105 6984 38117 6987
rect 37792 6956 38117 6984
rect 37792 6944 37798 6956
rect 38105 6953 38117 6956
rect 38151 6953 38163 6987
rect 38105 6947 38163 6953
rect 13722 6876 13728 6928
rect 13780 6916 13786 6928
rect 13780 6888 13860 6916
rect 13780 6876 13786 6888
rect 13832 6848 13860 6888
rect 13832 6820 14596 6848
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14568 6789 14596 6820
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14700 6820 14872 6848
rect 14700 6808 14706 6820
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14056 6752 14473 6780
rect 14056 6740 14062 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14734 6740 14740 6792
rect 14792 6740 14798 6792
rect 14844 6789 14872 6820
rect 15654 6808 15660 6860
rect 15712 6808 15718 6860
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6848 17923 6851
rect 17954 6848 17960 6860
rect 17911 6820 17960 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18414 6848 18420 6860
rect 18064 6820 18420 6848
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15528 6752 15853 6780
rect 15528 6740 15534 6752
rect 15841 6749 15853 6752
rect 15887 6780 15899 6783
rect 15930 6780 15936 6792
rect 15887 6752 15936 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16482 6740 16488 6792
rect 16540 6740 16546 6792
rect 18064 6789 18092 6820
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 20732 6820 22416 6848
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 20027 6752 20300 6780
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 18340 6712 18368 6740
rect 16500 6684 18368 6712
rect 16500 6653 16528 6684
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6613 16543 6647
rect 20272 6644 20300 6752
rect 20622 6740 20628 6792
rect 20680 6740 20686 6792
rect 20732 6789 20760 6820
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 22186 6780 22192 6792
rect 21600 6752 22192 6780
rect 21600 6740 21606 6752
rect 22186 6740 22192 6752
rect 22244 6780 22250 6792
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 22244 6752 22293 6780
rect 22244 6740 22250 6752
rect 22281 6749 22293 6752
rect 22327 6749 22339 6783
rect 22388 6780 22416 6820
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 24946 6848 24952 6860
rect 24176 6820 24952 6848
rect 24176 6808 24182 6820
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 25406 6808 25412 6860
rect 25464 6848 25470 6860
rect 25869 6851 25927 6857
rect 25869 6848 25881 6851
rect 25464 6820 25881 6848
rect 25464 6808 25470 6820
rect 25869 6817 25881 6820
rect 25915 6817 25927 6851
rect 27525 6851 27583 6857
rect 25869 6811 25927 6817
rect 25976 6820 27476 6848
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 22388 6752 24685 6780
rect 22281 6743 22339 6749
rect 24673 6749 24685 6752
rect 24719 6780 24731 6783
rect 25976 6780 26004 6820
rect 24719 6752 26004 6780
rect 24719 6749 24731 6752
rect 24673 6743 24731 6749
rect 26050 6740 26056 6792
rect 26108 6780 26114 6792
rect 26973 6783 27031 6789
rect 26973 6780 26985 6783
rect 26108 6752 26985 6780
rect 26108 6740 26114 6752
rect 26973 6749 26985 6752
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6749 27123 6783
rect 27448 6780 27476 6820
rect 27525 6817 27537 6851
rect 27571 6848 27583 6851
rect 28258 6848 28264 6860
rect 27571 6820 28264 6848
rect 27571 6817 27583 6820
rect 27525 6811 27583 6817
rect 28258 6808 28264 6820
rect 28316 6808 28322 6860
rect 28810 6808 28816 6860
rect 28868 6848 28874 6860
rect 29454 6848 29460 6860
rect 28868 6820 29460 6848
rect 28868 6808 28874 6820
rect 29454 6808 29460 6820
rect 29512 6808 29518 6860
rect 29546 6808 29552 6860
rect 29604 6848 29610 6860
rect 29733 6851 29791 6857
rect 29733 6848 29745 6851
rect 29604 6820 29745 6848
rect 29604 6808 29610 6820
rect 29733 6817 29745 6820
rect 29779 6817 29791 6851
rect 30558 6848 30564 6860
rect 29733 6811 29791 6817
rect 30208 6820 30564 6848
rect 29270 6780 29276 6792
rect 27448 6752 29276 6780
rect 27065 6743 27123 6749
rect 21082 6672 21088 6724
rect 21140 6712 21146 6724
rect 21266 6712 21272 6724
rect 21140 6684 21272 6712
rect 21140 6672 21146 6684
rect 21266 6672 21272 6684
rect 21324 6672 21330 6724
rect 22548 6715 22606 6721
rect 21376 6684 21772 6712
rect 21376 6644 21404 6684
rect 20272 6616 21404 6644
rect 16485 6607 16543 6613
rect 21450 6604 21456 6656
rect 21508 6653 21514 6656
rect 21508 6647 21527 6653
rect 21515 6613 21527 6647
rect 21508 6607 21527 6613
rect 21508 6604 21514 6607
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 21744 6644 21772 6684
rect 22548 6681 22560 6715
rect 22594 6712 22606 6715
rect 23198 6712 23204 6724
rect 22594 6684 23204 6712
rect 22594 6681 22606 6684
rect 22548 6675 22606 6681
rect 23198 6672 23204 6684
rect 23256 6672 23262 6724
rect 25225 6715 25283 6721
rect 25225 6681 25237 6715
rect 25271 6712 25283 6715
rect 25314 6712 25320 6724
rect 25271 6684 25320 6712
rect 25271 6681 25283 6684
rect 25225 6675 25283 6681
rect 25314 6672 25320 6684
rect 25372 6712 25378 6724
rect 25372 6684 26096 6712
rect 25372 6672 25378 6684
rect 23750 6644 23756 6656
rect 21744 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 25406 6604 25412 6656
rect 25464 6644 25470 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25464 6616 25973 6644
rect 25464 6604 25470 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 26068 6644 26096 6684
rect 26142 6672 26148 6724
rect 26200 6672 26206 6724
rect 26234 6672 26240 6724
rect 26292 6712 26298 6724
rect 27080 6712 27108 6743
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 30208 6789 30236 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 33689 6851 33747 6857
rect 33689 6848 33701 6851
rect 33192 6820 33701 6848
rect 33192 6808 33198 6820
rect 33689 6817 33701 6820
rect 33735 6817 33747 6851
rect 33689 6811 33747 6817
rect 30193 6783 30251 6789
rect 30193 6749 30205 6783
rect 30239 6749 30251 6783
rect 30193 6743 30251 6749
rect 30374 6740 30380 6792
rect 30432 6740 30438 6792
rect 30469 6783 30527 6789
rect 30469 6749 30481 6783
rect 30515 6749 30527 6783
rect 30469 6743 30527 6749
rect 36725 6783 36783 6789
rect 36725 6749 36737 6783
rect 36771 6780 36783 6783
rect 36814 6780 36820 6792
rect 36771 6752 36820 6780
rect 36771 6749 36783 6752
rect 36725 6743 36783 6749
rect 26292 6684 27108 6712
rect 26292 6672 26298 6684
rect 29914 6672 29920 6724
rect 29972 6712 29978 6724
rect 30484 6712 30512 6743
rect 36814 6740 36820 6752
rect 36872 6740 36878 6792
rect 29972 6684 30512 6712
rect 33505 6715 33563 6721
rect 29972 6672 29978 6684
rect 33505 6681 33517 6715
rect 33551 6712 33563 6715
rect 34054 6712 34060 6724
rect 33551 6684 34060 6712
rect 33551 6681 33563 6684
rect 33505 6675 33563 6681
rect 34054 6672 34060 6684
rect 34112 6672 34118 6724
rect 36992 6715 37050 6721
rect 36992 6681 37004 6715
rect 37038 6712 37050 6715
rect 37458 6712 37464 6724
rect 37038 6684 37464 6712
rect 37038 6681 37050 6684
rect 36992 6675 37050 6681
rect 37458 6672 37464 6684
rect 37516 6672 37522 6724
rect 28810 6644 28816 6656
rect 26068 6616 28816 6644
rect 25961 6607 26019 6613
rect 28810 6604 28816 6616
rect 28868 6604 28874 6656
rect 33597 6647 33655 6653
rect 33597 6613 33609 6647
rect 33643 6644 33655 6647
rect 37918 6644 37924 6656
rect 33643 6616 37924 6644
rect 33643 6613 33655 6616
rect 33597 6607 33655 6613
rect 37918 6604 37924 6616
rect 37976 6604 37982 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 20680 6412 23152 6440
rect 20680 6400 20686 6412
rect 19334 6372 19340 6384
rect 19182 6344 19340 6372
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 21450 6372 21456 6384
rect 20088 6344 21456 6372
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18322 6304 18328 6316
rect 18095 6276 18328 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 18506 6264 18512 6316
rect 18564 6264 18570 6316
rect 15562 6196 15568 6248
rect 15620 6196 15626 6248
rect 16206 6196 16212 6248
rect 16264 6196 16270 6248
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 20088 6245 20116 6344
rect 21450 6332 21456 6344
rect 21508 6372 21514 6384
rect 22094 6372 22100 6384
rect 21508 6344 22100 6372
rect 21508 6332 21514 6344
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 23124 6372 23152 6412
rect 23198 6400 23204 6452
rect 23256 6400 23262 6452
rect 23569 6443 23627 6449
rect 23569 6409 23581 6443
rect 23615 6440 23627 6443
rect 23934 6440 23940 6452
rect 23615 6412 23940 6440
rect 23615 6409 23627 6412
rect 23569 6403 23627 6409
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 24495 6443 24553 6449
rect 24495 6409 24507 6443
rect 24541 6440 24553 6443
rect 26142 6440 26148 6452
rect 24541 6412 26148 6440
rect 24541 6409 24553 6412
rect 24495 6403 24553 6409
rect 26142 6400 26148 6412
rect 26200 6400 26206 6452
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 28721 6443 28779 6449
rect 28721 6440 28733 6443
rect 28316 6412 28733 6440
rect 28316 6400 28322 6412
rect 28721 6409 28733 6412
rect 28767 6440 28779 6443
rect 29549 6443 29607 6449
rect 29549 6440 29561 6443
rect 28767 6412 29561 6440
rect 28767 6409 28779 6412
rect 28721 6403 28779 6409
rect 29549 6409 29561 6412
rect 29595 6409 29607 6443
rect 29549 6403 29607 6409
rect 29914 6400 29920 6452
rect 29972 6400 29978 6452
rect 30374 6400 30380 6452
rect 30432 6400 30438 6452
rect 34333 6443 34391 6449
rect 30668 6412 34284 6440
rect 24118 6372 24124 6384
rect 23124 6344 24124 6372
rect 24118 6332 24124 6344
rect 24176 6332 24182 6384
rect 24302 6332 24308 6384
rect 24360 6372 24366 6384
rect 24397 6375 24455 6381
rect 24397 6372 24409 6375
rect 24360 6344 24409 6372
rect 24360 6332 24366 6344
rect 24397 6341 24409 6344
rect 24443 6341 24455 6375
rect 24397 6335 24455 6341
rect 24946 6332 24952 6384
rect 25004 6372 25010 6384
rect 25004 6344 26188 6372
rect 25004 6332 25010 6344
rect 26160 6316 26188 6344
rect 20346 6264 20352 6316
rect 20404 6264 20410 6316
rect 21082 6264 21088 6316
rect 21140 6264 21146 6316
rect 21634 6264 21640 6316
rect 21692 6304 21698 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21692 6276 22017 6304
rect 21692 6264 21698 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6273 22247 6307
rect 24210 6304 24216 6316
rect 22189 6267 22247 6273
rect 23676 6276 24216 6304
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 19208 6208 20085 6236
rect 19208 6196 19214 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 22204 6236 22232 6267
rect 23676 6248 23704 6276
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 24673 6307 24731 6313
rect 24673 6273 24685 6307
rect 24719 6304 24731 6307
rect 25314 6304 25320 6316
rect 24719 6276 25320 6304
rect 24719 6273 24731 6276
rect 24673 6267 24731 6273
rect 25314 6264 25320 6276
rect 25372 6264 25378 6316
rect 25961 6307 26019 6313
rect 25961 6273 25973 6307
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 20073 6199 20131 6205
rect 20824 6208 22232 6236
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 20824 6177 20852 6208
rect 23658 6196 23664 6248
rect 23716 6196 23722 6248
rect 23845 6239 23903 6245
rect 23845 6205 23857 6239
rect 23891 6205 23903 6239
rect 25976 6236 26004 6267
rect 26142 6264 26148 6316
rect 26200 6264 26206 6316
rect 26234 6264 26240 6316
rect 26292 6264 26298 6316
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 27246 6304 27252 6316
rect 26476 6276 27252 6304
rect 26476 6264 26482 6276
rect 27246 6264 27252 6276
rect 27304 6304 27310 6316
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 27304 6276 27353 6304
rect 27304 6264 27310 6276
rect 27341 6273 27353 6276
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 27608 6307 27666 6313
rect 27608 6273 27620 6307
rect 27654 6304 27666 6307
rect 27890 6304 27896 6316
rect 27654 6276 27896 6304
rect 27654 6273 27666 6276
rect 27608 6267 27666 6273
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 28626 6264 28632 6316
rect 28684 6304 28690 6316
rect 29457 6307 29515 6313
rect 29457 6304 29469 6307
rect 28684 6276 29469 6304
rect 28684 6264 28690 6276
rect 29457 6273 29469 6276
rect 29503 6273 29515 6307
rect 29457 6267 29515 6273
rect 26050 6236 26056 6248
rect 25976 6208 26056 6236
rect 23845 6199 23903 6205
rect 20809 6171 20867 6177
rect 20809 6168 20821 6171
rect 14792 6140 20821 6168
rect 14792 6128 14798 6140
rect 20809 6137 20821 6140
rect 20855 6137 20867 6171
rect 23860 6168 23888 6199
rect 26050 6196 26056 6208
rect 26108 6196 26114 6248
rect 29270 6196 29276 6248
rect 29328 6236 29334 6248
rect 29365 6239 29423 6245
rect 29365 6236 29377 6239
rect 29328 6208 29377 6236
rect 29328 6196 29334 6208
rect 29365 6205 29377 6208
rect 29411 6236 29423 6239
rect 30668 6236 30696 6412
rect 34054 6332 34060 6384
rect 34112 6372 34118 6384
rect 34149 6375 34207 6381
rect 34149 6372 34161 6375
rect 34112 6344 34161 6372
rect 34112 6332 34118 6344
rect 34149 6341 34161 6344
rect 34195 6341 34207 6375
rect 34256 6372 34284 6412
rect 34333 6409 34345 6443
rect 34379 6440 34391 6443
rect 34698 6440 34704 6452
rect 34379 6412 34704 6440
rect 34379 6409 34391 6412
rect 34333 6403 34391 6409
rect 34698 6400 34704 6412
rect 34756 6400 34762 6452
rect 35434 6400 35440 6452
rect 35492 6400 35498 6452
rect 37458 6400 37464 6452
rect 37516 6400 37522 6452
rect 37734 6400 37740 6452
rect 37792 6440 37798 6452
rect 37829 6443 37887 6449
rect 37829 6440 37841 6443
rect 37792 6412 37841 6440
rect 37792 6400 37798 6412
rect 37829 6409 37841 6412
rect 37875 6409 37887 6443
rect 37829 6403 37887 6409
rect 37918 6400 37924 6452
rect 37976 6400 37982 6452
rect 34514 6372 34520 6384
rect 34256 6344 34520 6372
rect 34149 6335 34207 6341
rect 34514 6332 34520 6344
rect 34572 6332 34578 6384
rect 30742 6264 30748 6316
rect 30800 6264 30806 6316
rect 33965 6307 34023 6313
rect 33965 6273 33977 6307
rect 34011 6304 34023 6307
rect 34238 6304 34244 6316
rect 34011 6276 34244 6304
rect 34011 6273 34023 6276
rect 33965 6267 34023 6273
rect 34238 6264 34244 6276
rect 34296 6264 34302 6316
rect 34790 6264 34796 6316
rect 34848 6264 34854 6316
rect 34882 6264 34888 6316
rect 34940 6304 34946 6316
rect 34977 6307 35035 6313
rect 34977 6304 34989 6307
rect 34940 6276 34989 6304
rect 34940 6264 34946 6276
rect 34977 6273 34989 6276
rect 35023 6273 35035 6307
rect 34977 6267 35035 6273
rect 35069 6307 35127 6313
rect 35069 6273 35081 6307
rect 35115 6273 35127 6307
rect 35069 6267 35127 6273
rect 35161 6307 35219 6313
rect 35161 6273 35173 6307
rect 35207 6304 35219 6307
rect 37734 6304 37740 6316
rect 35207 6276 37740 6304
rect 35207 6273 35219 6276
rect 35161 6267 35219 6273
rect 29411 6208 30696 6236
rect 29411 6205 29423 6208
rect 29365 6199 29423 6205
rect 30834 6196 30840 6248
rect 30892 6196 30898 6248
rect 31021 6239 31079 6245
rect 31021 6205 31033 6239
rect 31067 6236 31079 6239
rect 34606 6236 34612 6248
rect 31067 6208 34612 6236
rect 31067 6205 31079 6208
rect 31021 6199 31079 6205
rect 23860 6140 26234 6168
rect 20809 6131 20867 6137
rect 20990 6060 20996 6112
rect 21048 6100 21054 6112
rect 22005 6103 22063 6109
rect 22005 6100 22017 6103
rect 21048 6072 22017 6100
rect 21048 6060 21054 6072
rect 22005 6069 22017 6072
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 25498 6060 25504 6112
rect 25556 6100 25562 6112
rect 25777 6103 25835 6109
rect 25777 6100 25789 6103
rect 25556 6072 25789 6100
rect 25556 6060 25562 6072
rect 25777 6069 25789 6072
rect 25823 6069 25835 6103
rect 26206 6100 26234 6140
rect 29454 6128 29460 6180
rect 29512 6168 29518 6180
rect 31036 6168 31064 6199
rect 34606 6196 34612 6208
rect 34664 6236 34670 6248
rect 35084 6236 35112 6267
rect 37734 6264 37740 6276
rect 37792 6264 37798 6316
rect 34664 6208 35112 6236
rect 34664 6196 34670 6208
rect 38010 6196 38016 6248
rect 38068 6196 38074 6248
rect 29512 6140 31064 6168
rect 29512 6128 29518 6140
rect 28442 6100 28448 6112
rect 26206 6072 28448 6100
rect 25777 6063 25835 6069
rect 28442 6060 28448 6072
rect 28500 6060 28506 6112
rect 30006 6060 30012 6112
rect 30064 6100 30070 6112
rect 37826 6100 37832 6112
rect 30064 6072 37832 6100
rect 30064 6060 30070 6072
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 19242 5896 19248 5908
rect 18104 5868 19248 5896
rect 18104 5856 18110 5868
rect 19242 5856 19248 5868
rect 19300 5896 19306 5908
rect 19300 5868 19564 5896
rect 19300 5856 19306 5868
rect 19334 5828 19340 5840
rect 17328 5800 19340 5828
rect 16206 5720 16212 5772
rect 16264 5760 16270 5772
rect 16482 5760 16488 5772
rect 16264 5732 16488 5760
rect 16264 5720 16270 5732
rect 16482 5720 16488 5732
rect 16540 5760 16546 5772
rect 17328 5769 17356 5800
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 19536 5837 19564 5868
rect 22094 5856 22100 5908
rect 22152 5856 22158 5908
rect 25314 5856 25320 5908
rect 25372 5856 25378 5908
rect 25406 5856 25412 5908
rect 25464 5856 25470 5908
rect 27890 5856 27896 5908
rect 27948 5856 27954 5908
rect 30558 5856 30564 5908
rect 30616 5896 30622 5908
rect 30616 5868 35112 5896
rect 30616 5856 30622 5868
rect 19521 5831 19579 5837
rect 19521 5797 19533 5831
rect 19567 5797 19579 5831
rect 19521 5791 19579 5797
rect 17313 5763 17371 5769
rect 16540 5732 17080 5760
rect 16540 5720 16546 5732
rect 17052 5701 17080 5732
rect 17313 5729 17325 5763
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5760 17647 5763
rect 18046 5760 18052 5772
rect 17635 5732 18052 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5760 18199 5763
rect 19150 5760 19156 5772
rect 18187 5732 19156 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 19150 5720 19156 5732
rect 19208 5720 19214 5772
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19484 5732 19901 5760
rect 19484 5720 19490 5732
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 22186 5760 22192 5772
rect 20772 5732 22192 5760
rect 20772 5720 20778 5732
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 25498 5720 25504 5772
rect 25556 5720 25562 5772
rect 28166 5720 28172 5772
rect 28224 5760 28230 5772
rect 28353 5763 28411 5769
rect 28353 5760 28365 5763
rect 28224 5732 28365 5760
rect 28224 5720 28230 5732
rect 28353 5729 28365 5732
rect 28399 5729 28411 5763
rect 28353 5723 28411 5729
rect 28442 5720 28448 5772
rect 28500 5720 28506 5772
rect 32398 5720 32404 5772
rect 32456 5760 32462 5772
rect 33045 5763 33103 5769
rect 33045 5760 33057 5763
rect 32456 5732 33057 5760
rect 32456 5720 32462 5732
rect 33045 5729 33057 5732
rect 33091 5729 33103 5763
rect 33045 5723 33103 5729
rect 33134 5720 33140 5772
rect 33192 5720 33198 5772
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 17770 5652 17776 5704
rect 17828 5652 17834 5704
rect 20990 5652 20996 5704
rect 21048 5652 21054 5704
rect 25222 5652 25228 5704
rect 25280 5652 25286 5704
rect 28258 5652 28264 5704
rect 28316 5652 28322 5704
rect 29730 5652 29736 5704
rect 29788 5692 29794 5704
rect 30193 5695 30251 5701
rect 30193 5692 30205 5695
rect 29788 5664 30205 5692
rect 29788 5652 29794 5664
rect 30193 5661 30205 5664
rect 30239 5692 30251 5695
rect 31754 5692 31760 5704
rect 30239 5664 31760 5692
rect 30239 5661 30251 5664
rect 30193 5655 30251 5661
rect 31754 5652 31760 5664
rect 31812 5652 31818 5704
rect 32953 5695 33011 5701
rect 32953 5661 32965 5695
rect 32999 5692 33011 5695
rect 33686 5692 33692 5704
rect 32999 5664 33692 5692
rect 32999 5661 33011 5664
rect 32953 5655 33011 5661
rect 33686 5652 33692 5664
rect 33744 5692 33750 5704
rect 35084 5701 35112 5868
rect 35526 5856 35532 5908
rect 35584 5856 35590 5908
rect 33965 5695 34023 5701
rect 33965 5692 33977 5695
rect 33744 5664 33977 5692
rect 33744 5652 33750 5664
rect 33965 5661 33977 5664
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 34149 5695 34207 5701
rect 34149 5661 34161 5695
rect 34195 5692 34207 5695
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34195 5664 34897 5692
rect 34195 5661 34207 5664
rect 34149 5655 34207 5661
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35069 5695 35127 5701
rect 35069 5661 35081 5695
rect 35115 5661 35127 5695
rect 35069 5655 35127 5661
rect 35161 5695 35219 5701
rect 35161 5661 35173 5695
rect 35207 5661 35219 5695
rect 35161 5655 35219 5661
rect 35253 5695 35311 5701
rect 35253 5661 35265 5695
rect 35299 5692 35311 5695
rect 36446 5692 36452 5704
rect 35299 5664 36452 5692
rect 35299 5661 35311 5664
rect 35253 5655 35311 5661
rect 30466 5633 30472 5636
rect 30460 5587 30472 5633
rect 30466 5584 30472 5587
rect 30524 5584 30530 5636
rect 33781 5627 33839 5633
rect 33781 5593 33793 5627
rect 33827 5624 33839 5627
rect 34238 5624 34244 5636
rect 33827 5596 34244 5624
rect 33827 5593 33839 5596
rect 33781 5587 33839 5593
rect 34238 5584 34244 5596
rect 34296 5584 34302 5636
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 35176 5624 35204 5655
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 37826 5652 37832 5704
rect 37884 5652 37890 5704
rect 34572 5596 35204 5624
rect 34572 5584 34578 5596
rect 38102 5584 38108 5636
rect 38160 5584 38166 5636
rect 19426 5516 19432 5568
rect 19484 5516 19490 5568
rect 30742 5516 30748 5568
rect 30800 5556 30806 5568
rect 31573 5559 31631 5565
rect 31573 5556 31585 5559
rect 30800 5528 31585 5556
rect 30800 5516 30806 5528
rect 31573 5525 31585 5528
rect 31619 5525 31631 5559
rect 31573 5519 31631 5525
rect 32582 5516 32588 5568
rect 32640 5516 32646 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 23566 5312 23572 5364
rect 23624 5352 23630 5364
rect 24578 5352 24584 5364
rect 23624 5324 24584 5352
rect 23624 5312 23630 5324
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 30377 5355 30435 5361
rect 30377 5321 30389 5355
rect 30423 5352 30435 5355
rect 30466 5352 30472 5364
rect 30423 5324 30472 5352
rect 30423 5321 30435 5324
rect 30377 5315 30435 5321
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 30742 5312 30748 5364
rect 30800 5312 30806 5364
rect 33686 5312 33692 5364
rect 33744 5312 33750 5364
rect 34517 5355 34575 5361
rect 34517 5321 34529 5355
rect 34563 5352 34575 5355
rect 34790 5352 34796 5364
rect 34563 5324 34796 5352
rect 34563 5321 34575 5324
rect 34517 5315 34575 5321
rect 34790 5312 34796 5324
rect 34848 5312 34854 5364
rect 36446 5312 36452 5364
rect 36504 5312 36510 5364
rect 37734 5312 37740 5364
rect 37792 5352 37798 5364
rect 37829 5355 37887 5361
rect 37829 5352 37841 5355
rect 37792 5324 37841 5352
rect 37792 5312 37798 5324
rect 37829 5321 37841 5324
rect 37875 5321 37887 5355
rect 37829 5315 37887 5321
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 17129 5287 17187 5293
rect 17129 5284 17141 5287
rect 16724 5256 17141 5284
rect 16724 5244 16730 5256
rect 17129 5253 17141 5256
rect 17175 5253 17187 5287
rect 17129 5247 17187 5253
rect 20901 5287 20959 5293
rect 20901 5253 20913 5287
rect 20947 5284 20959 5287
rect 23474 5284 23480 5296
rect 20947 5256 23480 5284
rect 20947 5253 20959 5256
rect 20901 5247 20959 5253
rect 23474 5244 23480 5256
rect 23532 5244 23538 5296
rect 31754 5244 31760 5296
rect 31812 5284 31818 5296
rect 32950 5284 32956 5296
rect 31812 5256 32956 5284
rect 31812 5244 31818 5256
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 19245 5219 19303 5225
rect 19245 5216 19257 5219
rect 18831 5188 19257 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19245 5185 19257 5188
rect 19291 5216 19303 5219
rect 20714 5216 20720 5228
rect 19291 5188 20720 5216
rect 19291 5185 19303 5188
rect 19245 5179 19303 5185
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 22456 5219 22514 5225
rect 22456 5185 22468 5219
rect 22502 5216 22514 5219
rect 23014 5216 23020 5228
rect 22502 5188 23020 5216
rect 22502 5185 22514 5188
rect 22456 5179 22514 5185
rect 23014 5176 23020 5188
rect 23072 5176 23078 5228
rect 24857 5219 24915 5225
rect 24857 5185 24869 5219
rect 24903 5216 24915 5219
rect 25222 5216 25228 5228
rect 24903 5188 25228 5216
rect 24903 5185 24915 5188
rect 24857 5179 24915 5185
rect 25222 5176 25228 5188
rect 25280 5216 25286 5228
rect 25958 5216 25964 5228
rect 25280 5188 25964 5216
rect 25280 5176 25286 5188
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 30558 5216 30564 5228
rect 28224 5188 30564 5216
rect 28224 5176 28230 5188
rect 30558 5176 30564 5188
rect 30616 5216 30622 5228
rect 32324 5225 32352 5256
rect 32950 5244 32956 5256
rect 33008 5244 33014 5296
rect 34149 5287 34207 5293
rect 34149 5253 34161 5287
rect 34195 5284 34207 5287
rect 34238 5284 34244 5296
rect 34195 5256 34244 5284
rect 34195 5253 34207 5256
rect 34149 5247 34207 5253
rect 34238 5244 34244 5256
rect 34296 5244 34302 5296
rect 36814 5284 36820 5296
rect 35084 5256 36820 5284
rect 32582 5225 32588 5228
rect 30837 5219 30895 5225
rect 30837 5216 30849 5219
rect 30616 5188 30849 5216
rect 30616 5176 30622 5188
rect 30837 5185 30849 5188
rect 30883 5185 30895 5219
rect 30837 5179 30895 5185
rect 32309 5219 32367 5225
rect 32309 5185 32321 5219
rect 32355 5185 32367 5219
rect 32576 5216 32588 5225
rect 32543 5188 32588 5216
rect 32309 5179 32367 5185
rect 32576 5179 32588 5188
rect 32582 5176 32588 5179
rect 32640 5176 32646 5228
rect 34330 5176 34336 5228
rect 34388 5176 34394 5228
rect 35084 5225 35112 5256
rect 36814 5244 36820 5256
rect 36872 5244 36878 5296
rect 37642 5244 37648 5296
rect 37700 5284 37706 5296
rect 37921 5287 37979 5293
rect 37921 5284 37933 5287
rect 37700 5256 37933 5284
rect 37700 5244 37706 5256
rect 37921 5253 37933 5256
rect 37967 5253 37979 5287
rect 37921 5247 37979 5253
rect 35342 5225 35348 5228
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5185 35127 5219
rect 35069 5179 35127 5185
rect 35336 5179 35348 5225
rect 35342 5176 35348 5179
rect 35400 5176 35406 5228
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 19426 5148 19432 5160
rect 18555 5120 19432 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19518 5108 19524 5160
rect 19576 5108 19582 5160
rect 22186 5108 22192 5160
rect 22244 5108 22250 5160
rect 24946 5108 24952 5160
rect 25004 5108 25010 5160
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 30650 5148 30656 5160
rect 25096 5120 30656 5148
rect 25096 5108 25102 5120
rect 30650 5108 30656 5120
rect 30708 5148 30714 5160
rect 31021 5151 31079 5157
rect 31021 5148 31033 5151
rect 30708 5120 31033 5148
rect 30708 5108 30714 5120
rect 31021 5117 31033 5120
rect 31067 5148 31079 5151
rect 31202 5148 31208 5160
rect 31067 5120 31208 5148
rect 31067 5117 31079 5120
rect 31021 5111 31079 5117
rect 31202 5108 31208 5120
rect 31260 5108 31266 5160
rect 38010 5108 38016 5160
rect 38068 5108 38074 5160
rect 37550 5040 37556 5092
rect 37608 5080 37614 5092
rect 38028 5080 38056 5108
rect 37608 5052 38056 5080
rect 37608 5040 37614 5052
rect 24489 5015 24547 5021
rect 24489 4981 24501 5015
rect 24535 5012 24547 5015
rect 24670 5012 24676 5024
rect 24535 4984 24676 5012
rect 24535 4981 24547 4984
rect 24489 4975 24547 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 37458 4972 37464 5024
rect 37516 4972 37522 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 20070 4808 20076 4820
rect 17819 4780 20076 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 23014 4768 23020 4820
rect 23072 4768 23078 4820
rect 24596 4780 28948 4808
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 11112 4644 16221 4672
rect 11112 4632 11118 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 16482 4632 16488 4684
rect 16540 4632 16546 4684
rect 23661 4675 23719 4681
rect 23661 4641 23673 4675
rect 23707 4672 23719 4675
rect 24596 4672 24624 4780
rect 25958 4700 25964 4752
rect 26016 4700 26022 4752
rect 26050 4700 26056 4752
rect 26108 4740 26114 4752
rect 26421 4743 26479 4749
rect 26421 4740 26433 4743
rect 26108 4712 26433 4740
rect 26108 4700 26114 4712
rect 26421 4709 26433 4712
rect 26467 4709 26479 4743
rect 26421 4703 26479 4709
rect 23707 4644 24624 4672
rect 23707 4641 23719 4644
rect 23661 4635 23719 4641
rect 28166 4632 28172 4684
rect 28224 4672 28230 4684
rect 28920 4681 28948 4780
rect 30834 4768 30840 4820
rect 30892 4808 30898 4820
rect 31113 4811 31171 4817
rect 31113 4808 31125 4811
rect 30892 4780 31125 4808
rect 30892 4768 30898 4780
rect 31113 4777 31125 4780
rect 31159 4777 31171 4811
rect 31113 4771 31171 4777
rect 31202 4768 31208 4820
rect 31260 4808 31266 4820
rect 31260 4780 34284 4808
rect 31260 4768 31266 4780
rect 28721 4675 28779 4681
rect 28721 4672 28733 4675
rect 28224 4644 28733 4672
rect 28224 4632 28230 4644
rect 28721 4641 28733 4644
rect 28767 4641 28779 4675
rect 28721 4635 28779 4641
rect 28905 4675 28963 4681
rect 28905 4641 28917 4675
rect 28951 4672 28963 4675
rect 29178 4672 29184 4684
rect 28951 4644 29184 4672
rect 28951 4641 28963 4644
rect 28905 4635 28963 4641
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 29730 4632 29736 4684
rect 29788 4632 29794 4684
rect 32950 4632 32956 4684
rect 33008 4632 33014 4684
rect 34256 4672 34284 4780
rect 34330 4768 34336 4820
rect 34388 4768 34394 4820
rect 35342 4768 35348 4820
rect 35400 4808 35406 4820
rect 35529 4811 35587 4817
rect 35529 4808 35541 4811
rect 35400 4780 35541 4808
rect 35400 4768 35406 4780
rect 35529 4777 35541 4780
rect 35575 4777 35587 4811
rect 37550 4808 37556 4820
rect 35529 4771 35587 4777
rect 36096 4780 37556 4808
rect 36096 4681 36124 4780
rect 37550 4768 37556 4780
rect 37608 4768 37614 4820
rect 37734 4768 37740 4820
rect 37792 4808 37798 4820
rect 38197 4811 38255 4817
rect 38197 4808 38209 4811
rect 37792 4780 38209 4808
rect 37792 4768 37798 4780
rect 38197 4777 38209 4780
rect 38243 4777 38255 4811
rect 38197 4771 38255 4777
rect 36081 4675 36139 4681
rect 36081 4672 36093 4675
rect 34256 4644 36093 4672
rect 36081 4641 36093 4644
rect 36127 4641 36139 4675
rect 36081 4635 36139 4641
rect 36814 4632 36820 4684
rect 36872 4632 36878 4684
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 22244 4576 24593 4604
rect 22244 4564 22250 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 24670 4564 24676 4616
rect 24728 4604 24734 4616
rect 24837 4607 24895 4613
rect 24837 4604 24849 4607
rect 24728 4576 24849 4604
rect 24728 4564 24734 4576
rect 24837 4573 24849 4576
rect 24883 4573 24895 4607
rect 24837 4567 24895 4573
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27304 4576 27813 4604
rect 27304 4564 27310 4576
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 28626 4564 28632 4616
rect 28684 4564 28690 4616
rect 35897 4607 35955 4613
rect 35897 4573 35909 4607
rect 35943 4604 35955 4607
rect 36446 4604 36452 4616
rect 35943 4576 36452 4604
rect 35943 4573 35955 4576
rect 35897 4567 35955 4573
rect 36446 4564 36452 4576
rect 36504 4564 36510 4616
rect 37084 4607 37142 4613
rect 37084 4573 37096 4607
rect 37130 4604 37142 4607
rect 37458 4604 37464 4616
rect 37130 4576 37464 4604
rect 37130 4573 37142 4576
rect 37084 4567 37142 4573
rect 37458 4564 37464 4576
rect 37516 4564 37522 4616
rect 23385 4539 23443 4545
rect 23385 4505 23397 4539
rect 23431 4536 23443 4539
rect 23566 4536 23572 4548
rect 23431 4508 23572 4536
rect 23431 4505 23443 4508
rect 23385 4499 23443 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 26510 4496 26516 4548
rect 26568 4536 26574 4548
rect 27534 4539 27592 4545
rect 27534 4536 27546 4539
rect 26568 4508 27546 4536
rect 26568 4496 26574 4508
rect 27534 4505 27546 4508
rect 27580 4505 27592 4539
rect 27534 4499 27592 4505
rect 30000 4539 30058 4545
rect 30000 4505 30012 4539
rect 30046 4536 30058 4539
rect 30098 4536 30104 4548
rect 30046 4508 30104 4536
rect 30046 4505 30058 4508
rect 30000 4499 30058 4505
rect 30098 4496 30104 4508
rect 30156 4496 30162 4548
rect 33220 4539 33278 4545
rect 33220 4505 33232 4539
rect 33266 4536 33278 4539
rect 33410 4536 33416 4548
rect 33266 4508 33416 4536
rect 33266 4505 33278 4508
rect 33220 4499 33278 4505
rect 33410 4496 33416 4508
rect 33468 4496 33474 4548
rect 35986 4496 35992 4548
rect 36044 4496 36050 4548
rect 23477 4471 23535 4477
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 23658 4468 23664 4480
rect 23523 4440 23664 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 23658 4428 23664 4440
rect 23716 4468 23722 4480
rect 24946 4468 24952 4480
rect 23716 4440 24952 4468
rect 23716 4428 23722 4440
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 28258 4428 28264 4480
rect 28316 4428 28322 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 26050 4224 26056 4276
rect 26108 4264 26114 4276
rect 26145 4267 26203 4273
rect 26145 4264 26157 4267
rect 26108 4236 26157 4264
rect 26108 4224 26114 4236
rect 26145 4233 26157 4236
rect 26191 4233 26203 4267
rect 26145 4227 26203 4233
rect 26510 4224 26516 4276
rect 26568 4224 26574 4276
rect 28626 4224 28632 4276
rect 28684 4264 28690 4276
rect 28905 4267 28963 4273
rect 28905 4264 28917 4267
rect 28684 4236 28917 4264
rect 28684 4224 28690 4236
rect 28905 4233 28917 4236
rect 28951 4233 28963 4267
rect 28905 4227 28963 4233
rect 30098 4224 30104 4276
rect 30156 4224 30162 4276
rect 30469 4267 30527 4273
rect 30469 4233 30481 4267
rect 30515 4264 30527 4267
rect 30834 4264 30840 4276
rect 30515 4236 30840 4264
rect 30515 4233 30527 4236
rect 30469 4227 30527 4233
rect 30834 4224 30840 4236
rect 30892 4224 30898 4276
rect 33410 4224 33416 4276
rect 33468 4224 33474 4276
rect 33781 4267 33839 4273
rect 33781 4233 33793 4267
rect 33827 4264 33839 4267
rect 34330 4264 34336 4276
rect 33827 4236 34336 4264
rect 33827 4233 33839 4236
rect 33781 4227 33839 4233
rect 34330 4224 34336 4236
rect 34388 4224 34394 4276
rect 27792 4199 27850 4205
rect 27792 4165 27804 4199
rect 27838 4196 27850 4199
rect 28258 4196 28264 4208
rect 27838 4168 28264 4196
rect 27838 4165 27850 4168
rect 27792 4159 27850 4165
rect 28258 4156 28264 4168
rect 28316 4156 28322 4208
rect 30558 4156 30564 4208
rect 30616 4156 30622 4208
rect 24946 4088 24952 4140
rect 25004 4128 25010 4140
rect 26053 4131 26111 4137
rect 26053 4128 26065 4131
rect 25004 4100 26065 4128
rect 25004 4088 25010 4100
rect 26053 4097 26065 4100
rect 26099 4097 26111 4131
rect 26053 4091 26111 4097
rect 27246 4088 27252 4140
rect 27304 4128 27310 4140
rect 27525 4131 27583 4137
rect 27525 4128 27537 4131
rect 27304 4100 27537 4128
rect 27304 4088 27310 4100
rect 27525 4097 27537 4100
rect 27571 4097 27583 4131
rect 27525 4091 27583 4097
rect 33870 4088 33876 4140
rect 33928 4088 33934 4140
rect 37829 4131 37887 4137
rect 37829 4097 37841 4131
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 38105 4131 38163 4137
rect 38105 4097 38117 4131
rect 38151 4128 38163 4131
rect 39022 4128 39028 4140
rect 38151 4100 39028 4128
rect 38151 4097 38163 4100
rect 38105 4091 38163 4097
rect 25866 4020 25872 4072
rect 25924 4020 25930 4072
rect 30745 4063 30803 4069
rect 30745 4029 30757 4063
rect 30791 4029 30803 4063
rect 30745 4023 30803 4029
rect 33965 4063 34023 4069
rect 33965 4029 33977 4063
rect 34011 4029 34023 4063
rect 33965 4023 34023 4029
rect 30760 3992 30788 4023
rect 33134 3992 33140 4004
rect 30760 3964 33140 3992
rect 33134 3952 33140 3964
rect 33192 3992 33198 4004
rect 33980 3992 34008 4023
rect 33192 3964 34008 3992
rect 33192 3952 33198 3964
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 37844 3924 37872 4091
rect 39022 4088 39028 4100
rect 39080 4088 39086 4140
rect 29696 3896 37872 3924
rect 29696 3884 29702 3896
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 37826 3000 37832 3052
rect 37884 3000 37890 3052
rect 38102 2932 38108 2984
rect 38160 2932 38166 2984
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 37829 2431 37887 2437
rect 37829 2428 37841 2431
rect 28132 2400 37841 2428
rect 28132 2388 28138 2400
rect 37829 2397 37841 2400
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38102 2320 38108 2372
rect 38160 2320 38166 2372
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 5080 39108 5132 39160
rect 6644 39108 6696 39160
rect 21640 39108 21692 39160
rect 22100 39108 22152 39160
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5816 37315 5868 37324
rect 5816 37281 5825 37315
rect 5825 37281 5859 37315
rect 5859 37281 5868 37315
rect 5816 37272 5868 37281
rect 9312 37272 9364 37324
rect 36636 37272 36688 37324
rect 39028 37272 39080 37324
rect 1768 37204 1820 37256
rect 6644 37247 6696 37256
rect 6644 37213 6653 37247
rect 6653 37213 6687 37247
rect 6687 37213 6696 37247
rect 6644 37204 6696 37213
rect 8392 37204 8444 37256
rect 11704 37204 11756 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 18328 37204 18380 37256
rect 5540 37179 5592 37188
rect 5540 37145 5549 37179
rect 5549 37145 5583 37179
rect 5583 37145 5592 37179
rect 5540 37136 5592 37145
rect 7012 37179 7064 37188
rect 7012 37145 7021 37179
rect 7021 37145 7055 37179
rect 7055 37145 7064 37179
rect 7012 37136 7064 37145
rect 7380 37136 7432 37188
rect 9680 37136 9732 37188
rect 5172 37111 5224 37120
rect 5172 37077 5181 37111
rect 5181 37077 5215 37111
rect 5215 37077 5224 37111
rect 5172 37068 5224 37077
rect 5632 37111 5684 37120
rect 5632 37077 5641 37111
rect 5641 37077 5675 37111
rect 5675 37077 5684 37111
rect 5632 37068 5684 37077
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 9588 37111 9640 37120
rect 9588 37077 9597 37111
rect 9597 37077 9631 37111
rect 9631 37077 9640 37111
rect 9588 37068 9640 37077
rect 12072 37136 12124 37188
rect 16212 37136 16264 37188
rect 18788 37179 18840 37188
rect 18788 37145 18797 37179
rect 18797 37145 18831 37179
rect 18831 37145 18840 37179
rect 18788 37136 18840 37145
rect 20168 37247 20220 37256
rect 20168 37213 20177 37247
rect 20177 37213 20211 37247
rect 20211 37213 20220 37247
rect 20168 37204 20220 37213
rect 22100 37247 22152 37256
rect 22100 37213 22109 37247
rect 22109 37213 22143 37247
rect 22143 37213 22152 37247
rect 22100 37204 22152 37213
rect 24952 37204 25004 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 27712 37204 27764 37256
rect 28264 37204 28316 37256
rect 31760 37204 31812 37256
rect 36912 37247 36964 37256
rect 36912 37213 36921 37247
rect 36921 37213 36955 37247
rect 36955 37213 36964 37247
rect 36912 37204 36964 37213
rect 38200 37247 38252 37256
rect 38200 37213 38209 37247
rect 38209 37213 38243 37247
rect 38243 37213 38252 37247
rect 38200 37204 38252 37213
rect 17040 37068 17092 37120
rect 19432 37068 19484 37120
rect 20996 37136 21048 37188
rect 22284 37136 22336 37188
rect 22928 37136 22980 37188
rect 31024 37136 31076 37188
rect 31852 37136 31904 37188
rect 23664 37068 23716 37120
rect 26608 37068 26660 37120
rect 28540 37111 28592 37120
rect 28540 37077 28549 37111
rect 28549 37077 28583 37111
rect 28583 37077 28592 37111
rect 28540 37068 28592 37077
rect 36820 37136 36872 37188
rect 39028 37068 39080 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 5632 36864 5684 36916
rect 9588 36907 9640 36916
rect 9588 36873 9597 36907
rect 9597 36873 9631 36907
rect 9631 36873 9640 36907
rect 9588 36864 9640 36873
rect 11060 36864 11112 36916
rect 14188 36864 14240 36916
rect 5172 36796 5224 36848
rect 9128 36796 9180 36848
rect 13176 36771 13228 36780
rect 13176 36737 13194 36771
rect 13194 36737 13228 36771
rect 13176 36728 13228 36737
rect 13360 36728 13412 36780
rect 15200 36796 15252 36848
rect 15936 36796 15988 36848
rect 17040 36771 17092 36780
rect 17040 36737 17049 36771
rect 17049 36737 17083 36771
rect 17083 36737 17092 36771
rect 17040 36728 17092 36737
rect 19432 36796 19484 36848
rect 20628 36728 20680 36780
rect 20996 36771 21048 36780
rect 20996 36737 21005 36771
rect 21005 36737 21039 36771
rect 21039 36737 21048 36771
rect 20996 36728 21048 36737
rect 21548 36728 21600 36780
rect 4620 36703 4672 36712
rect 4620 36669 4629 36703
rect 4629 36669 4663 36703
rect 4663 36669 4672 36703
rect 4620 36660 4672 36669
rect 14556 36703 14608 36712
rect 14556 36669 14565 36703
rect 14565 36669 14599 36703
rect 14599 36669 14608 36703
rect 14556 36660 14608 36669
rect 15108 36660 15160 36712
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 19984 36703 20036 36712
rect 19984 36669 19993 36703
rect 19993 36669 20027 36703
rect 20027 36669 20036 36703
rect 19984 36660 20036 36669
rect 23756 36796 23808 36848
rect 25596 36796 25648 36848
rect 22376 36771 22428 36780
rect 22376 36737 22410 36771
rect 22410 36737 22428 36771
rect 22376 36728 22428 36737
rect 26332 36771 26384 36780
rect 26332 36737 26341 36771
rect 26341 36737 26375 36771
rect 26375 36737 26384 36771
rect 26332 36728 26384 36737
rect 26608 36771 26660 36780
rect 26608 36737 26617 36771
rect 26617 36737 26651 36771
rect 26651 36737 26660 36771
rect 26608 36728 26660 36737
rect 28816 36796 28868 36848
rect 24860 36660 24912 36712
rect 26148 36660 26200 36712
rect 28264 36728 28316 36780
rect 32772 36796 32824 36848
rect 32404 36728 32456 36780
rect 33968 36728 34020 36780
rect 36728 36728 36780 36780
rect 37924 36728 37976 36780
rect 31852 36660 31904 36712
rect 34244 36660 34296 36712
rect 36636 36703 36688 36712
rect 36636 36669 36645 36703
rect 36645 36669 36679 36703
rect 36679 36669 36688 36703
rect 36636 36660 36688 36669
rect 39028 36660 39080 36712
rect 9128 36524 9180 36576
rect 12716 36524 12768 36576
rect 16028 36567 16080 36576
rect 16028 36533 16037 36567
rect 16037 36533 16071 36567
rect 16071 36533 16080 36567
rect 16028 36524 16080 36533
rect 16948 36567 17000 36576
rect 16948 36533 16957 36567
rect 16957 36533 16991 36567
rect 16991 36533 17000 36567
rect 16948 36524 17000 36533
rect 20168 36524 20220 36576
rect 20536 36524 20588 36576
rect 23020 36524 23072 36576
rect 26424 36524 26476 36576
rect 28724 36524 28776 36576
rect 30104 36524 30156 36576
rect 33416 36524 33468 36576
rect 35716 36567 35768 36576
rect 35716 36533 35725 36567
rect 35725 36533 35759 36567
rect 35759 36533 35768 36567
rect 35716 36524 35768 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 13176 36320 13228 36372
rect 15200 36363 15252 36372
rect 15200 36329 15209 36363
rect 15209 36329 15243 36363
rect 15243 36329 15252 36363
rect 15200 36320 15252 36329
rect 9220 36295 9272 36304
rect 9220 36261 9229 36295
rect 9229 36261 9263 36295
rect 9263 36261 9272 36295
rect 9220 36252 9272 36261
rect 14188 36252 14240 36304
rect 5632 36184 5684 36236
rect 5908 36227 5960 36236
rect 5908 36193 5917 36227
rect 5917 36193 5951 36227
rect 5951 36193 5960 36227
rect 5908 36184 5960 36193
rect 9680 36184 9732 36236
rect 12900 36227 12952 36236
rect 12900 36193 12909 36227
rect 12909 36193 12943 36227
rect 12943 36193 12952 36227
rect 12900 36184 12952 36193
rect 15936 36184 15988 36236
rect 16028 36184 16080 36236
rect 22284 36320 22336 36372
rect 24952 36320 25004 36372
rect 25596 36363 25648 36372
rect 25596 36329 25605 36363
rect 25605 36329 25639 36363
rect 25639 36329 25648 36363
rect 25596 36320 25648 36329
rect 18972 36252 19024 36304
rect 21272 36252 21324 36304
rect 27160 36320 27212 36372
rect 28264 36363 28316 36372
rect 28264 36329 28273 36363
rect 28273 36329 28307 36363
rect 28307 36329 28316 36363
rect 28264 36320 28316 36329
rect 30104 36363 30156 36372
rect 30104 36329 30113 36363
rect 30113 36329 30147 36363
rect 30147 36329 30156 36363
rect 30104 36320 30156 36329
rect 32404 36320 32456 36372
rect 33968 36363 34020 36372
rect 33968 36329 33977 36363
rect 33977 36329 34011 36363
rect 34011 36329 34020 36363
rect 33968 36320 34020 36329
rect 36820 36320 36872 36372
rect 4620 36116 4672 36168
rect 9128 36116 9180 36168
rect 12716 36116 12768 36168
rect 13268 36116 13320 36168
rect 15108 36159 15160 36168
rect 15108 36125 15117 36159
rect 15117 36125 15151 36159
rect 15151 36125 15160 36159
rect 15108 36116 15160 36125
rect 16120 36159 16172 36168
rect 16120 36125 16129 36159
rect 16129 36125 16163 36159
rect 16163 36125 16172 36159
rect 16120 36116 16172 36125
rect 5540 36048 5592 36100
rect 7104 36048 7156 36100
rect 9588 36048 9640 36100
rect 10140 36048 10192 36100
rect 11704 36048 11756 36100
rect 16948 36048 17000 36100
rect 5264 36023 5316 36032
rect 5264 35989 5273 36023
rect 5273 35989 5307 36023
rect 5307 35989 5316 36023
rect 5264 35980 5316 35989
rect 7840 36023 7892 36032
rect 7840 35989 7849 36023
rect 7849 35989 7883 36023
rect 7883 35989 7892 36023
rect 7840 35980 7892 35989
rect 11888 36023 11940 36032
rect 11888 35989 11897 36023
rect 11897 35989 11931 36023
rect 11931 35989 11940 36023
rect 11888 35980 11940 35989
rect 13452 35980 13504 36032
rect 18696 36048 18748 36100
rect 18972 36048 19024 36100
rect 20260 36116 20312 36168
rect 20352 36116 20404 36168
rect 20720 36159 20772 36168
rect 20720 36125 20729 36159
rect 20729 36125 20763 36159
rect 20763 36125 20772 36159
rect 20720 36116 20772 36125
rect 22284 36184 22336 36236
rect 22468 36184 22520 36236
rect 26148 36227 26200 36236
rect 26148 36193 26157 36227
rect 26157 36193 26191 36227
rect 26191 36193 26200 36227
rect 26148 36184 26200 36193
rect 26332 36184 26384 36236
rect 26424 36227 26476 36236
rect 26424 36193 26433 36227
rect 26433 36193 26467 36227
rect 26467 36193 26476 36227
rect 26424 36184 26476 36193
rect 23020 36116 23072 36168
rect 23388 36116 23440 36168
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 23664 36048 23716 36100
rect 31484 36227 31536 36236
rect 31484 36193 31493 36227
rect 31493 36193 31527 36227
rect 31527 36193 31536 36227
rect 31484 36184 31536 36193
rect 24860 36091 24912 36100
rect 24860 36057 24869 36091
rect 24869 36057 24903 36091
rect 24903 36057 24912 36091
rect 24860 36048 24912 36057
rect 27712 36048 27764 36100
rect 30196 36159 30248 36168
rect 30196 36125 30205 36159
rect 30205 36125 30239 36159
rect 30239 36125 30248 36159
rect 30196 36116 30248 36125
rect 33048 36184 33100 36236
rect 34244 36184 34296 36236
rect 32680 36116 32732 36168
rect 31852 36048 31904 36100
rect 32496 36048 32548 36100
rect 36360 36116 36412 36168
rect 34520 36048 34572 36100
rect 37464 36048 37516 36100
rect 19432 35980 19484 36032
rect 20444 36023 20496 36032
rect 20444 35989 20453 36023
rect 20453 35989 20487 36023
rect 20487 35989 20496 36023
rect 20444 35980 20496 35989
rect 22928 35980 22980 36032
rect 28724 35980 28776 36032
rect 29184 35980 29236 36032
rect 36084 35980 36136 36032
rect 37832 35980 37884 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 7104 35819 7156 35828
rect 7104 35785 7113 35819
rect 7113 35785 7147 35819
rect 7147 35785 7156 35819
rect 7104 35776 7156 35785
rect 7564 35819 7616 35828
rect 7564 35785 7573 35819
rect 7573 35785 7607 35819
rect 7607 35785 7616 35819
rect 7564 35776 7616 35785
rect 7840 35776 7892 35828
rect 11704 35819 11756 35828
rect 11704 35785 11713 35819
rect 11713 35785 11747 35819
rect 11747 35785 11756 35819
rect 11704 35776 11756 35785
rect 18420 35776 18472 35828
rect 20720 35776 20772 35828
rect 21364 35776 21416 35828
rect 22376 35776 22428 35828
rect 23020 35776 23072 35828
rect 33048 35776 33100 35828
rect 34520 35776 34572 35828
rect 36912 35776 36964 35828
rect 37464 35819 37516 35828
rect 37464 35785 37473 35819
rect 37473 35785 37507 35819
rect 37507 35785 37516 35819
rect 37464 35776 37516 35785
rect 7472 35683 7524 35692
rect 7472 35649 7481 35683
rect 7481 35649 7515 35683
rect 7515 35649 7524 35683
rect 7472 35640 7524 35649
rect 5816 35572 5868 35624
rect 9312 35708 9364 35760
rect 9864 35683 9916 35692
rect 9864 35649 9873 35683
rect 9873 35649 9907 35683
rect 9907 35649 9916 35683
rect 9864 35640 9916 35649
rect 9956 35615 10008 35624
rect 9956 35581 9965 35615
rect 9965 35581 9999 35615
rect 9999 35581 10008 35615
rect 9956 35572 10008 35581
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 11796 35572 11848 35624
rect 12900 35708 12952 35760
rect 15108 35640 15160 35692
rect 17040 35683 17092 35692
rect 17040 35649 17049 35683
rect 17049 35649 17083 35683
rect 17083 35649 17092 35683
rect 17040 35640 17092 35649
rect 18420 35640 18472 35692
rect 18604 35683 18656 35692
rect 18604 35649 18613 35683
rect 18613 35649 18647 35683
rect 18647 35649 18656 35683
rect 18604 35640 18656 35649
rect 18972 35683 19024 35692
rect 18972 35649 18981 35683
rect 18981 35649 19015 35683
rect 19015 35649 19024 35683
rect 18972 35640 19024 35649
rect 18696 35572 18748 35624
rect 20352 35640 20404 35692
rect 20536 35683 20588 35692
rect 20536 35649 20545 35683
rect 20545 35649 20579 35683
rect 20579 35649 20588 35683
rect 20536 35640 20588 35649
rect 21272 35708 21324 35760
rect 23388 35708 23440 35760
rect 23572 35708 23624 35760
rect 20812 35615 20864 35624
rect 20812 35581 20821 35615
rect 20821 35581 20855 35615
rect 20855 35581 20864 35615
rect 20812 35572 20864 35581
rect 9864 35504 9916 35556
rect 16212 35504 16264 35556
rect 22928 35640 22980 35692
rect 23664 35683 23716 35692
rect 23664 35649 23673 35683
rect 23673 35649 23707 35683
rect 23707 35649 23716 35683
rect 23664 35640 23716 35649
rect 23756 35640 23808 35692
rect 25228 35640 25280 35692
rect 25136 35572 25188 35624
rect 25504 35615 25556 35624
rect 25504 35581 25513 35615
rect 25513 35581 25547 35615
rect 25547 35581 25556 35615
rect 25504 35572 25556 35581
rect 27252 35683 27304 35692
rect 27252 35649 27261 35683
rect 27261 35649 27295 35683
rect 27295 35649 27304 35683
rect 27252 35640 27304 35649
rect 28816 35683 28868 35692
rect 28816 35649 28825 35683
rect 28825 35649 28859 35683
rect 28859 35649 28868 35683
rect 28816 35640 28868 35649
rect 29092 35683 29144 35692
rect 29092 35649 29126 35683
rect 29126 35649 29144 35683
rect 29092 35640 29144 35649
rect 32496 35683 32548 35692
rect 32496 35649 32505 35683
rect 32505 35649 32539 35683
rect 32539 35649 32548 35683
rect 32496 35640 32548 35649
rect 32680 35683 32732 35692
rect 32680 35649 32689 35683
rect 32689 35649 32723 35683
rect 32723 35649 32732 35683
rect 32680 35640 32732 35649
rect 33508 35683 33560 35692
rect 33508 35649 33517 35683
rect 33517 35649 33551 35683
rect 33551 35649 33560 35683
rect 33508 35640 33560 35649
rect 36728 35683 36780 35692
rect 36728 35649 36737 35683
rect 36737 35649 36771 35683
rect 36771 35649 36780 35683
rect 36728 35640 36780 35649
rect 37648 35640 37700 35692
rect 37832 35683 37884 35692
rect 37832 35649 37841 35683
rect 37841 35649 37875 35683
rect 37875 35649 37884 35683
rect 37832 35640 37884 35649
rect 27712 35615 27764 35624
rect 27712 35581 27721 35615
rect 27721 35581 27755 35615
rect 27755 35581 27764 35615
rect 27712 35572 27764 35581
rect 37924 35615 37976 35624
rect 37924 35581 37933 35615
rect 37933 35581 37967 35615
rect 37967 35581 37976 35615
rect 37924 35572 37976 35581
rect 38016 35615 38068 35624
rect 38016 35581 38025 35615
rect 38025 35581 38059 35615
rect 38059 35581 38068 35615
rect 38016 35572 38068 35581
rect 26056 35504 26108 35556
rect 9404 35436 9456 35488
rect 14740 35436 14792 35488
rect 16948 35479 17000 35488
rect 16948 35445 16957 35479
rect 16957 35445 16991 35479
rect 16991 35445 17000 35479
rect 16948 35436 17000 35445
rect 18236 35479 18288 35488
rect 18236 35445 18245 35479
rect 18245 35445 18279 35479
rect 18279 35445 18288 35479
rect 18236 35436 18288 35445
rect 23388 35436 23440 35488
rect 25044 35479 25096 35488
rect 25044 35445 25053 35479
rect 25053 35445 25087 35479
rect 25087 35445 25096 35479
rect 25044 35436 25096 35445
rect 30196 35479 30248 35488
rect 30196 35445 30205 35479
rect 30205 35445 30239 35479
rect 30239 35445 30248 35479
rect 30196 35436 30248 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 10600 35164 10652 35216
rect 5816 35139 5868 35148
rect 5816 35105 5825 35139
rect 5825 35105 5859 35139
rect 5859 35105 5868 35139
rect 5816 35096 5868 35105
rect 12072 35096 12124 35148
rect 13452 35096 13504 35148
rect 15936 35096 15988 35148
rect 16212 35096 16264 35148
rect 9128 35071 9180 35080
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 9404 35071 9456 35080
rect 9404 35037 9438 35071
rect 9438 35037 9456 35071
rect 9404 35028 9456 35037
rect 10140 35028 10192 35080
rect 6368 34960 6420 35012
rect 7012 34960 7064 35012
rect 11796 35003 11848 35012
rect 11796 34969 11805 35003
rect 11805 34969 11839 35003
rect 11839 34969 11848 35003
rect 11796 34960 11848 34969
rect 12624 35003 12676 35012
rect 12624 34969 12633 35003
rect 12633 34969 12667 35003
rect 12667 34969 12676 35003
rect 12624 34960 12676 34969
rect 5172 34935 5224 34944
rect 5172 34901 5181 34935
rect 5181 34901 5215 34935
rect 5215 34901 5224 34935
rect 5172 34892 5224 34901
rect 5632 34935 5684 34944
rect 5632 34901 5641 34935
rect 5641 34901 5675 34935
rect 5675 34901 5684 34935
rect 5632 34892 5684 34901
rect 9956 34892 10008 34944
rect 13268 35071 13320 35080
rect 13268 35037 13277 35071
rect 13277 35037 13311 35071
rect 13311 35037 13320 35071
rect 13268 35028 13320 35037
rect 16948 35028 17000 35080
rect 15844 35003 15896 35012
rect 15844 34969 15853 35003
rect 15853 34969 15887 35003
rect 15887 34969 15896 35003
rect 15844 34960 15896 34969
rect 22468 35164 22520 35216
rect 20260 35096 20312 35148
rect 17960 35028 18012 35080
rect 18328 35028 18380 35080
rect 18604 35028 18656 35080
rect 18696 35003 18748 35012
rect 18696 34969 18730 35003
rect 18730 34969 18748 35003
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 21088 35096 21140 35148
rect 20444 35071 20496 35080
rect 20444 35037 20453 35071
rect 20453 35037 20487 35071
rect 20487 35037 20496 35071
rect 20444 35028 20496 35037
rect 20628 35071 20680 35080
rect 20628 35037 20637 35071
rect 20637 35037 20671 35071
rect 20671 35037 20680 35071
rect 20628 35028 20680 35037
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 25228 35232 25280 35284
rect 25964 35232 26016 35284
rect 23480 35207 23532 35216
rect 23480 35173 23489 35207
rect 23489 35173 23523 35207
rect 23523 35173 23532 35207
rect 23480 35164 23532 35173
rect 24860 35164 24912 35216
rect 25504 35164 25556 35216
rect 27344 35164 27396 35216
rect 29092 35275 29144 35284
rect 29092 35241 29101 35275
rect 29101 35241 29135 35275
rect 29135 35241 29144 35275
rect 29092 35232 29144 35241
rect 32496 35232 32548 35284
rect 33508 35232 33560 35284
rect 31208 35164 31260 35216
rect 23664 35028 23716 35080
rect 23848 35071 23900 35080
rect 23848 35037 23857 35071
rect 23857 35037 23891 35071
rect 23891 35037 23900 35071
rect 23848 35028 23900 35037
rect 25228 35096 25280 35148
rect 26148 35096 26200 35148
rect 18696 34960 18748 34969
rect 20536 35003 20588 35012
rect 20536 34969 20545 35003
rect 20545 34969 20579 35003
rect 20579 34969 20588 35003
rect 20536 34960 20588 34969
rect 21180 34960 21232 35012
rect 18420 34892 18472 34944
rect 20352 34892 20404 34944
rect 23020 35003 23072 35012
rect 23020 34969 23029 35003
rect 23029 34969 23063 35003
rect 23063 34969 23072 35003
rect 23020 34960 23072 34969
rect 23388 34892 23440 34944
rect 25136 35028 25188 35080
rect 26608 35071 26660 35080
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26608 35028 26660 35037
rect 29184 35139 29236 35148
rect 29184 35105 29193 35139
rect 29193 35105 29227 35139
rect 29227 35105 29236 35139
rect 29184 35096 29236 35105
rect 28908 35071 28960 35080
rect 28908 35037 28917 35071
rect 28917 35037 28951 35071
rect 28951 35037 28960 35071
rect 28908 35028 28960 35037
rect 29276 35028 29328 35080
rect 30840 35071 30892 35080
rect 30840 35037 30849 35071
rect 30849 35037 30883 35071
rect 30883 35037 30892 35071
rect 30840 35028 30892 35037
rect 30932 35071 30984 35080
rect 30932 35037 30942 35071
rect 30942 35037 30976 35071
rect 30976 35037 30984 35071
rect 35716 35096 35768 35148
rect 35900 35096 35952 35148
rect 36360 35139 36412 35148
rect 36360 35105 36369 35139
rect 36369 35105 36403 35139
rect 36403 35105 36412 35139
rect 36360 35096 36412 35105
rect 30932 35028 30984 35037
rect 31576 35028 31628 35080
rect 32956 35071 33008 35080
rect 32956 35037 32965 35071
rect 32965 35037 32999 35071
rect 32999 35037 33008 35071
rect 32956 35028 33008 35037
rect 24860 34892 24912 34944
rect 25504 34960 25556 35012
rect 26056 34960 26108 35012
rect 26884 35003 26936 35012
rect 26884 34969 26893 35003
rect 26893 34969 26927 35003
rect 26927 34969 26936 35003
rect 26884 34960 26936 34969
rect 25044 34892 25096 34944
rect 25596 34892 25648 34944
rect 25688 34935 25740 34944
rect 25688 34901 25697 34935
rect 25697 34901 25731 34935
rect 25731 34901 25740 34935
rect 25688 34892 25740 34901
rect 28632 34892 28684 34944
rect 30932 34892 30984 34944
rect 31208 35003 31260 35012
rect 31208 34969 31217 35003
rect 31217 34969 31251 35003
rect 31251 34969 31260 35003
rect 31208 34960 31260 34969
rect 32496 34960 32548 35012
rect 34796 34960 34848 35012
rect 37464 34960 37516 35012
rect 33048 34892 33100 34944
rect 37740 34935 37792 34944
rect 37740 34901 37749 34935
rect 37749 34901 37783 34935
rect 37783 34901 37792 34935
rect 37740 34892 37792 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4620 34688 4672 34740
rect 5632 34688 5684 34740
rect 7104 34688 7156 34740
rect 9864 34731 9916 34740
rect 9864 34697 9873 34731
rect 9873 34697 9907 34731
rect 9907 34697 9916 34731
rect 9864 34688 9916 34697
rect 9956 34731 10008 34740
rect 9956 34697 9965 34731
rect 9965 34697 9999 34731
rect 9999 34697 10008 34731
rect 9956 34688 10008 34697
rect 20076 34688 20128 34740
rect 5540 34620 5592 34672
rect 5908 34620 5960 34672
rect 20628 34688 20680 34740
rect 22100 34688 22152 34740
rect 24492 34688 24544 34740
rect 27252 34688 27304 34740
rect 28908 34688 28960 34740
rect 31484 34688 31536 34740
rect 5172 34552 5224 34604
rect 7564 34595 7616 34604
rect 7564 34561 7573 34595
rect 7573 34561 7607 34595
rect 7607 34561 7616 34595
rect 7564 34552 7616 34561
rect 13360 34595 13412 34604
rect 13360 34561 13369 34595
rect 13369 34561 13403 34595
rect 13403 34561 13412 34595
rect 13360 34552 13412 34561
rect 14740 34552 14792 34604
rect 19984 34595 20036 34604
rect 19984 34561 19993 34595
rect 19993 34561 20027 34595
rect 20027 34561 20036 34595
rect 19984 34552 20036 34561
rect 20444 34620 20496 34672
rect 20628 34552 20680 34604
rect 21088 34595 21140 34604
rect 21088 34561 21097 34595
rect 21097 34561 21131 34595
rect 21131 34561 21140 34595
rect 21088 34552 21140 34561
rect 7472 34527 7524 34536
rect 7472 34493 7481 34527
rect 7481 34493 7515 34527
rect 7515 34493 7524 34527
rect 7472 34484 7524 34493
rect 7932 34484 7984 34536
rect 8208 34527 8260 34536
rect 8208 34493 8217 34527
rect 8217 34493 8251 34527
rect 8251 34493 8260 34527
rect 8208 34484 8260 34493
rect 10140 34527 10192 34536
rect 10140 34493 10149 34527
rect 10149 34493 10183 34527
rect 10183 34493 10192 34527
rect 10140 34484 10192 34493
rect 12072 34484 12124 34536
rect 13176 34484 13228 34536
rect 13636 34527 13688 34536
rect 13636 34493 13645 34527
rect 13645 34493 13679 34527
rect 13679 34493 13688 34527
rect 13636 34484 13688 34493
rect 15016 34484 15068 34536
rect 20352 34484 20404 34536
rect 20536 34484 20588 34536
rect 20812 34484 20864 34536
rect 26148 34620 26200 34672
rect 21272 34595 21324 34604
rect 21272 34561 21281 34595
rect 21281 34561 21315 34595
rect 21315 34561 21324 34595
rect 21272 34552 21324 34561
rect 21364 34552 21416 34604
rect 25044 34552 25096 34604
rect 25136 34595 25188 34604
rect 25136 34561 25145 34595
rect 25145 34561 25179 34595
rect 25179 34561 25188 34595
rect 25136 34552 25188 34561
rect 26056 34552 26108 34604
rect 26884 34620 26936 34672
rect 29460 34595 29512 34604
rect 29460 34561 29469 34595
rect 29469 34561 29503 34595
rect 29503 34561 29512 34595
rect 29460 34552 29512 34561
rect 30196 34595 30248 34604
rect 30196 34561 30205 34595
rect 30205 34561 30239 34595
rect 30239 34561 30248 34595
rect 30196 34552 30248 34561
rect 30656 34595 30708 34604
rect 30656 34561 30665 34595
rect 30665 34561 30699 34595
rect 30699 34561 30708 34595
rect 30656 34552 30708 34561
rect 30748 34595 30800 34604
rect 30748 34561 30758 34595
rect 30758 34561 30792 34595
rect 30792 34561 30800 34595
rect 30748 34552 30800 34561
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 31024 34595 31076 34604
rect 31024 34561 31033 34595
rect 31033 34561 31067 34595
rect 31067 34561 31076 34595
rect 31024 34552 31076 34561
rect 31576 34552 31628 34604
rect 32496 34663 32548 34672
rect 32496 34629 32521 34663
rect 32521 34629 32548 34663
rect 32680 34731 32732 34740
rect 32680 34697 32689 34731
rect 32689 34697 32723 34731
rect 32723 34697 32732 34731
rect 32680 34688 32732 34697
rect 37464 34731 37516 34740
rect 37464 34697 37473 34731
rect 37473 34697 37507 34731
rect 37507 34697 37516 34731
rect 37464 34688 37516 34697
rect 32496 34620 32548 34629
rect 33416 34620 33468 34672
rect 33048 34552 33100 34604
rect 34244 34595 34296 34604
rect 34244 34561 34253 34595
rect 34253 34561 34287 34595
rect 34287 34561 34296 34595
rect 34244 34552 34296 34561
rect 22376 34484 22428 34536
rect 23480 34484 23532 34536
rect 23848 34527 23900 34536
rect 23848 34493 23857 34527
rect 23857 34493 23891 34527
rect 23891 34493 23900 34527
rect 23848 34484 23900 34493
rect 24952 34527 25004 34536
rect 24952 34493 24961 34527
rect 24961 34493 24995 34527
rect 24995 34493 25004 34527
rect 24952 34484 25004 34493
rect 27620 34527 27672 34536
rect 27620 34493 27629 34527
rect 27629 34493 27663 34527
rect 27663 34493 27672 34527
rect 27620 34484 27672 34493
rect 32220 34484 32272 34536
rect 20168 34416 20220 34468
rect 20260 34416 20312 34468
rect 17040 34348 17092 34400
rect 22192 34348 22244 34400
rect 22560 34391 22612 34400
rect 22560 34357 22569 34391
rect 22569 34357 22603 34391
rect 22603 34357 22612 34391
rect 22560 34348 22612 34357
rect 22744 34391 22796 34400
rect 22744 34357 22753 34391
rect 22753 34357 22787 34391
rect 22787 34357 22796 34391
rect 22744 34348 22796 34357
rect 23204 34459 23256 34468
rect 23204 34425 23213 34459
rect 23213 34425 23247 34459
rect 23247 34425 23256 34459
rect 23204 34416 23256 34425
rect 23388 34416 23440 34468
rect 23664 34416 23716 34468
rect 31392 34416 31444 34468
rect 24676 34348 24728 34400
rect 25228 34348 25280 34400
rect 29184 34391 29236 34400
rect 29184 34357 29193 34391
rect 29193 34357 29227 34391
rect 29227 34357 29236 34391
rect 29184 34348 29236 34357
rect 32404 34348 32456 34400
rect 32956 34484 33008 34536
rect 37740 34552 37792 34604
rect 37832 34416 37884 34468
rect 38016 34527 38068 34536
rect 38016 34493 38025 34527
rect 38025 34493 38059 34527
rect 38059 34493 38068 34527
rect 38016 34484 38068 34493
rect 35348 34348 35400 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 8300 34144 8352 34196
rect 15016 34076 15068 34128
rect 5540 34051 5592 34060
rect 5540 34017 5549 34051
rect 5549 34017 5583 34051
rect 5583 34017 5592 34051
rect 5540 34008 5592 34017
rect 5632 34051 5684 34060
rect 5632 34017 5641 34051
rect 5641 34017 5675 34051
rect 5675 34017 5684 34051
rect 5632 34008 5684 34017
rect 7380 33940 7432 33992
rect 10600 34051 10652 34060
rect 10600 34017 10609 34051
rect 10609 34017 10643 34051
rect 10643 34017 10652 34051
rect 10600 34008 10652 34017
rect 15292 34008 15344 34060
rect 7840 33983 7892 33992
rect 7840 33949 7849 33983
rect 7849 33949 7883 33983
rect 7883 33949 7892 33983
rect 7840 33940 7892 33949
rect 8208 33940 8260 33992
rect 9404 33983 9456 33992
rect 9404 33949 9413 33983
rect 9413 33949 9447 33983
rect 9447 33949 9456 33983
rect 9404 33940 9456 33949
rect 11520 33940 11572 33992
rect 11888 33940 11940 33992
rect 12532 33940 12584 33992
rect 14740 33940 14792 33992
rect 16212 33940 16264 33992
rect 6368 33872 6420 33924
rect 9864 33872 9916 33924
rect 13728 33872 13780 33924
rect 17040 33983 17092 33992
rect 17040 33949 17049 33983
rect 17049 33949 17083 33983
rect 17083 33949 17092 33983
rect 17040 33940 17092 33949
rect 20444 34187 20496 34196
rect 20444 34153 20453 34187
rect 20453 34153 20487 34187
rect 20487 34153 20496 34187
rect 20444 34144 20496 34153
rect 21272 34144 21324 34196
rect 22744 34144 22796 34196
rect 23572 34144 23624 34196
rect 23848 34144 23900 34196
rect 30840 34144 30892 34196
rect 32496 34144 32548 34196
rect 33140 34144 33192 34196
rect 37648 34144 37700 34196
rect 19984 34076 20036 34128
rect 20260 34076 20312 34128
rect 20536 34076 20588 34128
rect 22652 34076 22704 34128
rect 24952 34076 25004 34128
rect 28080 34076 28132 34128
rect 28724 34119 28776 34128
rect 28724 34085 28733 34119
rect 28733 34085 28767 34119
rect 28767 34085 28776 34119
rect 28724 34076 28776 34085
rect 28908 34076 28960 34128
rect 18604 33983 18656 33992
rect 18604 33949 18613 33983
rect 18613 33949 18647 33983
rect 18647 33949 18656 33983
rect 18604 33940 18656 33949
rect 17776 33915 17828 33924
rect 17776 33881 17785 33915
rect 17785 33881 17819 33915
rect 17819 33881 17828 33915
rect 17776 33872 17828 33881
rect 17868 33872 17920 33924
rect 19248 33872 19300 33924
rect 21364 34008 21416 34060
rect 20260 33983 20312 33992
rect 20260 33949 20269 33983
rect 20269 33949 20303 33983
rect 20303 33949 20312 33983
rect 20260 33940 20312 33949
rect 20444 33983 20496 33992
rect 20444 33949 20453 33983
rect 20453 33949 20487 33983
rect 20487 33949 20496 33983
rect 20444 33940 20496 33949
rect 20720 33940 20772 33992
rect 24308 34008 24360 34060
rect 22376 33983 22428 33992
rect 22376 33949 22385 33983
rect 22385 33949 22419 33983
rect 22419 33949 22428 33983
rect 22376 33940 22428 33949
rect 21548 33915 21600 33924
rect 21548 33881 21557 33915
rect 21557 33881 21591 33915
rect 21591 33881 21600 33915
rect 21548 33872 21600 33881
rect 21640 33915 21692 33924
rect 21640 33881 21649 33915
rect 21649 33881 21683 33915
rect 21683 33881 21692 33915
rect 21640 33872 21692 33881
rect 22560 33983 22612 33992
rect 22560 33949 22569 33983
rect 22569 33949 22603 33983
rect 22603 33949 22612 33983
rect 22560 33940 22612 33949
rect 23020 33940 23072 33992
rect 23480 33940 23532 33992
rect 23388 33872 23440 33924
rect 24676 33983 24728 33992
rect 24676 33949 24685 33983
rect 24685 33949 24719 33983
rect 24719 33949 24728 33983
rect 24676 33940 24728 33949
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 25596 33940 25648 33992
rect 26700 34008 26752 34060
rect 25228 33872 25280 33924
rect 25688 33872 25740 33924
rect 26884 33940 26936 33992
rect 29184 33940 29236 33992
rect 29736 33983 29788 33992
rect 29736 33949 29745 33983
rect 29745 33949 29779 33983
rect 29779 33949 29788 33983
rect 29736 33940 29788 33949
rect 29828 33983 29880 33992
rect 29828 33949 29838 33983
rect 29838 33949 29872 33983
rect 29872 33949 29880 33983
rect 35716 34076 35768 34128
rect 29828 33940 29880 33949
rect 30288 33940 30340 33992
rect 31208 33983 31260 33992
rect 31208 33949 31217 33983
rect 31217 33949 31251 33983
rect 31251 33949 31260 33983
rect 31208 33940 31260 33949
rect 33232 34008 33284 34060
rect 36084 34008 36136 34060
rect 38108 34051 38160 34060
rect 38108 34017 38117 34051
rect 38117 34017 38151 34051
rect 38151 34017 38160 34051
rect 38108 34008 38160 34017
rect 31668 33983 31720 33992
rect 31668 33949 31682 33983
rect 31682 33949 31716 33983
rect 31716 33949 31720 33983
rect 31668 33940 31720 33949
rect 37832 33983 37884 33992
rect 37832 33949 37841 33983
rect 37841 33949 37875 33983
rect 37875 33949 37884 33983
rect 37832 33940 37884 33949
rect 26516 33915 26568 33924
rect 26516 33881 26525 33915
rect 26525 33881 26559 33915
rect 26559 33881 26568 33915
rect 26516 33872 26568 33881
rect 27620 33872 27672 33924
rect 30012 33915 30064 33924
rect 30012 33881 30021 33915
rect 30021 33881 30055 33915
rect 30055 33881 30064 33915
rect 30012 33872 30064 33881
rect 30104 33915 30156 33924
rect 30104 33881 30113 33915
rect 30113 33881 30147 33915
rect 30147 33881 30156 33915
rect 30104 33872 30156 33881
rect 6092 33847 6144 33856
rect 6092 33813 6101 33847
rect 6101 33813 6135 33847
rect 6135 33813 6144 33847
rect 6092 33804 6144 33813
rect 8760 33804 8812 33856
rect 14188 33804 14240 33856
rect 15476 33847 15528 33856
rect 15476 33813 15485 33847
rect 15485 33813 15519 33847
rect 15519 33813 15528 33847
rect 15476 33804 15528 33813
rect 17592 33804 17644 33856
rect 18512 33847 18564 33856
rect 18512 33813 18521 33847
rect 18521 33813 18555 33847
rect 18555 33813 18564 33847
rect 18512 33804 18564 33813
rect 19340 33804 19392 33856
rect 30932 33872 30984 33924
rect 31760 33872 31812 33924
rect 32128 33804 32180 33856
rect 32680 33804 32732 33856
rect 35348 33804 35400 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 13636 33643 13688 33652
rect 13636 33609 13645 33643
rect 13645 33609 13679 33643
rect 13679 33609 13688 33643
rect 13636 33600 13688 33609
rect 14740 33643 14792 33652
rect 14740 33609 14749 33643
rect 14749 33609 14783 33643
rect 14783 33609 14792 33643
rect 14740 33600 14792 33609
rect 7104 33575 7156 33584
rect 7104 33541 7113 33575
rect 7113 33541 7147 33575
rect 7147 33541 7156 33575
rect 7104 33532 7156 33541
rect 9404 33532 9456 33584
rect 6552 33464 6604 33516
rect 6000 33439 6052 33448
rect 6000 33405 6009 33439
rect 6009 33405 6043 33439
rect 6043 33405 6052 33439
rect 6000 33396 6052 33405
rect 6828 33396 6880 33448
rect 7380 33328 7432 33380
rect 8392 33328 8444 33380
rect 8760 33507 8812 33516
rect 8760 33473 8769 33507
rect 8769 33473 8803 33507
rect 8803 33473 8812 33507
rect 8760 33464 8812 33473
rect 9680 33507 9732 33516
rect 9680 33473 9689 33507
rect 9689 33473 9723 33507
rect 9723 33473 9732 33507
rect 9680 33464 9732 33473
rect 10600 33507 10652 33516
rect 10600 33473 10609 33507
rect 10609 33473 10643 33507
rect 10643 33473 10652 33507
rect 10600 33464 10652 33473
rect 11520 33464 11572 33516
rect 12256 33464 12308 33516
rect 14096 33507 14148 33516
rect 9312 33396 9364 33448
rect 10048 33396 10100 33448
rect 14096 33473 14105 33507
rect 14105 33473 14139 33507
rect 14139 33473 14148 33507
rect 14096 33464 14148 33473
rect 14556 33507 14608 33516
rect 14556 33473 14565 33507
rect 14565 33473 14599 33507
rect 14599 33473 14608 33507
rect 14556 33464 14608 33473
rect 15200 33464 15252 33516
rect 15384 33507 15436 33516
rect 15384 33473 15393 33507
rect 15393 33473 15427 33507
rect 15427 33473 15436 33507
rect 15384 33464 15436 33473
rect 16120 33600 16172 33652
rect 16764 33600 16816 33652
rect 17868 33600 17920 33652
rect 17960 33600 18012 33652
rect 18972 33600 19024 33652
rect 19432 33600 19484 33652
rect 20352 33600 20404 33652
rect 21640 33600 21692 33652
rect 16212 33532 16264 33584
rect 13544 33396 13596 33448
rect 14464 33439 14516 33448
rect 14464 33405 14473 33439
rect 14473 33405 14507 33439
rect 14507 33405 14516 33439
rect 14464 33396 14516 33405
rect 15660 33439 15712 33448
rect 15660 33405 15669 33439
rect 15669 33405 15703 33439
rect 15703 33405 15712 33439
rect 15660 33396 15712 33405
rect 15568 33328 15620 33380
rect 16948 33464 17000 33516
rect 17776 33464 17828 33516
rect 17960 33396 18012 33448
rect 18696 33464 18748 33516
rect 18880 33464 18932 33516
rect 20536 33532 20588 33584
rect 25688 33600 25740 33652
rect 22376 33532 22428 33584
rect 19432 33507 19484 33516
rect 19432 33473 19441 33507
rect 19441 33473 19475 33507
rect 19475 33473 19484 33507
rect 19432 33464 19484 33473
rect 19616 33507 19668 33516
rect 19616 33473 19625 33507
rect 19625 33473 19659 33507
rect 19659 33473 19668 33507
rect 19616 33464 19668 33473
rect 19708 33507 19760 33516
rect 19708 33473 19717 33507
rect 19717 33473 19751 33507
rect 19751 33473 19760 33507
rect 19708 33464 19760 33473
rect 19984 33464 20036 33516
rect 20168 33507 20220 33516
rect 20168 33473 20177 33507
rect 20177 33473 20211 33507
rect 20211 33473 20220 33507
rect 20168 33464 20220 33473
rect 18420 33396 18472 33448
rect 19892 33396 19944 33448
rect 22836 33464 22888 33516
rect 23388 33464 23440 33516
rect 25596 33532 25648 33584
rect 26608 33600 26660 33652
rect 27436 33600 27488 33652
rect 30104 33600 30156 33652
rect 26516 33532 26568 33584
rect 29460 33532 29512 33584
rect 23204 33439 23256 33448
rect 23204 33405 23213 33439
rect 23213 33405 23247 33439
rect 23247 33405 23256 33439
rect 23204 33396 23256 33405
rect 23572 33396 23624 33448
rect 19616 33328 19668 33380
rect 25136 33396 25188 33448
rect 26148 33507 26200 33516
rect 26148 33473 26157 33507
rect 26157 33473 26191 33507
rect 26191 33473 26200 33507
rect 26148 33464 26200 33473
rect 5632 33260 5684 33312
rect 6552 33260 6604 33312
rect 14188 33303 14240 33312
rect 14188 33269 14197 33303
rect 14197 33269 14231 33303
rect 14231 33269 14240 33303
rect 14188 33260 14240 33269
rect 15476 33303 15528 33312
rect 15476 33269 15485 33303
rect 15485 33269 15519 33303
rect 15519 33269 15528 33303
rect 15476 33260 15528 33269
rect 18328 33260 18380 33312
rect 19984 33260 20036 33312
rect 22192 33260 22244 33312
rect 22652 33260 22704 33312
rect 24860 33260 24912 33312
rect 25780 33328 25832 33380
rect 25228 33260 25280 33312
rect 25872 33260 25924 33312
rect 28632 33507 28684 33516
rect 28632 33473 28641 33507
rect 28641 33473 28675 33507
rect 28675 33473 28684 33507
rect 28632 33464 28684 33473
rect 30932 33532 30984 33584
rect 32404 33600 32456 33652
rect 33416 33575 33468 33584
rect 33416 33541 33425 33575
rect 33425 33541 33459 33575
rect 33459 33541 33468 33575
rect 33416 33532 33468 33541
rect 34428 33600 34480 33652
rect 35992 33600 36044 33652
rect 37832 33600 37884 33652
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 26332 33396 26384 33448
rect 27160 33396 27212 33448
rect 29000 33439 29052 33448
rect 29000 33405 29009 33439
rect 29009 33405 29043 33439
rect 29043 33405 29052 33439
rect 29000 33396 29052 33405
rect 30288 33439 30340 33448
rect 30288 33405 30297 33439
rect 30297 33405 30331 33439
rect 30331 33405 30340 33439
rect 30288 33396 30340 33405
rect 31392 33507 31444 33516
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 31576 33464 31628 33516
rect 33048 33507 33100 33516
rect 33048 33473 33057 33507
rect 33057 33473 33091 33507
rect 33091 33473 33100 33507
rect 33048 33464 33100 33473
rect 33140 33507 33192 33516
rect 33140 33473 33150 33507
rect 33150 33473 33184 33507
rect 33184 33473 33192 33507
rect 33140 33464 33192 33473
rect 28632 33328 28684 33380
rect 32680 33396 32732 33448
rect 34428 33464 34480 33516
rect 37924 33532 37976 33584
rect 34704 33507 34756 33516
rect 34704 33473 34713 33507
rect 34713 33473 34747 33507
rect 34747 33473 34756 33507
rect 34704 33464 34756 33473
rect 34796 33507 34848 33516
rect 34796 33473 34805 33507
rect 34805 33473 34839 33507
rect 34839 33473 34848 33507
rect 34796 33464 34848 33473
rect 34704 33328 34756 33380
rect 35808 33507 35860 33516
rect 35808 33473 35817 33507
rect 35817 33473 35851 33507
rect 35851 33473 35860 33507
rect 35808 33464 35860 33473
rect 35900 33507 35952 33516
rect 35900 33473 35909 33507
rect 35909 33473 35943 33507
rect 35943 33473 35952 33507
rect 35900 33464 35952 33473
rect 35992 33464 36044 33516
rect 36268 33464 36320 33516
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 35716 33396 35768 33448
rect 37740 33396 37792 33448
rect 37924 33439 37976 33448
rect 37924 33405 37933 33439
rect 37933 33405 37967 33439
rect 37967 33405 37976 33439
rect 37924 33396 37976 33405
rect 38016 33439 38068 33448
rect 38016 33405 38025 33439
rect 38025 33405 38059 33439
rect 38059 33405 38068 33439
rect 38016 33396 38068 33405
rect 35808 33260 35860 33312
rect 37096 33260 37148 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4988 33056 5040 33108
rect 8760 33056 8812 33108
rect 13728 33056 13780 33108
rect 14096 33056 14148 33108
rect 15292 33099 15344 33108
rect 15292 33065 15301 33099
rect 15301 33065 15335 33099
rect 15335 33065 15344 33099
rect 15292 33056 15344 33065
rect 15844 33056 15896 33108
rect 9680 32988 9732 33040
rect 10140 32988 10192 33040
rect 18052 33056 18104 33108
rect 18236 33056 18288 33108
rect 4528 32852 4580 32904
rect 6000 32920 6052 32972
rect 10600 32920 10652 32972
rect 5264 32895 5316 32904
rect 5264 32861 5273 32895
rect 5273 32861 5307 32895
rect 5307 32861 5316 32895
rect 5264 32852 5316 32861
rect 6552 32852 6604 32904
rect 7380 32852 7432 32904
rect 6184 32784 6236 32836
rect 7564 32852 7616 32904
rect 7840 32852 7892 32904
rect 8116 32784 8168 32836
rect 8392 32895 8444 32904
rect 8392 32861 8401 32895
rect 8401 32861 8435 32895
rect 8435 32861 8444 32895
rect 8392 32852 8444 32861
rect 9864 32895 9916 32904
rect 9864 32861 9873 32895
rect 9873 32861 9907 32895
rect 9907 32861 9916 32895
rect 9864 32852 9916 32861
rect 10048 32852 10100 32904
rect 11520 32852 11572 32904
rect 12440 32895 12492 32904
rect 12440 32861 12449 32895
rect 12449 32861 12483 32895
rect 12483 32861 12492 32895
rect 12440 32852 12492 32861
rect 12532 32895 12584 32904
rect 12532 32861 12541 32895
rect 12541 32861 12575 32895
rect 12575 32861 12584 32895
rect 12532 32852 12584 32861
rect 13544 32895 13596 32904
rect 13544 32861 13553 32895
rect 13553 32861 13587 32895
rect 13587 32861 13596 32895
rect 13544 32852 13596 32861
rect 14832 32920 14884 32972
rect 14740 32895 14792 32904
rect 14740 32861 14749 32895
rect 14749 32861 14783 32895
rect 14783 32861 14792 32895
rect 15476 32920 15528 32972
rect 17224 32920 17276 32972
rect 19340 32988 19392 33040
rect 14740 32852 14792 32861
rect 15200 32852 15252 32904
rect 9496 32716 9548 32768
rect 10600 32716 10652 32768
rect 12808 32784 12860 32836
rect 14556 32784 14608 32836
rect 15568 32852 15620 32904
rect 17592 32895 17644 32904
rect 17592 32861 17601 32895
rect 17601 32861 17635 32895
rect 17635 32861 17644 32895
rect 17592 32852 17644 32861
rect 18328 32852 18380 32904
rect 18604 32920 18656 32972
rect 22744 33056 22796 33108
rect 25688 33056 25740 33108
rect 30656 33056 30708 33108
rect 31208 33056 31260 33108
rect 31300 33056 31352 33108
rect 20352 32988 20404 33040
rect 20720 32988 20772 33040
rect 25412 33031 25464 33040
rect 25412 32997 25421 33031
rect 25421 32997 25455 33031
rect 25455 32997 25464 33031
rect 25412 32988 25464 32997
rect 20260 32920 20312 32972
rect 20352 32852 20404 32904
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 21640 32920 21692 32972
rect 22836 32920 22888 32972
rect 22560 32852 22612 32904
rect 22928 32895 22980 32904
rect 22928 32861 22937 32895
rect 22937 32861 22971 32895
rect 22971 32861 22980 32895
rect 22928 32852 22980 32861
rect 23388 32920 23440 32972
rect 24952 32920 25004 32972
rect 27620 32988 27672 33040
rect 24584 32852 24636 32904
rect 25228 32895 25280 32904
rect 25228 32861 25237 32895
rect 25237 32861 25271 32895
rect 25271 32861 25280 32895
rect 25228 32852 25280 32861
rect 20812 32827 20864 32836
rect 20812 32793 20821 32827
rect 20821 32793 20855 32827
rect 20855 32793 20864 32827
rect 20812 32784 20864 32793
rect 26240 32895 26292 32904
rect 13636 32716 13688 32768
rect 14280 32716 14332 32768
rect 14372 32716 14424 32768
rect 18420 32716 18472 32768
rect 19340 32716 19392 32768
rect 19432 32716 19484 32768
rect 19892 32716 19944 32768
rect 20260 32759 20312 32768
rect 20260 32725 20269 32759
rect 20269 32725 20303 32759
rect 20303 32725 20312 32759
rect 20260 32716 20312 32725
rect 20904 32716 20956 32768
rect 22744 32759 22796 32768
rect 22744 32725 22753 32759
rect 22753 32725 22787 32759
rect 22787 32725 22796 32759
rect 22744 32716 22796 32725
rect 23572 32716 23624 32768
rect 26240 32861 26249 32895
rect 26249 32861 26283 32895
rect 26283 32861 26292 32895
rect 26240 32852 26292 32861
rect 26700 32895 26752 32904
rect 26700 32861 26709 32895
rect 26709 32861 26743 32895
rect 26743 32861 26752 32895
rect 26700 32852 26752 32861
rect 26056 32784 26108 32836
rect 28172 32895 28224 32904
rect 28172 32861 28181 32895
rect 28181 32861 28215 32895
rect 28215 32861 28224 32895
rect 28172 32852 28224 32861
rect 28724 32895 28776 32904
rect 28724 32861 28733 32895
rect 28733 32861 28767 32895
rect 28767 32861 28776 32895
rect 28724 32852 28776 32861
rect 30288 32988 30340 33040
rect 31944 32988 31996 33040
rect 33048 33056 33100 33108
rect 37832 33056 37884 33108
rect 28816 32784 28868 32836
rect 26148 32716 26200 32768
rect 26608 32716 26660 32768
rect 29920 32852 29972 32904
rect 30288 32852 30340 32904
rect 31300 32895 31352 32904
rect 31300 32861 31345 32895
rect 31345 32861 31352 32895
rect 31300 32852 31352 32861
rect 31484 32895 31536 32904
rect 31484 32861 31493 32895
rect 31493 32861 31527 32895
rect 31527 32861 31536 32895
rect 31484 32852 31536 32861
rect 32588 32920 32640 32972
rect 32220 32895 32272 32904
rect 32220 32861 32229 32895
rect 32229 32861 32263 32895
rect 32263 32861 32272 32895
rect 32220 32852 32272 32861
rect 32312 32895 32364 32904
rect 32312 32861 32321 32895
rect 32321 32861 32355 32895
rect 32355 32861 32364 32895
rect 32312 32852 32364 32861
rect 35440 32852 35492 32904
rect 36360 32920 36412 32972
rect 36084 32895 36136 32904
rect 36084 32861 36093 32895
rect 36093 32861 36127 32895
rect 36127 32861 36136 32895
rect 36084 32852 36136 32861
rect 36268 32852 36320 32904
rect 37096 32895 37148 32904
rect 37096 32861 37130 32895
rect 37130 32861 37148 32895
rect 37096 32852 37148 32861
rect 30012 32827 30064 32836
rect 30012 32793 30021 32827
rect 30021 32793 30055 32827
rect 30055 32793 30064 32827
rect 30012 32784 30064 32793
rect 31116 32827 31168 32836
rect 31116 32793 31125 32827
rect 31125 32793 31159 32827
rect 31159 32793 31168 32827
rect 31116 32784 31168 32793
rect 31668 32784 31720 32836
rect 31760 32716 31812 32768
rect 35808 32716 35860 32768
rect 35900 32716 35952 32768
rect 37924 32716 37976 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 13728 32512 13780 32564
rect 4528 32419 4580 32428
rect 4528 32385 4537 32419
rect 4537 32385 4571 32419
rect 4571 32385 4580 32419
rect 4528 32376 4580 32385
rect 4988 32376 5040 32428
rect 5816 32376 5868 32428
rect 9128 32444 9180 32496
rect 9680 32444 9732 32496
rect 6092 32308 6144 32360
rect 7380 32376 7432 32428
rect 8760 32419 8812 32428
rect 8760 32385 8769 32419
rect 8769 32385 8803 32419
rect 8803 32385 8812 32419
rect 8760 32376 8812 32385
rect 9772 32419 9824 32428
rect 9772 32385 9781 32419
rect 9781 32385 9815 32419
rect 9815 32385 9824 32419
rect 9772 32376 9824 32385
rect 9864 32376 9916 32428
rect 10140 32419 10192 32428
rect 10140 32385 10149 32419
rect 10149 32385 10183 32419
rect 10183 32385 10192 32419
rect 10140 32376 10192 32385
rect 13636 32444 13688 32496
rect 14372 32512 14424 32564
rect 14464 32512 14516 32564
rect 14280 32487 14332 32496
rect 14280 32453 14289 32487
rect 14289 32453 14323 32487
rect 14323 32453 14332 32487
rect 14280 32444 14332 32453
rect 17592 32512 17644 32564
rect 18328 32512 18380 32564
rect 20904 32512 20956 32564
rect 23480 32512 23532 32564
rect 24124 32512 24176 32564
rect 12072 32419 12124 32428
rect 12072 32385 12081 32419
rect 12081 32385 12115 32419
rect 12115 32385 12124 32419
rect 12072 32376 12124 32385
rect 12164 32419 12216 32428
rect 12164 32385 12173 32419
rect 12173 32385 12207 32419
rect 12207 32385 12216 32419
rect 12164 32376 12216 32385
rect 14556 32419 14608 32428
rect 14556 32385 14565 32419
rect 14565 32385 14599 32419
rect 14599 32385 14608 32419
rect 14556 32376 14608 32385
rect 14924 32376 14976 32428
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 16304 32419 16356 32428
rect 16304 32385 16313 32419
rect 16313 32385 16347 32419
rect 16347 32385 16356 32419
rect 16304 32376 16356 32385
rect 20260 32444 20312 32496
rect 21548 32444 21600 32496
rect 25228 32512 25280 32564
rect 9680 32308 9732 32360
rect 11520 32308 11572 32360
rect 15108 32308 15160 32360
rect 17316 32419 17368 32428
rect 17316 32385 17325 32419
rect 17325 32385 17359 32419
rect 17359 32385 17368 32419
rect 17316 32376 17368 32385
rect 20444 32419 20496 32428
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 5632 32240 5684 32292
rect 7012 32240 7064 32292
rect 9312 32240 9364 32292
rect 4896 32172 4948 32224
rect 5724 32172 5776 32224
rect 8024 32172 8076 32224
rect 10600 32172 10652 32224
rect 11888 32283 11940 32292
rect 11888 32249 11897 32283
rect 11897 32249 11931 32283
rect 11931 32249 11940 32283
rect 11888 32240 11940 32249
rect 12992 32240 13044 32292
rect 17132 32308 17184 32360
rect 20720 32308 20772 32360
rect 21916 32308 21968 32360
rect 23480 32419 23532 32428
rect 23480 32385 23489 32419
rect 23489 32385 23523 32419
rect 23523 32385 23532 32419
rect 23480 32376 23532 32385
rect 23848 32419 23900 32428
rect 23848 32385 23857 32419
rect 23857 32385 23891 32419
rect 23891 32385 23900 32419
rect 23848 32376 23900 32385
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 24492 32419 24544 32428
rect 24492 32385 24501 32419
rect 24501 32385 24535 32419
rect 24535 32385 24544 32419
rect 24492 32376 24544 32385
rect 24676 32419 24728 32428
rect 24676 32385 24685 32419
rect 24685 32385 24719 32419
rect 24719 32385 24728 32419
rect 24676 32376 24728 32385
rect 26056 32376 26108 32428
rect 26240 32419 26292 32428
rect 26240 32385 26249 32419
rect 26249 32385 26283 32419
rect 26283 32385 26292 32419
rect 26240 32376 26292 32385
rect 25228 32308 25280 32360
rect 16028 32240 16080 32292
rect 28724 32555 28776 32564
rect 28724 32521 28743 32555
rect 28743 32521 28776 32555
rect 28724 32512 28776 32521
rect 27896 32376 27948 32428
rect 27988 32419 28040 32428
rect 27988 32385 27997 32419
rect 27997 32385 28031 32419
rect 28031 32385 28040 32419
rect 27988 32376 28040 32385
rect 27712 32308 27764 32360
rect 29736 32376 29788 32428
rect 30012 32444 30064 32496
rect 31024 32512 31076 32564
rect 31668 32512 31720 32564
rect 34520 32512 34572 32564
rect 28264 32308 28316 32360
rect 29460 32308 29512 32360
rect 30472 32419 30524 32428
rect 30472 32385 30481 32419
rect 30481 32385 30515 32419
rect 30515 32385 30524 32419
rect 30472 32376 30524 32385
rect 31116 32444 31168 32496
rect 35440 32555 35492 32564
rect 35440 32521 35449 32555
rect 35449 32521 35483 32555
rect 35483 32521 35492 32555
rect 35440 32512 35492 32521
rect 30288 32308 30340 32360
rect 30380 32308 30432 32360
rect 31484 32376 31536 32428
rect 32864 32376 32916 32428
rect 35532 32444 35584 32496
rect 35716 32444 35768 32496
rect 38108 32487 38160 32496
rect 38108 32453 38117 32487
rect 38117 32453 38151 32487
rect 38151 32453 38160 32487
rect 38108 32444 38160 32453
rect 31852 32308 31904 32360
rect 32772 32351 32824 32360
rect 32772 32317 32781 32351
rect 32781 32317 32815 32351
rect 32815 32317 32824 32351
rect 32772 32308 32824 32317
rect 35256 32419 35308 32428
rect 35256 32385 35265 32419
rect 35265 32385 35299 32419
rect 35299 32385 35308 32419
rect 35256 32376 35308 32385
rect 37924 32376 37976 32428
rect 35624 32308 35676 32360
rect 27988 32240 28040 32292
rect 31300 32240 31352 32292
rect 12440 32172 12492 32224
rect 12716 32172 12768 32224
rect 13820 32172 13872 32224
rect 14372 32172 14424 32224
rect 14924 32172 14976 32224
rect 15292 32215 15344 32224
rect 15292 32181 15301 32215
rect 15301 32181 15335 32215
rect 15335 32181 15344 32215
rect 15292 32172 15344 32181
rect 15936 32172 15988 32224
rect 16120 32215 16172 32224
rect 16120 32181 16129 32215
rect 16129 32181 16163 32215
rect 16163 32181 16172 32215
rect 16120 32172 16172 32181
rect 16948 32215 17000 32224
rect 16948 32181 16957 32215
rect 16957 32181 16991 32215
rect 16991 32181 17000 32215
rect 16948 32172 17000 32181
rect 17408 32172 17460 32224
rect 20444 32172 20496 32224
rect 20812 32172 20864 32224
rect 21456 32172 21508 32224
rect 22284 32215 22336 32224
rect 22284 32181 22293 32215
rect 22293 32181 22327 32215
rect 22327 32181 22336 32215
rect 22284 32172 22336 32181
rect 23848 32215 23900 32224
rect 23848 32181 23857 32215
rect 23857 32181 23891 32215
rect 23891 32181 23900 32215
rect 23848 32172 23900 32181
rect 25136 32172 25188 32224
rect 28172 32172 28224 32224
rect 28356 32172 28408 32224
rect 28816 32172 28868 32224
rect 32312 32172 32364 32224
rect 34704 32240 34756 32292
rect 35256 32240 35308 32292
rect 34152 32215 34204 32224
rect 34152 32181 34161 32215
rect 34161 32181 34195 32215
rect 34195 32181 34204 32215
rect 34152 32172 34204 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 5724 31968 5776 32020
rect 3424 31900 3476 31952
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 8024 31968 8076 32020
rect 9680 31968 9732 32020
rect 9772 31968 9824 32020
rect 10324 31968 10376 32020
rect 9588 31900 9640 31952
rect 11980 31900 12032 31952
rect 12716 32011 12768 32020
rect 12716 31977 12725 32011
rect 12725 31977 12759 32011
rect 12759 31977 12768 32011
rect 12716 31968 12768 31977
rect 14740 31968 14792 32020
rect 14832 32011 14884 32020
rect 14832 31977 14841 32011
rect 14841 31977 14875 32011
rect 14875 31977 14884 32011
rect 14832 31968 14884 31977
rect 15200 32011 15252 32020
rect 15200 31977 15209 32011
rect 15209 31977 15243 32011
rect 15243 31977 15252 32011
rect 15200 31968 15252 31977
rect 12992 31943 13044 31952
rect 12992 31909 13001 31943
rect 13001 31909 13035 31943
rect 13035 31909 13044 31943
rect 12992 31900 13044 31909
rect 15568 31900 15620 31952
rect 15844 32011 15896 32020
rect 15844 31977 15853 32011
rect 15853 31977 15887 32011
rect 15887 31977 15896 32011
rect 15844 31968 15896 31977
rect 18052 31968 18104 32020
rect 22100 31968 22152 32020
rect 22560 31968 22612 32020
rect 22836 31968 22888 32020
rect 26700 31968 26752 32020
rect 6092 31832 6144 31884
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 4988 31696 5040 31748
rect 6920 31764 6972 31816
rect 7012 31807 7064 31816
rect 7012 31773 7021 31807
rect 7021 31773 7055 31807
rect 7055 31773 7064 31807
rect 7012 31764 7064 31773
rect 8024 31807 8076 31816
rect 8024 31773 8033 31807
rect 8033 31773 8067 31807
rect 8067 31773 8076 31807
rect 8024 31764 8076 31773
rect 8116 31764 8168 31816
rect 10324 31832 10376 31884
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 9312 31764 9364 31816
rect 9496 31807 9548 31816
rect 9496 31773 9505 31807
rect 9505 31773 9539 31807
rect 9539 31773 9548 31807
rect 9496 31764 9548 31773
rect 9772 31764 9824 31816
rect 11796 31832 11848 31884
rect 10508 31807 10560 31816
rect 10508 31773 10517 31807
rect 10517 31773 10551 31807
rect 10551 31773 10560 31807
rect 10508 31764 10560 31773
rect 11612 31807 11664 31816
rect 11612 31773 11621 31807
rect 11621 31773 11655 31807
rect 11655 31773 11664 31807
rect 11612 31764 11664 31773
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 12072 31832 12124 31884
rect 10140 31696 10192 31748
rect 4068 31671 4120 31680
rect 4068 31637 4077 31671
rect 4077 31637 4111 31671
rect 4111 31637 4120 31671
rect 4068 31628 4120 31637
rect 7012 31628 7064 31680
rect 7748 31671 7800 31680
rect 7748 31637 7757 31671
rect 7757 31637 7791 31671
rect 7791 31637 7800 31671
rect 7748 31628 7800 31637
rect 9588 31671 9640 31680
rect 9588 31637 9597 31671
rect 9597 31637 9631 31671
rect 9631 31637 9640 31671
rect 9588 31628 9640 31637
rect 11704 31628 11756 31680
rect 12348 31764 12400 31816
rect 12808 31807 12860 31816
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 14556 31832 14608 31884
rect 14832 31875 14884 31884
rect 14832 31841 14841 31875
rect 14841 31841 14875 31875
rect 14875 31841 14884 31875
rect 14832 31832 14884 31841
rect 15936 31875 15988 31884
rect 15936 31841 15945 31875
rect 15945 31841 15979 31875
rect 15979 31841 15988 31875
rect 15936 31832 15988 31841
rect 12808 31764 12860 31773
rect 16028 31807 16080 31816
rect 16028 31773 16037 31807
rect 16037 31773 16071 31807
rect 16071 31773 16080 31807
rect 16028 31764 16080 31773
rect 17592 31832 17644 31884
rect 18880 31900 18932 31952
rect 19800 31943 19852 31952
rect 19800 31909 19809 31943
rect 19809 31909 19843 31943
rect 19843 31909 19852 31943
rect 19800 31900 19852 31909
rect 20352 31900 20404 31952
rect 20536 31900 20588 31952
rect 21456 31900 21508 31952
rect 16856 31807 16908 31816
rect 16856 31773 16865 31807
rect 16865 31773 16899 31807
rect 16899 31773 16908 31807
rect 16856 31764 16908 31773
rect 17132 31764 17184 31816
rect 19340 31764 19392 31816
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 21272 31832 21324 31884
rect 22560 31832 22612 31884
rect 23112 31900 23164 31952
rect 25688 31900 25740 31952
rect 26148 31900 26200 31952
rect 29184 31900 29236 31952
rect 24308 31832 24360 31884
rect 21364 31807 21416 31816
rect 21364 31773 21373 31807
rect 21373 31773 21407 31807
rect 21407 31773 21416 31807
rect 21364 31764 21416 31773
rect 22928 31807 22980 31816
rect 22928 31773 22937 31807
rect 22937 31773 22971 31807
rect 22971 31773 22980 31807
rect 22928 31764 22980 31773
rect 13544 31671 13596 31680
rect 13544 31637 13553 31671
rect 13553 31637 13587 31671
rect 13587 31637 13596 31671
rect 13544 31628 13596 31637
rect 15200 31628 15252 31680
rect 15752 31628 15804 31680
rect 16120 31628 16172 31680
rect 18696 31628 18748 31680
rect 20260 31628 20312 31680
rect 21180 31671 21232 31680
rect 21180 31637 21189 31671
rect 21189 31637 21223 31671
rect 21223 31637 21232 31671
rect 21180 31628 21232 31637
rect 23388 31696 23440 31748
rect 23848 31807 23900 31816
rect 23848 31773 23857 31807
rect 23857 31773 23891 31807
rect 23891 31773 23900 31807
rect 23848 31764 23900 31773
rect 24492 31764 24544 31816
rect 25688 31764 25740 31816
rect 25872 31807 25924 31816
rect 25872 31773 25881 31807
rect 25881 31773 25915 31807
rect 25915 31773 25924 31807
rect 25872 31764 25924 31773
rect 25044 31696 25096 31748
rect 27896 31875 27948 31884
rect 27896 31841 27905 31875
rect 27905 31841 27939 31875
rect 27939 31841 27948 31875
rect 27896 31832 27948 31841
rect 28264 31875 28316 31884
rect 28264 31841 28273 31875
rect 28273 31841 28307 31875
rect 28307 31841 28316 31875
rect 28264 31832 28316 31841
rect 27160 31807 27212 31816
rect 27160 31773 27169 31807
rect 27169 31773 27203 31807
rect 27203 31773 27212 31807
rect 27160 31764 27212 31773
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 27988 31807 28040 31816
rect 27988 31773 27997 31807
rect 27997 31773 28031 31807
rect 28031 31773 28040 31807
rect 27988 31764 28040 31773
rect 30288 31968 30340 32020
rect 30288 31832 30340 31884
rect 28632 31764 28684 31816
rect 27068 31696 27120 31748
rect 22468 31628 22520 31680
rect 29368 31696 29420 31748
rect 32036 31807 32088 31816
rect 32036 31773 32045 31807
rect 32045 31773 32079 31807
rect 32079 31773 32088 31807
rect 32036 31764 32088 31773
rect 32864 31968 32916 32020
rect 36544 31968 36596 32020
rect 32956 31807 33008 31816
rect 32956 31773 32965 31807
rect 32965 31773 32999 31807
rect 32999 31773 33008 31807
rect 32956 31764 33008 31773
rect 35256 31807 35308 31816
rect 35256 31773 35265 31807
rect 35265 31773 35299 31807
rect 35299 31773 35308 31807
rect 35256 31764 35308 31773
rect 35440 31764 35492 31816
rect 35992 31832 36044 31884
rect 36360 31875 36412 31884
rect 36360 31841 36369 31875
rect 36369 31841 36403 31875
rect 36403 31841 36412 31875
rect 36360 31832 36412 31841
rect 32220 31696 32272 31748
rect 36268 31764 36320 31816
rect 36912 31696 36964 31748
rect 31116 31628 31168 31680
rect 31576 31628 31628 31680
rect 32404 31628 32456 31680
rect 35900 31671 35952 31680
rect 35900 31637 35909 31671
rect 35909 31637 35943 31671
rect 35943 31637 35952 31671
rect 35900 31628 35952 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5632 31424 5684 31476
rect 6000 31424 6052 31476
rect 6644 31424 6696 31476
rect 7380 31399 7432 31408
rect 7380 31365 7389 31399
rect 7389 31365 7423 31399
rect 7423 31365 7432 31399
rect 7380 31356 7432 31365
rect 8208 31399 8260 31408
rect 8208 31365 8217 31399
rect 8217 31365 8251 31399
rect 8251 31365 8260 31399
rect 8208 31356 8260 31365
rect 9680 31424 9732 31476
rect 11612 31424 11664 31476
rect 4896 31288 4948 31340
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 4988 31288 5040 31297
rect 5448 31288 5500 31340
rect 5816 31331 5868 31340
rect 5816 31297 5825 31331
rect 5825 31297 5859 31331
rect 5859 31297 5868 31331
rect 5816 31288 5868 31297
rect 6092 31288 6144 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 6828 31288 6880 31340
rect 7196 31288 7248 31340
rect 11796 31356 11848 31408
rect 13544 31424 13596 31476
rect 19432 31424 19484 31476
rect 19616 31424 19668 31476
rect 21180 31424 21232 31476
rect 12348 31356 12400 31408
rect 13360 31356 13412 31408
rect 5540 31220 5592 31272
rect 6736 31152 6788 31204
rect 7288 31152 7340 31204
rect 9312 31152 9364 31204
rect 5632 31084 5684 31136
rect 7196 31084 7248 31136
rect 7840 31084 7892 31136
rect 10232 31288 10284 31340
rect 12256 31288 12308 31340
rect 12992 31288 13044 31340
rect 13636 31288 13688 31340
rect 14280 31331 14332 31340
rect 14280 31297 14289 31331
rect 14289 31297 14323 31331
rect 14323 31297 14332 31331
rect 14280 31288 14332 31297
rect 15752 31399 15804 31408
rect 15752 31365 15761 31399
rect 15761 31365 15795 31399
rect 15795 31365 15804 31399
rect 15752 31356 15804 31365
rect 16856 31356 16908 31408
rect 15844 31288 15896 31340
rect 20260 31356 20312 31408
rect 23020 31424 23072 31476
rect 23848 31424 23900 31476
rect 24768 31424 24820 31476
rect 25688 31424 25740 31476
rect 25872 31424 25924 31476
rect 25964 31424 26016 31476
rect 10508 31220 10560 31272
rect 13728 31220 13780 31272
rect 18144 31288 18196 31340
rect 17316 31263 17368 31272
rect 17316 31229 17325 31263
rect 17325 31229 17359 31263
rect 17359 31229 17368 31263
rect 17316 31220 17368 31229
rect 17500 31220 17552 31272
rect 17776 31220 17828 31272
rect 18512 31331 18564 31340
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 18696 31331 18748 31340
rect 18696 31297 18705 31331
rect 18705 31297 18739 31331
rect 18739 31297 18748 31331
rect 18696 31288 18748 31297
rect 19156 31288 19208 31340
rect 20168 31288 20220 31340
rect 21272 31331 21324 31340
rect 21272 31297 21281 31331
rect 21281 31297 21315 31331
rect 21315 31297 21324 31331
rect 21272 31288 21324 31297
rect 22284 31288 22336 31340
rect 22376 31288 22428 31340
rect 23388 31331 23440 31340
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 24492 31288 24544 31340
rect 24860 31331 24912 31340
rect 24860 31297 24869 31331
rect 24869 31297 24903 31331
rect 24903 31297 24912 31331
rect 24860 31288 24912 31297
rect 25688 31288 25740 31340
rect 28264 31424 28316 31476
rect 32220 31424 32272 31476
rect 32956 31424 33008 31476
rect 35256 31424 35308 31476
rect 36544 31467 36596 31476
rect 36544 31433 36553 31467
rect 36553 31433 36587 31467
rect 36587 31433 36596 31467
rect 36544 31424 36596 31433
rect 36912 31467 36964 31476
rect 36912 31433 36921 31467
rect 36921 31433 36955 31467
rect 36955 31433 36964 31467
rect 36912 31424 36964 31433
rect 16672 31152 16724 31204
rect 20260 31220 20312 31272
rect 20812 31220 20864 31272
rect 23480 31263 23532 31272
rect 23480 31229 23489 31263
rect 23489 31229 23523 31263
rect 23523 31229 23532 31263
rect 23480 31220 23532 31229
rect 11796 31084 11848 31136
rect 14188 31084 14240 31136
rect 15292 31084 15344 31136
rect 16212 31084 16264 31136
rect 17776 31084 17828 31136
rect 20352 31152 20404 31204
rect 23388 31152 23440 31204
rect 23756 31220 23808 31272
rect 23940 31220 23992 31272
rect 24400 31220 24452 31272
rect 26240 31331 26292 31340
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 26332 31288 26384 31340
rect 26976 31288 27028 31340
rect 27252 31331 27304 31340
rect 27252 31297 27261 31331
rect 27261 31297 27295 31331
rect 27295 31297 27304 31331
rect 27252 31288 27304 31297
rect 27988 31288 28040 31340
rect 28632 31331 28684 31340
rect 28632 31297 28641 31331
rect 28641 31297 28675 31331
rect 28675 31297 28684 31331
rect 28632 31288 28684 31297
rect 29184 31331 29236 31340
rect 29184 31297 29193 31331
rect 29193 31297 29227 31331
rect 29227 31297 29236 31331
rect 29184 31288 29236 31297
rect 30932 31399 30984 31408
rect 30932 31365 30941 31399
rect 30941 31365 30975 31399
rect 30975 31365 30984 31399
rect 30932 31356 30984 31365
rect 31208 31356 31260 31408
rect 32312 31399 32364 31408
rect 32312 31365 32321 31399
rect 32321 31365 32355 31399
rect 32355 31365 32364 31399
rect 32312 31356 32364 31365
rect 38108 31399 38160 31408
rect 38108 31365 38117 31399
rect 38117 31365 38151 31399
rect 38151 31365 38160 31399
rect 38108 31356 38160 31365
rect 30656 31331 30708 31340
rect 30656 31297 30665 31331
rect 30665 31297 30699 31331
rect 30699 31297 30708 31331
rect 30656 31288 30708 31297
rect 30748 31331 30800 31340
rect 30748 31297 30758 31331
rect 30758 31297 30792 31331
rect 30792 31297 30800 31331
rect 30748 31288 30800 31297
rect 29000 31220 29052 31272
rect 31116 31331 31168 31340
rect 31116 31297 31130 31331
rect 31130 31297 31164 31331
rect 31164 31297 31168 31331
rect 31116 31288 31168 31297
rect 34336 31331 34388 31340
rect 34336 31297 34345 31331
rect 34345 31297 34379 31331
rect 34379 31297 34388 31331
rect 34336 31288 34388 31297
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 34152 31220 34204 31272
rect 31300 31152 31352 31204
rect 34704 31331 34756 31340
rect 34704 31297 34713 31331
rect 34713 31297 34747 31331
rect 34747 31297 34756 31331
rect 34704 31288 34756 31297
rect 35348 31288 35400 31340
rect 35900 31288 35952 31340
rect 38016 31220 38068 31272
rect 22560 31084 22612 31136
rect 22744 31084 22796 31136
rect 25228 31084 25280 31136
rect 25780 31127 25832 31136
rect 25780 31093 25789 31127
rect 25789 31093 25823 31127
rect 25823 31093 25832 31127
rect 25780 31084 25832 31093
rect 27804 31084 27856 31136
rect 32036 31084 32088 31136
rect 34152 31084 34204 31136
rect 35992 31084 36044 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 5264 30880 5316 30932
rect 6736 30923 6788 30932
rect 6736 30889 6745 30923
rect 6745 30889 6779 30923
rect 6779 30889 6788 30923
rect 6736 30880 6788 30889
rect 7012 30923 7064 30932
rect 7012 30889 7021 30923
rect 7021 30889 7055 30923
rect 7055 30889 7064 30923
rect 7012 30880 7064 30889
rect 11888 30880 11940 30932
rect 12164 30880 12216 30932
rect 14556 30923 14608 30932
rect 14556 30889 14565 30923
rect 14565 30889 14599 30923
rect 14599 30889 14608 30923
rect 14556 30880 14608 30889
rect 14648 30880 14700 30932
rect 19524 30880 19576 30932
rect 19984 30880 20036 30932
rect 20444 30923 20496 30932
rect 20444 30889 20453 30923
rect 20453 30889 20487 30923
rect 20487 30889 20496 30923
rect 20444 30880 20496 30889
rect 20812 30880 20864 30932
rect 22100 30880 22152 30932
rect 23296 30880 23348 30932
rect 25412 30880 25464 30932
rect 25872 30880 25924 30932
rect 26332 30923 26384 30932
rect 26332 30889 26341 30923
rect 26341 30889 26375 30923
rect 26375 30889 26384 30923
rect 26332 30880 26384 30889
rect 29736 30880 29788 30932
rect 4804 30812 4856 30864
rect 5816 30812 5868 30864
rect 6460 30744 6512 30796
rect 6552 30744 6604 30796
rect 7840 30855 7892 30864
rect 7840 30821 7849 30855
rect 7849 30821 7883 30855
rect 7883 30821 7892 30855
rect 7840 30812 7892 30821
rect 8116 30812 8168 30864
rect 9312 30812 9364 30864
rect 9588 30812 9640 30864
rect 9680 30744 9732 30796
rect 11612 30744 11664 30796
rect 13728 30787 13780 30796
rect 13728 30753 13737 30787
rect 13737 30753 13771 30787
rect 13771 30753 13780 30787
rect 13728 30744 13780 30753
rect 15476 30744 15528 30796
rect 15752 30812 15804 30864
rect 5816 30676 5868 30728
rect 5264 30651 5316 30660
rect 5264 30617 5273 30651
rect 5273 30617 5307 30651
rect 5307 30617 5316 30651
rect 5264 30608 5316 30617
rect 5908 30651 5960 30660
rect 5908 30617 5917 30651
rect 5917 30617 5951 30651
rect 5951 30617 5960 30651
rect 5908 30608 5960 30617
rect 6552 30651 6604 30660
rect 6552 30617 6561 30651
rect 6561 30617 6595 30651
rect 6595 30617 6604 30651
rect 6552 30608 6604 30617
rect 7288 30676 7340 30728
rect 7748 30719 7800 30728
rect 7748 30685 7757 30719
rect 7757 30685 7791 30719
rect 7791 30685 7800 30719
rect 7748 30676 7800 30685
rect 7840 30676 7892 30728
rect 9404 30719 9456 30728
rect 9404 30685 9413 30719
rect 9413 30685 9447 30719
rect 9447 30685 9456 30719
rect 9404 30676 9456 30685
rect 11060 30676 11112 30728
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 11980 30719 12032 30728
rect 11980 30685 11989 30719
rect 11989 30685 12023 30719
rect 12023 30685 12032 30719
rect 11980 30676 12032 30685
rect 7012 30608 7064 30660
rect 11612 30608 11664 30660
rect 12256 30676 12308 30728
rect 12992 30676 13044 30728
rect 14188 30676 14240 30728
rect 15108 30676 15160 30728
rect 4988 30540 5040 30592
rect 5632 30540 5684 30592
rect 7748 30540 7800 30592
rect 11980 30540 12032 30592
rect 13820 30540 13872 30592
rect 14740 30540 14792 30592
rect 15200 30583 15252 30592
rect 15200 30549 15209 30583
rect 15209 30549 15243 30583
rect 15243 30549 15252 30583
rect 15200 30540 15252 30549
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 15844 30676 15896 30728
rect 16304 30676 16356 30728
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 17684 30676 17736 30728
rect 17040 30608 17092 30660
rect 17868 30719 17920 30728
rect 17868 30685 17877 30719
rect 17877 30685 17911 30719
rect 17911 30685 17920 30719
rect 17868 30676 17920 30685
rect 18052 30651 18104 30660
rect 18052 30617 18061 30651
rect 18061 30617 18095 30651
rect 18095 30617 18104 30651
rect 18052 30608 18104 30617
rect 18604 30608 18656 30660
rect 19340 30744 19392 30796
rect 19616 30719 19668 30728
rect 19616 30685 19625 30719
rect 19625 30685 19659 30719
rect 19659 30685 19668 30719
rect 19616 30676 19668 30685
rect 25780 30812 25832 30864
rect 26240 30812 26292 30864
rect 27528 30812 27580 30864
rect 36728 30880 36780 30932
rect 32036 30812 32088 30864
rect 20444 30744 20496 30796
rect 20536 30676 20588 30728
rect 21088 30719 21140 30728
rect 21088 30685 21097 30719
rect 21097 30685 21131 30719
rect 21131 30685 21140 30719
rect 21088 30676 21140 30685
rect 21272 30676 21324 30728
rect 22744 30744 22796 30796
rect 25136 30744 25188 30796
rect 22652 30719 22704 30728
rect 22652 30685 22661 30719
rect 22661 30685 22695 30719
rect 22695 30685 22704 30719
rect 22652 30676 22704 30685
rect 23388 30676 23440 30728
rect 23572 30676 23624 30728
rect 23848 30719 23900 30728
rect 23848 30685 23857 30719
rect 23857 30685 23891 30719
rect 23891 30685 23900 30719
rect 23848 30676 23900 30685
rect 24216 30676 24268 30728
rect 16304 30540 16356 30592
rect 17868 30540 17920 30592
rect 18144 30540 18196 30592
rect 19432 30540 19484 30592
rect 22744 30608 22796 30660
rect 25504 30676 25556 30728
rect 25780 30676 25832 30728
rect 31116 30744 31168 30796
rect 33876 30744 33928 30796
rect 26056 30719 26108 30728
rect 26056 30685 26065 30719
rect 26065 30685 26099 30719
rect 26099 30685 26108 30719
rect 26056 30676 26108 30685
rect 27068 30676 27120 30728
rect 27528 30676 27580 30728
rect 28172 30676 28224 30728
rect 28264 30719 28316 30728
rect 28264 30685 28273 30719
rect 28273 30685 28307 30719
rect 28307 30685 28316 30719
rect 28264 30676 28316 30685
rect 29184 30676 29236 30728
rect 29828 30719 29880 30728
rect 29828 30685 29837 30719
rect 29837 30685 29871 30719
rect 29871 30685 29880 30719
rect 29828 30676 29880 30685
rect 26700 30608 26752 30660
rect 27252 30608 27304 30660
rect 30748 30719 30800 30728
rect 30748 30685 30757 30719
rect 30757 30685 30791 30719
rect 30791 30685 30800 30719
rect 30748 30676 30800 30685
rect 20904 30540 20956 30592
rect 22836 30583 22888 30592
rect 22836 30549 22845 30583
rect 22845 30549 22879 30583
rect 22879 30549 22888 30583
rect 22836 30540 22888 30549
rect 30472 30608 30524 30660
rect 30932 30676 30984 30728
rect 27528 30540 27580 30592
rect 28908 30540 28960 30592
rect 31484 30676 31536 30728
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 37832 30719 37884 30728
rect 37832 30685 37841 30719
rect 37841 30685 37875 30719
rect 37875 30685 37884 30719
rect 37832 30676 37884 30685
rect 31116 30651 31168 30660
rect 31116 30617 31125 30651
rect 31125 30617 31159 30651
rect 31159 30617 31168 30651
rect 31116 30608 31168 30617
rect 32680 30608 32732 30660
rect 39028 30608 39080 30660
rect 31300 30540 31352 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5908 30336 5960 30388
rect 7380 30268 7432 30320
rect 8392 30268 8444 30320
rect 2780 30243 2832 30252
rect 2780 30209 2789 30243
rect 2789 30209 2823 30243
rect 2823 30209 2832 30243
rect 2780 30200 2832 30209
rect 3976 30200 4028 30252
rect 4804 30243 4856 30252
rect 4804 30209 4813 30243
rect 4813 30209 4847 30243
rect 4847 30209 4856 30243
rect 4804 30200 4856 30209
rect 5080 30200 5132 30252
rect 5540 30243 5592 30252
rect 5540 30209 5549 30243
rect 5549 30209 5583 30243
rect 5583 30209 5592 30243
rect 5540 30200 5592 30209
rect 5816 30243 5868 30252
rect 5816 30209 5825 30243
rect 5825 30209 5859 30243
rect 5859 30209 5868 30243
rect 5816 30200 5868 30209
rect 6460 30200 6512 30252
rect 4896 30132 4948 30184
rect 7104 30132 7156 30184
rect 7472 30200 7524 30252
rect 9404 30268 9456 30320
rect 7656 30132 7708 30184
rect 8760 30243 8812 30252
rect 8760 30209 8769 30243
rect 8769 30209 8803 30243
rect 8803 30209 8812 30243
rect 8760 30200 8812 30209
rect 9036 30200 9088 30252
rect 9680 30243 9732 30252
rect 9680 30209 9689 30243
rect 9689 30209 9723 30243
rect 9723 30209 9732 30243
rect 9680 30200 9732 30209
rect 14372 30336 14424 30388
rect 15568 30336 15620 30388
rect 18328 30336 18380 30388
rect 20352 30336 20404 30388
rect 24216 30336 24268 30388
rect 9864 30311 9916 30320
rect 9864 30277 9873 30311
rect 9873 30277 9907 30311
rect 9907 30277 9916 30311
rect 9864 30268 9916 30277
rect 10324 30311 10376 30320
rect 10324 30277 10333 30311
rect 10333 30277 10367 30311
rect 10367 30277 10376 30311
rect 10324 30268 10376 30277
rect 10692 30268 10744 30320
rect 15752 30268 15804 30320
rect 16488 30268 16540 30320
rect 18144 30268 18196 30320
rect 9312 30132 9364 30184
rect 11796 30243 11848 30252
rect 11796 30209 11805 30243
rect 11805 30209 11839 30243
rect 11839 30209 11848 30243
rect 11796 30200 11848 30209
rect 4620 29996 4672 30048
rect 4804 30039 4856 30048
rect 4804 30005 4813 30039
rect 4813 30005 4847 30039
rect 4847 30005 4856 30039
rect 4804 29996 4856 30005
rect 6000 30039 6052 30048
rect 6000 30005 6009 30039
rect 6009 30005 6043 30039
rect 6043 30005 6052 30039
rect 6000 29996 6052 30005
rect 6092 29996 6144 30048
rect 9036 29996 9088 30048
rect 10508 30064 10560 30116
rect 11612 30064 11664 30116
rect 11888 30064 11940 30116
rect 12992 30132 13044 30184
rect 15384 30243 15436 30252
rect 15384 30209 15393 30243
rect 15393 30209 15427 30243
rect 15427 30209 15436 30243
rect 15384 30200 15436 30209
rect 16672 30200 16724 30252
rect 17776 30243 17828 30252
rect 17776 30209 17785 30243
rect 17785 30209 17819 30243
rect 17819 30209 17828 30243
rect 17776 30200 17828 30209
rect 17868 30243 17920 30252
rect 17868 30209 17877 30243
rect 17877 30209 17911 30243
rect 17911 30209 17920 30243
rect 17868 30200 17920 30209
rect 18328 30243 18380 30252
rect 18328 30209 18337 30243
rect 18337 30209 18371 30243
rect 18371 30209 18380 30243
rect 18328 30200 18380 30209
rect 20260 30200 20312 30252
rect 20352 30243 20404 30252
rect 20352 30209 20361 30243
rect 20361 30209 20395 30243
rect 20395 30209 20404 30243
rect 20352 30200 20404 30209
rect 23204 30200 23256 30252
rect 23572 30200 23624 30252
rect 14740 30132 14792 30184
rect 18604 30132 18656 30184
rect 21456 30132 21508 30184
rect 23296 30132 23348 30184
rect 15292 30064 15344 30116
rect 15660 30064 15712 30116
rect 17408 30064 17460 30116
rect 17776 30064 17828 30116
rect 12532 29996 12584 30048
rect 14464 30039 14516 30048
rect 14464 30005 14473 30039
rect 14473 30005 14507 30039
rect 14507 30005 14516 30039
rect 14464 29996 14516 30005
rect 14556 29996 14608 30048
rect 17592 29996 17644 30048
rect 18512 30039 18564 30048
rect 18512 30005 18521 30039
rect 18521 30005 18555 30039
rect 18555 30005 18564 30039
rect 18512 29996 18564 30005
rect 20720 29996 20772 30048
rect 22652 29996 22704 30048
rect 22928 30107 22980 30116
rect 22928 30073 22937 30107
rect 22937 30073 22971 30107
rect 22971 30073 22980 30107
rect 22928 30064 22980 30073
rect 23112 29996 23164 30048
rect 24308 30200 24360 30252
rect 24492 30268 24544 30320
rect 25964 30336 26016 30388
rect 27252 30336 27304 30388
rect 27712 30336 27764 30388
rect 29368 30336 29420 30388
rect 30656 30336 30708 30388
rect 25504 30268 25556 30320
rect 27436 30268 27488 30320
rect 25412 30243 25464 30252
rect 25412 30209 25421 30243
rect 25421 30209 25455 30243
rect 25455 30209 25464 30243
rect 25412 30200 25464 30209
rect 25596 30243 25648 30252
rect 25596 30209 25605 30243
rect 25605 30209 25639 30243
rect 25639 30209 25648 30243
rect 25596 30200 25648 30209
rect 25964 30243 26016 30252
rect 25964 30209 25973 30243
rect 25973 30209 26007 30243
rect 26007 30209 26016 30243
rect 25964 30200 26016 30209
rect 27620 30243 27672 30252
rect 27620 30209 27629 30243
rect 27629 30209 27663 30243
rect 27663 30209 27672 30243
rect 27620 30200 27672 30209
rect 29092 30268 29144 30320
rect 30012 30311 30064 30320
rect 30012 30277 30021 30311
rect 30021 30277 30055 30311
rect 30055 30277 30064 30311
rect 30012 30268 30064 30277
rect 30472 30268 30524 30320
rect 33876 30311 33928 30320
rect 33876 30277 33910 30311
rect 33910 30277 33928 30311
rect 33876 30268 33928 30277
rect 35900 30336 35952 30388
rect 29736 30243 29788 30252
rect 29736 30209 29745 30243
rect 29745 30209 29779 30243
rect 29779 30209 29788 30243
rect 29736 30200 29788 30209
rect 24768 30132 24820 30184
rect 25320 30132 25372 30184
rect 26148 30132 26200 30184
rect 27436 30132 27488 30184
rect 29092 30132 29144 30184
rect 30104 30243 30156 30252
rect 30104 30209 30113 30243
rect 30113 30209 30147 30243
rect 30147 30209 30156 30243
rect 30104 30200 30156 30209
rect 30288 30200 30340 30252
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 32680 30243 32732 30252
rect 32680 30209 32689 30243
rect 32689 30209 32723 30243
rect 32723 30209 32732 30243
rect 32680 30200 32732 30209
rect 33324 30132 33376 30184
rect 35440 30200 35492 30252
rect 38200 30268 38252 30320
rect 35992 30243 36044 30252
rect 35992 30209 36001 30243
rect 36001 30209 36035 30243
rect 36035 30209 36044 30243
rect 35992 30200 36044 30209
rect 36268 30200 36320 30252
rect 25412 30064 25464 30116
rect 29000 30039 29052 30048
rect 29000 30005 29009 30039
rect 29009 30005 29043 30039
rect 29043 30005 29052 30039
rect 29000 29996 29052 30005
rect 30104 30064 30156 30116
rect 33416 30064 33468 30116
rect 35992 30064 36044 30116
rect 37832 30064 37884 30116
rect 38016 30175 38068 30184
rect 38016 30141 38025 30175
rect 38025 30141 38059 30175
rect 38059 30141 38068 30175
rect 38016 30132 38068 30141
rect 31024 29996 31076 30048
rect 33140 29996 33192 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3976 29835 4028 29844
rect 3976 29801 3985 29835
rect 3985 29801 4019 29835
rect 4019 29801 4028 29835
rect 3976 29792 4028 29801
rect 3424 29699 3476 29708
rect 3424 29665 3433 29699
rect 3433 29665 3467 29699
rect 3467 29665 3476 29699
rect 3424 29656 3476 29665
rect 10140 29792 10192 29844
rect 11152 29792 11204 29844
rect 12072 29835 12124 29844
rect 12072 29801 12081 29835
rect 12081 29801 12115 29835
rect 12115 29801 12124 29835
rect 12072 29792 12124 29801
rect 17224 29835 17276 29844
rect 17224 29801 17233 29835
rect 17233 29801 17267 29835
rect 17267 29801 17276 29835
rect 17224 29792 17276 29801
rect 6000 29724 6052 29776
rect 13820 29724 13872 29776
rect 16212 29724 16264 29776
rect 19984 29792 20036 29844
rect 17592 29724 17644 29776
rect 3148 29631 3200 29640
rect 3148 29597 3157 29631
rect 3157 29597 3191 29631
rect 3191 29597 3200 29631
rect 3148 29588 3200 29597
rect 3332 29631 3384 29640
rect 3332 29597 3341 29631
rect 3341 29597 3375 29631
rect 3375 29597 3384 29631
rect 3332 29588 3384 29597
rect 13268 29656 13320 29708
rect 15476 29656 15528 29708
rect 18512 29656 18564 29708
rect 19432 29656 19484 29708
rect 4620 29452 4672 29504
rect 5632 29588 5684 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 7380 29588 7432 29640
rect 7564 29631 7616 29640
rect 7564 29597 7573 29631
rect 7573 29597 7607 29631
rect 7607 29597 7616 29631
rect 7564 29588 7616 29597
rect 7656 29588 7708 29640
rect 9404 29588 9456 29640
rect 14096 29588 14148 29640
rect 16488 29631 16540 29640
rect 16488 29597 16497 29631
rect 16497 29597 16531 29631
rect 16531 29597 16540 29631
rect 16488 29588 16540 29597
rect 16764 29588 16816 29640
rect 17408 29631 17460 29640
rect 17408 29597 17417 29631
rect 17417 29597 17451 29631
rect 17451 29597 17460 29631
rect 17408 29588 17460 29597
rect 17868 29588 17920 29640
rect 20260 29588 20312 29640
rect 21732 29792 21784 29844
rect 22468 29792 22520 29844
rect 22744 29724 22796 29776
rect 23020 29792 23072 29844
rect 23296 29792 23348 29844
rect 23388 29835 23440 29844
rect 23388 29801 23397 29835
rect 23397 29801 23431 29835
rect 23431 29801 23440 29835
rect 23388 29792 23440 29801
rect 25780 29792 25832 29844
rect 29000 29792 29052 29844
rect 30748 29792 30800 29844
rect 31024 29792 31076 29844
rect 31668 29792 31720 29844
rect 32496 29792 32548 29844
rect 21640 29699 21692 29708
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 24032 29724 24084 29776
rect 26424 29724 26476 29776
rect 28908 29724 28960 29776
rect 34612 29792 34664 29844
rect 35440 29835 35492 29844
rect 35440 29801 35449 29835
rect 35449 29801 35483 29835
rect 35483 29801 35492 29835
rect 35440 29792 35492 29801
rect 36268 29835 36320 29844
rect 36268 29801 36277 29835
rect 36277 29801 36311 29835
rect 36311 29801 36320 29835
rect 36268 29792 36320 29801
rect 38200 29835 38252 29844
rect 38200 29801 38209 29835
rect 38209 29801 38243 29835
rect 38243 29801 38252 29835
rect 38200 29792 38252 29801
rect 5080 29452 5132 29504
rect 5632 29452 5684 29504
rect 8208 29520 8260 29572
rect 10140 29520 10192 29572
rect 11796 29520 11848 29572
rect 11888 29563 11940 29572
rect 11888 29529 11897 29563
rect 11897 29529 11931 29563
rect 11931 29529 11940 29563
rect 11888 29520 11940 29529
rect 12348 29520 12400 29572
rect 14188 29520 14240 29572
rect 14464 29520 14516 29572
rect 16120 29520 16172 29572
rect 17684 29563 17736 29572
rect 17684 29529 17693 29563
rect 17693 29529 17727 29563
rect 17727 29529 17736 29563
rect 17684 29520 17736 29529
rect 7564 29495 7616 29504
rect 7564 29461 7573 29495
rect 7573 29461 7607 29495
rect 7607 29461 7616 29495
rect 7564 29452 7616 29461
rect 11704 29452 11756 29504
rect 14096 29452 14148 29504
rect 16580 29495 16632 29504
rect 16580 29461 16589 29495
rect 16589 29461 16623 29495
rect 16623 29461 16632 29495
rect 16580 29452 16632 29461
rect 20352 29452 20404 29504
rect 21732 29631 21784 29640
rect 21732 29597 21741 29631
rect 21741 29597 21775 29631
rect 21775 29597 21784 29631
rect 21732 29588 21784 29597
rect 21916 29588 21968 29640
rect 22192 29563 22244 29572
rect 22192 29529 22201 29563
rect 22201 29529 22235 29563
rect 22235 29529 22244 29563
rect 22192 29520 22244 29529
rect 22560 29588 22612 29640
rect 23112 29588 23164 29640
rect 23296 29631 23348 29640
rect 23296 29597 23305 29631
rect 23305 29597 23339 29631
rect 23339 29597 23348 29631
rect 23296 29588 23348 29597
rect 23388 29588 23440 29640
rect 22652 29452 22704 29504
rect 23756 29520 23808 29572
rect 26240 29588 26292 29640
rect 27436 29631 27488 29640
rect 27436 29597 27445 29631
rect 27445 29597 27479 29631
rect 27479 29597 27488 29631
rect 27436 29588 27488 29597
rect 28816 29699 28868 29708
rect 28816 29665 28825 29699
rect 28825 29665 28859 29699
rect 28859 29665 28868 29699
rect 28816 29656 28868 29665
rect 30748 29656 30800 29708
rect 25136 29452 25188 29504
rect 27252 29520 27304 29572
rect 29276 29588 29328 29640
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 29920 29631 29972 29640
rect 29920 29597 29927 29631
rect 29927 29597 29972 29631
rect 29920 29588 29972 29597
rect 30012 29631 30064 29640
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 30012 29588 30064 29597
rect 30288 29588 30340 29640
rect 30380 29588 30432 29640
rect 36360 29656 36412 29708
rect 27068 29495 27120 29504
rect 27068 29461 27077 29495
rect 27077 29461 27111 29495
rect 27111 29461 27120 29495
rect 29644 29520 29696 29572
rect 30104 29563 30156 29572
rect 30104 29529 30113 29563
rect 30113 29529 30147 29563
rect 30147 29529 30156 29563
rect 30104 29520 30156 29529
rect 27068 29452 27120 29461
rect 28448 29452 28500 29504
rect 31484 29631 31536 29640
rect 31484 29597 31498 29631
rect 31498 29597 31532 29631
rect 31532 29597 31536 29631
rect 31484 29588 31536 29597
rect 32404 29631 32456 29640
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 33416 29588 33468 29640
rect 35440 29588 35492 29640
rect 36084 29631 36136 29640
rect 36084 29597 36093 29631
rect 36093 29597 36127 29631
rect 36127 29597 36136 29631
rect 36084 29588 36136 29597
rect 37464 29588 37516 29640
rect 31300 29563 31352 29572
rect 31300 29529 31309 29563
rect 31309 29529 31343 29563
rect 31343 29529 31352 29563
rect 31300 29520 31352 29529
rect 31484 29452 31536 29504
rect 32496 29520 32548 29572
rect 33140 29563 33192 29572
rect 33140 29529 33174 29563
rect 33174 29529 33192 29563
rect 33140 29520 33192 29529
rect 33324 29520 33376 29572
rect 34520 29520 34572 29572
rect 35072 29563 35124 29572
rect 35072 29529 35081 29563
rect 35081 29529 35115 29563
rect 35115 29529 35124 29563
rect 35072 29520 35124 29529
rect 35164 29563 35216 29572
rect 35164 29529 35173 29563
rect 35173 29529 35207 29563
rect 35207 29529 35216 29563
rect 35164 29520 35216 29529
rect 32312 29495 32364 29504
rect 32312 29461 32321 29495
rect 32321 29461 32355 29495
rect 32355 29461 32364 29495
rect 32312 29452 32364 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5816 29248 5868 29300
rect 3332 29180 3384 29232
rect 3976 29180 4028 29232
rect 4804 29180 4856 29232
rect 3148 29112 3200 29164
rect 4896 29112 4948 29164
rect 5264 29155 5316 29164
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 6000 29112 6052 29164
rect 6828 29180 6880 29232
rect 6920 29223 6972 29232
rect 6920 29189 6929 29223
rect 6929 29189 6963 29223
rect 6963 29189 6972 29223
rect 6920 29180 6972 29189
rect 7012 29180 7064 29232
rect 7472 29112 7524 29164
rect 5172 29044 5224 29096
rect 5448 29087 5500 29096
rect 5448 29053 5457 29087
rect 5457 29053 5491 29087
rect 5491 29053 5500 29087
rect 5448 29044 5500 29053
rect 8760 29112 8812 29164
rect 11152 29291 11204 29300
rect 11152 29257 11161 29291
rect 11161 29257 11195 29291
rect 11195 29257 11204 29291
rect 11152 29248 11204 29257
rect 11980 29248 12032 29300
rect 11704 29223 11756 29232
rect 11704 29189 11713 29223
rect 11713 29189 11747 29223
rect 11747 29189 11756 29223
rect 11704 29180 11756 29189
rect 9496 29112 9548 29164
rect 9956 29155 10008 29164
rect 9956 29121 9965 29155
rect 9965 29121 9999 29155
rect 9999 29121 10008 29155
rect 9956 29112 10008 29121
rect 10048 29155 10100 29164
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 8208 29044 8260 29096
rect 4620 28976 4672 29028
rect 5080 29019 5132 29028
rect 5080 28985 5089 29019
rect 5089 28985 5123 29019
rect 5123 28985 5132 29019
rect 5080 28976 5132 28985
rect 7748 28976 7800 29028
rect 9588 29044 9640 29096
rect 11152 29155 11204 29164
rect 11152 29121 11161 29155
rect 11161 29121 11195 29155
rect 11195 29121 11204 29155
rect 11152 29112 11204 29121
rect 9680 28976 9732 29028
rect 10508 28976 10560 29028
rect 12440 29112 12492 29164
rect 14832 29248 14884 29300
rect 16212 29248 16264 29300
rect 18420 29248 18472 29300
rect 19340 29248 19392 29300
rect 13820 29180 13872 29232
rect 16580 29180 16632 29232
rect 12992 29112 13044 29164
rect 13268 29155 13320 29164
rect 13268 29121 13277 29155
rect 13277 29121 13311 29155
rect 13311 29121 13320 29155
rect 13268 29112 13320 29121
rect 13912 29112 13964 29164
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 16948 29112 17000 29164
rect 20168 29180 20220 29232
rect 5356 28951 5408 28960
rect 5356 28917 5365 28951
rect 5365 28917 5399 28951
rect 5399 28917 5408 28951
rect 5356 28908 5408 28917
rect 5908 28908 5960 28960
rect 6644 28951 6696 28960
rect 6644 28917 6653 28951
rect 6653 28917 6687 28951
rect 6687 28917 6696 28951
rect 6644 28908 6696 28917
rect 6828 28908 6880 28960
rect 9128 28908 9180 28960
rect 10140 28908 10192 28960
rect 11152 28908 11204 28960
rect 11980 28908 12032 28960
rect 13176 28908 13228 28960
rect 13452 28951 13504 28960
rect 13452 28917 13461 28951
rect 13461 28917 13495 28951
rect 13495 28917 13504 28951
rect 13452 28908 13504 28917
rect 14740 29044 14792 29096
rect 15844 29087 15896 29096
rect 15844 29053 15853 29087
rect 15853 29053 15887 29087
rect 15887 29053 15896 29087
rect 15844 29044 15896 29053
rect 17592 29112 17644 29164
rect 17960 29112 18012 29164
rect 13912 28976 13964 29028
rect 15108 28976 15160 29028
rect 17500 29044 17552 29096
rect 18972 29112 19024 29164
rect 19616 29155 19668 29164
rect 19616 29121 19625 29155
rect 19625 29121 19659 29155
rect 19659 29121 19668 29155
rect 19616 29112 19668 29121
rect 20444 29180 20496 29232
rect 18512 29044 18564 29096
rect 19156 29044 19208 29096
rect 19248 29044 19300 29096
rect 20996 29112 21048 29164
rect 22192 29112 22244 29164
rect 19800 29044 19852 29096
rect 20260 29044 20312 29096
rect 22468 29044 22520 29096
rect 23388 29291 23440 29300
rect 23388 29257 23397 29291
rect 23397 29257 23431 29291
rect 23431 29257 23440 29291
rect 23388 29248 23440 29257
rect 23664 29248 23716 29300
rect 24952 29291 25004 29300
rect 24952 29257 24961 29291
rect 24961 29257 24995 29291
rect 24995 29257 25004 29291
rect 24952 29248 25004 29257
rect 24308 29180 24360 29232
rect 25688 29248 25740 29300
rect 27160 29248 27212 29300
rect 30104 29248 30156 29300
rect 23756 29155 23808 29164
rect 23756 29121 23765 29155
rect 23765 29121 23799 29155
rect 23799 29121 23808 29155
rect 23756 29112 23808 29121
rect 23848 29155 23900 29164
rect 23848 29121 23857 29155
rect 23857 29121 23891 29155
rect 23891 29121 23900 29155
rect 25320 29180 25372 29232
rect 27068 29180 27120 29232
rect 27988 29180 28040 29232
rect 28264 29180 28316 29232
rect 28632 29180 28684 29232
rect 23848 29112 23900 29121
rect 24952 29112 25004 29164
rect 25504 29112 25556 29164
rect 27160 29155 27212 29164
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 27252 29112 27304 29164
rect 23388 29044 23440 29096
rect 25044 29044 25096 29096
rect 18880 28976 18932 29028
rect 19616 28976 19668 29028
rect 20720 28976 20772 29028
rect 21456 28976 21508 29028
rect 22100 28976 22152 29028
rect 23020 28976 23072 29028
rect 24860 28976 24912 29028
rect 25228 29087 25280 29096
rect 25228 29053 25237 29087
rect 25237 29053 25271 29087
rect 25271 29053 25280 29087
rect 25228 29044 25280 29053
rect 25320 29087 25372 29096
rect 25320 29053 25329 29087
rect 25329 29053 25363 29087
rect 25363 29053 25372 29087
rect 25320 29044 25372 29053
rect 25688 29044 25740 29096
rect 26056 29087 26108 29096
rect 26056 29053 26065 29087
rect 26065 29053 26099 29087
rect 26099 29053 26108 29087
rect 26056 29044 26108 29053
rect 26976 29044 27028 29096
rect 28264 29044 28316 29096
rect 29092 29112 29144 29164
rect 29000 29044 29052 29096
rect 30656 29112 30708 29164
rect 30932 29112 30984 29164
rect 31392 29112 31444 29164
rect 31484 29155 31536 29164
rect 31484 29121 31493 29155
rect 31493 29121 31527 29155
rect 31527 29121 31536 29155
rect 31484 29112 31536 29121
rect 32496 29291 32548 29300
rect 32496 29257 32505 29291
rect 32505 29257 32539 29291
rect 32539 29257 32548 29291
rect 32496 29248 32548 29257
rect 32680 29291 32732 29300
rect 32680 29257 32689 29291
rect 32689 29257 32723 29291
rect 32723 29257 32732 29291
rect 32680 29248 32732 29257
rect 32312 29223 32364 29232
rect 32312 29189 32321 29223
rect 32321 29189 32355 29223
rect 32355 29189 32364 29223
rect 32312 29180 32364 29189
rect 33048 29180 33100 29232
rect 35072 29223 35124 29232
rect 35072 29189 35081 29223
rect 35081 29189 35115 29223
rect 35115 29189 35124 29223
rect 35072 29180 35124 29189
rect 35348 29180 35400 29232
rect 38016 29180 38068 29232
rect 26240 28976 26292 29028
rect 28172 29019 28224 29028
rect 28172 28985 28181 29019
rect 28181 28985 28215 29019
rect 28215 28985 28224 29019
rect 28172 28976 28224 28985
rect 29092 28976 29144 29028
rect 35440 29112 35492 29164
rect 36176 29112 36228 29164
rect 37556 29155 37608 29164
rect 37556 29121 37565 29155
rect 37565 29121 37599 29155
rect 37599 29121 37608 29155
rect 37556 29112 37608 29121
rect 39028 29044 39080 29096
rect 21088 28908 21140 28960
rect 25044 28908 25096 28960
rect 25596 28908 25648 28960
rect 28908 28908 28960 28960
rect 31116 28908 31168 28960
rect 32404 28908 32456 28960
rect 35532 28908 35584 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3976 28704 4028 28756
rect 4988 28704 5040 28756
rect 5356 28704 5408 28756
rect 9220 28704 9272 28756
rect 5448 28543 5500 28552
rect 5448 28509 5457 28543
rect 5457 28509 5491 28543
rect 5491 28509 5500 28543
rect 5448 28500 5500 28509
rect 6644 28543 6696 28552
rect 6644 28509 6653 28543
rect 6653 28509 6687 28543
rect 6687 28509 6696 28543
rect 6644 28500 6696 28509
rect 9312 28636 9364 28688
rect 9496 28636 9548 28688
rect 10600 28636 10652 28688
rect 11060 28704 11112 28756
rect 11888 28747 11940 28756
rect 11888 28713 11897 28747
rect 11897 28713 11931 28747
rect 11931 28713 11940 28747
rect 11888 28704 11940 28713
rect 11980 28704 12032 28756
rect 15384 28704 15436 28756
rect 8024 28568 8076 28620
rect 7196 28500 7248 28552
rect 7472 28500 7524 28552
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 5356 28364 5408 28416
rect 6552 28475 6604 28484
rect 6552 28441 6561 28475
rect 6561 28441 6595 28475
rect 6595 28441 6604 28475
rect 6552 28432 6604 28441
rect 9680 28432 9732 28484
rect 10140 28432 10192 28484
rect 10508 28500 10560 28552
rect 11520 28500 11572 28552
rect 11796 28432 11848 28484
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 13452 28636 13504 28688
rect 16488 28704 16540 28756
rect 17684 28747 17736 28756
rect 17684 28713 17693 28747
rect 17693 28713 17727 28747
rect 17727 28713 17736 28747
rect 17684 28704 17736 28713
rect 19800 28747 19852 28756
rect 19800 28713 19809 28747
rect 19809 28713 19843 28747
rect 19843 28713 19852 28747
rect 19800 28704 19852 28713
rect 16764 28636 16816 28688
rect 14740 28543 14792 28552
rect 14740 28509 14749 28543
rect 14749 28509 14783 28543
rect 14783 28509 14792 28543
rect 14740 28500 14792 28509
rect 15108 28500 15160 28552
rect 15200 28543 15252 28552
rect 15200 28509 15209 28543
rect 15209 28509 15243 28543
rect 15243 28509 15252 28543
rect 15200 28500 15252 28509
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 16580 28500 16632 28509
rect 16856 28500 16908 28552
rect 17960 28568 18012 28620
rect 21456 28611 21508 28620
rect 21456 28577 21465 28611
rect 21465 28577 21499 28611
rect 21499 28577 21508 28611
rect 21456 28568 21508 28577
rect 5816 28364 5868 28416
rect 7380 28364 7432 28416
rect 7840 28364 7892 28416
rect 9588 28364 9640 28416
rect 10784 28407 10836 28416
rect 10784 28373 10793 28407
rect 10793 28373 10827 28407
rect 10827 28373 10836 28407
rect 10784 28364 10836 28373
rect 11704 28407 11756 28416
rect 11704 28373 11713 28407
rect 11713 28373 11747 28407
rect 11747 28373 11756 28407
rect 11704 28364 11756 28373
rect 12624 28364 12676 28416
rect 13360 28432 13412 28484
rect 17868 28500 17920 28552
rect 18236 28500 18288 28552
rect 21364 28500 21416 28552
rect 19248 28432 19300 28484
rect 19984 28432 20036 28484
rect 20444 28432 20496 28484
rect 27160 28704 27212 28756
rect 31300 28704 31352 28756
rect 31392 28704 31444 28756
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 23848 28636 23900 28688
rect 24952 28679 25004 28688
rect 24952 28645 24961 28679
rect 24961 28645 24995 28679
rect 24995 28645 25004 28679
rect 24952 28636 25004 28645
rect 25044 28679 25096 28688
rect 25044 28645 25053 28679
rect 25053 28645 25087 28679
rect 25087 28645 25096 28679
rect 25044 28636 25096 28645
rect 23480 28543 23532 28552
rect 23480 28509 23489 28543
rect 23489 28509 23523 28543
rect 23523 28509 23532 28543
rect 23480 28500 23532 28509
rect 26056 28568 26108 28620
rect 24124 28500 24176 28552
rect 27896 28568 27948 28620
rect 21916 28432 21968 28484
rect 22560 28475 22612 28484
rect 22560 28441 22569 28475
rect 22569 28441 22603 28475
rect 22603 28441 22612 28475
rect 22560 28432 22612 28441
rect 23296 28432 23348 28484
rect 14832 28364 14884 28416
rect 14924 28364 14976 28416
rect 21456 28364 21508 28416
rect 21824 28407 21876 28416
rect 21824 28373 21833 28407
rect 21833 28373 21867 28407
rect 21867 28373 21876 28407
rect 21824 28364 21876 28373
rect 22284 28364 22336 28416
rect 22836 28364 22888 28416
rect 27068 28500 27120 28552
rect 27988 28500 28040 28552
rect 28264 28543 28316 28552
rect 28264 28509 28273 28543
rect 28273 28509 28307 28543
rect 28307 28509 28316 28543
rect 28264 28500 28316 28509
rect 24768 28432 24820 28484
rect 25044 28364 25096 28416
rect 27252 28432 27304 28484
rect 27436 28432 27488 28484
rect 31116 28568 31168 28620
rect 29920 28500 29972 28552
rect 31208 28543 31260 28552
rect 31208 28509 31217 28543
rect 31217 28509 31251 28543
rect 31251 28509 31260 28543
rect 31208 28500 31260 28509
rect 31668 28543 31720 28552
rect 31668 28509 31677 28543
rect 31677 28509 31711 28543
rect 31711 28509 31720 28543
rect 31668 28500 31720 28509
rect 31760 28543 31812 28552
rect 31760 28509 31770 28543
rect 31770 28509 31804 28543
rect 31804 28509 31812 28543
rect 31760 28500 31812 28509
rect 32404 28704 32456 28756
rect 33416 28611 33468 28620
rect 33416 28577 33425 28611
rect 33425 28577 33459 28611
rect 33459 28577 33468 28611
rect 33416 28568 33468 28577
rect 33876 28568 33928 28620
rect 35992 28636 36044 28688
rect 33048 28543 33100 28552
rect 33048 28509 33057 28543
rect 33057 28509 33091 28543
rect 33091 28509 33100 28543
rect 33048 28500 33100 28509
rect 35532 28543 35584 28552
rect 35532 28509 35541 28543
rect 35541 28509 35575 28543
rect 35575 28509 35584 28543
rect 35532 28500 35584 28509
rect 36360 28568 36412 28620
rect 27620 28364 27672 28416
rect 31392 28432 31444 28484
rect 32036 28475 32088 28484
rect 32036 28441 32045 28475
rect 32045 28441 32079 28475
rect 32079 28441 32088 28475
rect 32036 28432 32088 28441
rect 28632 28364 28684 28416
rect 29920 28364 29972 28416
rect 35900 28543 35952 28552
rect 35900 28509 35909 28543
rect 35909 28509 35943 28543
rect 35943 28509 35952 28543
rect 35900 28500 35952 28509
rect 36268 28500 36320 28552
rect 36176 28407 36228 28416
rect 36176 28373 36185 28407
rect 36185 28373 36219 28407
rect 36219 28373 36228 28407
rect 36176 28364 36228 28373
rect 37464 28432 37516 28484
rect 37832 28364 37884 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4804 28160 4856 28212
rect 3884 27956 3936 28008
rect 11704 28160 11756 28212
rect 11796 28160 11848 28212
rect 6552 28092 6604 28144
rect 7196 28092 7248 28144
rect 10784 28092 10836 28144
rect 13360 28092 13412 28144
rect 14648 28203 14700 28212
rect 14648 28169 14657 28203
rect 14657 28169 14691 28203
rect 14691 28169 14700 28203
rect 14648 28160 14700 28169
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 20168 28160 20220 28212
rect 5172 28067 5224 28076
rect 5172 28033 5181 28067
rect 5181 28033 5215 28067
rect 5215 28033 5224 28067
rect 5172 28024 5224 28033
rect 5540 28024 5592 28076
rect 9220 28024 9272 28076
rect 10048 28024 10100 28076
rect 10140 28024 10192 28076
rect 10508 28067 10560 28076
rect 10508 28033 10517 28067
rect 10517 28033 10551 28067
rect 10551 28033 10560 28067
rect 10508 28024 10560 28033
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 7104 27956 7156 28008
rect 10600 27956 10652 28008
rect 13360 27999 13412 28008
rect 13360 27965 13369 27999
rect 13369 27965 13403 27999
rect 13403 27965 13412 27999
rect 13360 27956 13412 27965
rect 7748 27888 7800 27940
rect 8300 27888 8352 27940
rect 4804 27863 4856 27872
rect 4804 27829 4813 27863
rect 4813 27829 4847 27863
rect 4847 27829 4856 27863
rect 4804 27820 4856 27829
rect 6552 27820 6604 27872
rect 6828 27863 6880 27872
rect 6828 27829 6837 27863
rect 6837 27829 6871 27863
rect 6871 27829 6880 27863
rect 6828 27820 6880 27829
rect 9220 27820 9272 27872
rect 16488 28024 16540 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 16580 27956 16632 28008
rect 18328 28024 18380 28076
rect 19984 28024 20036 28076
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 20260 27999 20312 28008
rect 20260 27965 20269 27999
rect 20269 27965 20303 27999
rect 20303 27965 20312 27999
rect 20260 27956 20312 27965
rect 20996 28160 21048 28212
rect 24768 28160 24820 28212
rect 24860 28160 24912 28212
rect 25964 28203 26016 28212
rect 25964 28169 25973 28203
rect 25973 28169 26007 28203
rect 26007 28169 26016 28203
rect 25964 28160 26016 28169
rect 27896 28160 27948 28212
rect 28632 28160 28684 28212
rect 30380 28203 30432 28212
rect 30380 28169 30389 28203
rect 30389 28169 30423 28203
rect 30423 28169 30432 28203
rect 30380 28160 30432 28169
rect 20536 28092 20588 28144
rect 22284 28024 22336 28076
rect 22836 28092 22888 28144
rect 23296 28092 23348 28144
rect 24124 28092 24176 28144
rect 25136 28135 25188 28144
rect 25136 28101 25145 28135
rect 25145 28101 25179 28135
rect 25179 28101 25188 28135
rect 25136 28092 25188 28101
rect 23112 28024 23164 28076
rect 23204 28067 23256 28076
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 25044 28024 25096 28076
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 24952 27956 25004 28008
rect 25228 27956 25280 28008
rect 26240 28067 26292 28076
rect 26240 28033 26249 28067
rect 26249 28033 26283 28067
rect 26283 28033 26292 28067
rect 26240 28024 26292 28033
rect 27344 28067 27396 28076
rect 27344 28033 27353 28067
rect 27353 28033 27387 28067
rect 27387 28033 27396 28067
rect 27344 28024 27396 28033
rect 27804 28135 27856 28144
rect 27804 28101 27813 28135
rect 27813 28101 27847 28135
rect 27847 28101 27856 28135
rect 27804 28092 27856 28101
rect 30012 28135 30064 28144
rect 30012 28101 30021 28135
rect 30021 28101 30055 28135
rect 30055 28101 30064 28135
rect 30012 28092 30064 28101
rect 29736 28067 29788 28076
rect 29736 28033 29745 28067
rect 29745 28033 29779 28067
rect 29779 28033 29788 28067
rect 29736 28024 29788 28033
rect 27436 27999 27488 28008
rect 27436 27965 27445 27999
rect 27445 27965 27479 27999
rect 27479 27965 27488 27999
rect 27436 27956 27488 27965
rect 29552 27956 29604 28008
rect 30288 28024 30340 28076
rect 30380 27956 30432 28008
rect 14832 27888 14884 27940
rect 19340 27888 19392 27940
rect 19984 27888 20036 27940
rect 13176 27820 13228 27872
rect 20076 27820 20128 27872
rect 20536 27863 20588 27872
rect 20536 27829 20545 27863
rect 20545 27829 20579 27863
rect 20579 27829 20588 27863
rect 20536 27820 20588 27829
rect 22836 27888 22888 27940
rect 26976 27888 27028 27940
rect 27068 27888 27120 27940
rect 31760 28160 31812 28212
rect 31852 28092 31904 28144
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 32404 28067 32456 28076
rect 32404 28033 32413 28067
rect 32413 28033 32447 28067
rect 32447 28033 32456 28067
rect 32404 28024 32456 28033
rect 34244 28160 34296 28212
rect 37464 28203 37516 28212
rect 37464 28169 37473 28203
rect 37473 28169 37507 28203
rect 37507 28169 37516 28203
rect 37464 28160 37516 28169
rect 37832 28203 37884 28212
rect 37832 28169 37841 28203
rect 37841 28169 37875 28203
rect 37875 28169 37884 28203
rect 37832 28160 37884 28169
rect 33416 28092 33468 28144
rect 36176 28092 36228 28144
rect 33600 28024 33652 28076
rect 32588 27888 32640 27940
rect 23480 27820 23532 27872
rect 26424 27820 26476 27872
rect 27160 27863 27212 27872
rect 27160 27829 27169 27863
rect 27169 27829 27203 27863
rect 27203 27829 27212 27863
rect 27160 27820 27212 27829
rect 27528 27863 27580 27872
rect 27528 27829 27537 27863
rect 27537 27829 27571 27863
rect 27571 27829 27580 27863
rect 27528 27820 27580 27829
rect 33324 27956 33376 28008
rect 38016 27999 38068 28008
rect 38016 27965 38025 27999
rect 38025 27965 38059 27999
rect 38059 27965 38068 27999
rect 38016 27956 38068 27965
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4620 27548 4672 27600
rect 5632 27548 5684 27600
rect 7196 27548 7248 27600
rect 5356 27523 5408 27532
rect 5356 27489 5365 27523
rect 5365 27489 5399 27523
rect 5399 27489 5408 27523
rect 5356 27480 5408 27489
rect 7472 27548 7524 27600
rect 7748 27480 7800 27532
rect 9128 27548 9180 27600
rect 10692 27591 10744 27600
rect 10692 27557 10701 27591
rect 10701 27557 10735 27591
rect 10735 27557 10744 27591
rect 10692 27548 10744 27557
rect 17040 27548 17092 27600
rect 17684 27548 17736 27600
rect 18236 27548 18288 27600
rect 19340 27616 19392 27668
rect 20996 27616 21048 27668
rect 21180 27616 21232 27668
rect 23664 27616 23716 27668
rect 29736 27616 29788 27668
rect 30932 27616 30984 27668
rect 31116 27659 31168 27668
rect 31116 27625 31125 27659
rect 31125 27625 31159 27659
rect 31159 27625 31168 27659
rect 31116 27616 31168 27625
rect 31208 27616 31260 27668
rect 32312 27616 32364 27668
rect 4436 27455 4488 27464
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 4804 27344 4856 27396
rect 5080 27455 5132 27464
rect 5080 27421 5089 27455
rect 5089 27421 5123 27455
rect 5123 27421 5132 27455
rect 5080 27412 5132 27421
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 5724 27412 5776 27464
rect 7104 27455 7156 27464
rect 7104 27421 7113 27455
rect 7113 27421 7147 27455
rect 7147 27421 7156 27455
rect 7104 27412 7156 27421
rect 7840 27412 7892 27464
rect 6184 27344 6236 27396
rect 6276 27344 6328 27396
rect 8300 27412 8352 27464
rect 10232 27480 10284 27532
rect 17960 27480 18012 27532
rect 18604 27480 18656 27532
rect 10784 27412 10836 27464
rect 11888 27412 11940 27464
rect 12348 27455 12400 27464
rect 12348 27421 12357 27455
rect 12357 27421 12391 27455
rect 12391 27421 12400 27455
rect 12348 27412 12400 27421
rect 3976 27319 4028 27328
rect 3976 27285 3985 27319
rect 3985 27285 4019 27319
rect 4019 27285 4028 27319
rect 3976 27276 4028 27285
rect 5080 27276 5132 27328
rect 5540 27276 5592 27328
rect 5908 27276 5960 27328
rect 7748 27319 7800 27328
rect 7748 27285 7757 27319
rect 7757 27285 7791 27319
rect 7791 27285 7800 27319
rect 7748 27276 7800 27285
rect 9036 27276 9088 27328
rect 10324 27387 10376 27396
rect 10324 27353 10333 27387
rect 10333 27353 10367 27387
rect 10367 27353 10376 27387
rect 10324 27344 10376 27353
rect 12808 27344 12860 27396
rect 17132 27412 17184 27464
rect 17408 27344 17460 27396
rect 19064 27412 19116 27464
rect 20444 27480 20496 27532
rect 20076 27412 20128 27464
rect 22928 27548 22980 27600
rect 23204 27548 23256 27600
rect 23572 27591 23624 27600
rect 23572 27557 23581 27591
rect 23581 27557 23615 27591
rect 23615 27557 23624 27591
rect 23572 27548 23624 27557
rect 24124 27548 24176 27600
rect 27804 27548 27856 27600
rect 23480 27480 23532 27532
rect 24860 27480 24912 27532
rect 25780 27480 25832 27532
rect 21824 27412 21876 27464
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 22652 27412 22704 27421
rect 20720 27344 20772 27396
rect 21088 27387 21140 27396
rect 21088 27353 21097 27387
rect 21097 27353 21131 27387
rect 21131 27353 21140 27387
rect 21088 27344 21140 27353
rect 25320 27412 25372 27464
rect 26148 27412 26200 27464
rect 9864 27276 9916 27328
rect 12440 27276 12492 27328
rect 13452 27276 13504 27328
rect 14004 27276 14056 27328
rect 16580 27319 16632 27328
rect 16580 27285 16589 27319
rect 16589 27285 16623 27319
rect 16623 27285 16632 27319
rect 16580 27276 16632 27285
rect 17040 27276 17092 27328
rect 19340 27276 19392 27328
rect 19892 27276 19944 27328
rect 23940 27344 23992 27396
rect 22468 27276 22520 27328
rect 23112 27276 23164 27328
rect 24768 27276 24820 27328
rect 25136 27276 25188 27328
rect 25412 27387 25464 27396
rect 25412 27353 25421 27387
rect 25421 27353 25455 27387
rect 25455 27353 25464 27387
rect 25412 27344 25464 27353
rect 25504 27344 25556 27396
rect 26608 27455 26660 27464
rect 26608 27421 26617 27455
rect 26617 27421 26651 27455
rect 26651 27421 26660 27455
rect 26608 27412 26660 27421
rect 26240 27276 26292 27328
rect 27344 27412 27396 27464
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 30288 27548 30340 27600
rect 31668 27548 31720 27600
rect 33692 27548 33744 27600
rect 35440 27548 35492 27600
rect 26792 27344 26844 27396
rect 29920 27455 29972 27464
rect 29920 27421 29930 27455
rect 29930 27421 29964 27455
rect 29964 27421 29972 27455
rect 29920 27412 29972 27421
rect 30104 27455 30156 27464
rect 30104 27421 30113 27455
rect 30113 27421 30147 27455
rect 30147 27421 30156 27455
rect 30104 27412 30156 27421
rect 30656 27480 30708 27532
rect 33416 27480 33468 27532
rect 33600 27480 33652 27532
rect 27252 27276 27304 27328
rect 27804 27276 27856 27328
rect 30932 27344 30984 27396
rect 32956 27455 33008 27464
rect 32956 27421 32965 27455
rect 32965 27421 32999 27455
rect 32999 27421 33008 27455
rect 32956 27412 33008 27421
rect 33692 27455 33744 27464
rect 33692 27421 33701 27455
rect 33701 27421 33735 27455
rect 33735 27421 33744 27455
rect 33692 27412 33744 27421
rect 33968 27412 34020 27464
rect 34520 27412 34572 27464
rect 34980 27455 35032 27464
rect 34980 27421 34989 27455
rect 34989 27421 35023 27455
rect 35023 27421 35032 27455
rect 34980 27412 35032 27421
rect 35532 27412 35584 27464
rect 38936 27480 38988 27532
rect 30288 27276 30340 27328
rect 32036 27276 32088 27328
rect 33876 27387 33928 27396
rect 33876 27353 33885 27387
rect 33885 27353 33919 27387
rect 33919 27353 33928 27387
rect 33876 27344 33928 27353
rect 37924 27344 37976 27396
rect 39028 27344 39080 27396
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4436 27072 4488 27124
rect 3976 27004 4028 27056
rect 5540 27047 5592 27056
rect 5540 27013 5549 27047
rect 5549 27013 5583 27047
rect 5583 27013 5592 27047
rect 5540 27004 5592 27013
rect 7380 27072 7432 27124
rect 8208 27072 8260 27124
rect 12808 27115 12860 27124
rect 12808 27081 12817 27115
rect 12817 27081 12851 27115
rect 12851 27081 12860 27115
rect 12808 27072 12860 27081
rect 13176 27047 13228 27056
rect 13176 27013 13185 27047
rect 13185 27013 13219 27047
rect 13219 27013 13228 27047
rect 13176 27004 13228 27013
rect 2780 26979 2832 26988
rect 2780 26945 2789 26979
rect 2789 26945 2823 26979
rect 2823 26945 2832 26979
rect 2780 26936 2832 26945
rect 4804 26936 4856 26988
rect 5356 26936 5408 26988
rect 5908 26936 5960 26988
rect 6092 26936 6144 26988
rect 6644 26936 6696 26988
rect 6184 26868 6236 26920
rect 7288 26979 7340 26988
rect 7288 26945 7297 26979
rect 7297 26945 7331 26979
rect 7331 26945 7340 26979
rect 7288 26936 7340 26945
rect 7472 26979 7524 26988
rect 7472 26945 7481 26979
rect 7481 26945 7515 26979
rect 7515 26945 7524 26979
rect 7472 26936 7524 26945
rect 6920 26868 6972 26920
rect 8116 26936 8168 26988
rect 8208 26936 8260 26988
rect 8024 26843 8076 26852
rect 8024 26809 8033 26843
rect 8033 26809 8067 26843
rect 8067 26809 8076 26843
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 8760 26911 8812 26920
rect 8760 26877 8769 26911
rect 8769 26877 8803 26911
rect 8803 26877 8812 26911
rect 8760 26868 8812 26877
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 10232 26979 10284 26988
rect 10232 26945 10241 26979
rect 10241 26945 10275 26979
rect 10275 26945 10284 26979
rect 10232 26936 10284 26945
rect 10508 26936 10560 26988
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 14004 27004 14056 27056
rect 15108 27072 15160 27124
rect 17132 27072 17184 27124
rect 20260 27072 20312 27124
rect 16948 27004 17000 27056
rect 13360 26979 13412 26988
rect 13360 26945 13369 26979
rect 13369 26945 13403 26979
rect 13403 26945 13412 26979
rect 13360 26936 13412 26945
rect 14832 26979 14884 26988
rect 14832 26945 14866 26979
rect 14866 26945 14884 26979
rect 14832 26936 14884 26945
rect 8024 26800 8076 26809
rect 4712 26732 4764 26784
rect 8208 26732 8260 26784
rect 12440 26868 12492 26920
rect 14464 26868 14516 26920
rect 16764 26868 16816 26920
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 18236 26936 18288 26988
rect 19064 27004 19116 27056
rect 19800 26936 19852 26988
rect 18144 26911 18196 26920
rect 18144 26877 18153 26911
rect 18153 26877 18187 26911
rect 18187 26877 18196 26911
rect 18144 26868 18196 26877
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20536 27004 20588 27056
rect 20260 26936 20312 26945
rect 20996 26936 21048 26988
rect 22652 26936 22704 26988
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 14372 26800 14424 26852
rect 17040 26843 17092 26852
rect 17040 26809 17049 26843
rect 17049 26809 17083 26843
rect 17083 26809 17092 26843
rect 17040 26800 17092 26809
rect 17224 26800 17276 26852
rect 18328 26800 18380 26852
rect 20904 26911 20956 26920
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 21732 26868 21784 26920
rect 10232 26775 10284 26784
rect 10232 26741 10241 26775
rect 10241 26741 10275 26775
rect 10275 26741 10284 26775
rect 10232 26732 10284 26741
rect 10416 26732 10468 26784
rect 16396 26732 16448 26784
rect 16488 26732 16540 26784
rect 20720 26732 20772 26784
rect 21088 26732 21140 26784
rect 21548 26732 21600 26784
rect 22100 26732 22152 26784
rect 23020 26775 23072 26784
rect 23020 26741 23029 26775
rect 23029 26741 23063 26775
rect 23063 26741 23072 26775
rect 23020 26732 23072 26741
rect 24584 27115 24636 27124
rect 24584 27081 24593 27115
rect 24593 27081 24627 27115
rect 24627 27081 24636 27115
rect 24584 27072 24636 27081
rect 24952 27072 25004 27124
rect 23940 26979 23992 26988
rect 23940 26945 23949 26979
rect 23949 26945 23983 26979
rect 23983 26945 23992 26979
rect 23940 26936 23992 26945
rect 24124 26979 24176 26988
rect 24124 26945 24133 26979
rect 24133 26945 24167 26979
rect 24167 26945 24176 26979
rect 24124 26936 24176 26945
rect 24768 26979 24820 26988
rect 24768 26945 24777 26979
rect 24777 26945 24811 26979
rect 24811 26945 24820 26979
rect 24768 26936 24820 26945
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 25504 27004 25556 27056
rect 26148 27047 26200 27056
rect 26148 27013 26157 27047
rect 26157 27013 26191 27047
rect 26191 27013 26200 27047
rect 26148 27004 26200 27013
rect 27160 27072 27212 27124
rect 27620 27072 27672 27124
rect 31116 27072 31168 27124
rect 32956 27072 33008 27124
rect 37556 27072 37608 27124
rect 37924 27115 37976 27124
rect 37924 27081 37933 27115
rect 37933 27081 37967 27115
rect 37967 27081 37976 27115
rect 37924 27072 37976 27081
rect 25136 26936 25188 26988
rect 27344 26936 27396 26988
rect 27436 26868 27488 26920
rect 27620 26979 27672 26988
rect 27620 26945 27629 26979
rect 27629 26945 27663 26979
rect 27663 26945 27672 26979
rect 27620 26936 27672 26945
rect 32220 27004 32272 27056
rect 34796 27047 34848 27056
rect 34796 27013 34805 27047
rect 34805 27013 34839 27047
rect 34839 27013 34848 27047
rect 34796 27004 34848 27013
rect 36360 27004 36412 27056
rect 29000 26936 29052 26988
rect 29736 26979 29788 26988
rect 29736 26945 29745 26979
rect 29745 26945 29779 26979
rect 29779 26945 29788 26979
rect 29736 26936 29788 26945
rect 30104 26936 30156 26988
rect 31484 26936 31536 26988
rect 32588 26979 32640 26988
rect 32588 26945 32597 26979
rect 32597 26945 32631 26979
rect 32631 26945 32640 26979
rect 32588 26936 32640 26945
rect 33048 26936 33100 26988
rect 34152 26979 34204 26988
rect 34152 26945 34161 26979
rect 34161 26945 34195 26979
rect 34195 26945 34204 26979
rect 34152 26936 34204 26945
rect 34704 26936 34756 26988
rect 37832 26979 37884 26988
rect 37832 26945 37841 26979
rect 37841 26945 37875 26979
rect 37875 26945 37884 26979
rect 37832 26936 37884 26945
rect 31392 26868 31444 26920
rect 32680 26868 32732 26920
rect 33324 26911 33376 26920
rect 33324 26877 33333 26911
rect 33333 26877 33367 26911
rect 33367 26877 33376 26911
rect 33324 26868 33376 26877
rect 33416 26868 33468 26920
rect 38108 26868 38160 26920
rect 23572 26800 23624 26852
rect 24860 26800 24912 26852
rect 24952 26843 25004 26852
rect 24952 26809 24961 26843
rect 24961 26809 24995 26843
rect 24995 26809 25004 26843
rect 24952 26800 25004 26809
rect 32956 26800 33008 26852
rect 34980 26800 35032 26852
rect 35808 26800 35860 26852
rect 25044 26732 25096 26784
rect 26332 26775 26384 26784
rect 26332 26741 26341 26775
rect 26341 26741 26375 26775
rect 26375 26741 26384 26775
rect 26332 26732 26384 26741
rect 36268 26732 36320 26784
rect 36820 26732 36872 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8116 26528 8168 26580
rect 10324 26528 10376 26580
rect 12256 26528 12308 26580
rect 14832 26528 14884 26580
rect 16396 26528 16448 26580
rect 19432 26528 19484 26580
rect 23020 26528 23072 26580
rect 23664 26528 23716 26580
rect 25872 26528 25924 26580
rect 26516 26528 26568 26580
rect 6368 26460 6420 26512
rect 10416 26460 10468 26512
rect 14096 26460 14148 26512
rect 5448 26392 5500 26444
rect 8392 26392 8444 26444
rect 14372 26392 14424 26444
rect 17224 26392 17276 26444
rect 4896 26324 4948 26376
rect 5632 26324 5684 26376
rect 5908 26367 5960 26376
rect 5908 26333 5917 26367
rect 5917 26333 5951 26367
rect 5951 26333 5960 26367
rect 5908 26324 5960 26333
rect 6092 26367 6144 26376
rect 6092 26333 6101 26367
rect 6101 26333 6135 26367
rect 6135 26333 6144 26367
rect 6092 26324 6144 26333
rect 8300 26367 8352 26376
rect 8300 26333 8309 26367
rect 8309 26333 8343 26367
rect 8343 26333 8352 26367
rect 8300 26324 8352 26333
rect 8760 26324 8812 26376
rect 5724 26256 5776 26308
rect 6184 26256 6236 26308
rect 4620 26188 4672 26240
rect 9496 26299 9548 26308
rect 9496 26265 9505 26299
rect 9505 26265 9539 26299
rect 9539 26265 9548 26299
rect 9496 26256 9548 26265
rect 11152 26256 11204 26308
rect 15108 26367 15160 26376
rect 15108 26333 15117 26367
rect 15117 26333 15151 26367
rect 15151 26333 15160 26367
rect 15108 26324 15160 26333
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 17960 26392 18012 26444
rect 20444 26460 20496 26512
rect 21272 26460 21324 26512
rect 21456 26460 21508 26512
rect 21732 26460 21784 26512
rect 13636 26256 13688 26308
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 20352 26392 20404 26444
rect 18328 26324 18380 26376
rect 17224 26256 17276 26308
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 19800 26324 19852 26376
rect 20536 26324 20588 26376
rect 21640 26392 21692 26444
rect 21180 26324 21232 26376
rect 21456 26324 21508 26376
rect 23848 26392 23900 26444
rect 24032 26460 24084 26512
rect 22008 26367 22060 26376
rect 22008 26333 22017 26367
rect 22017 26333 22051 26367
rect 22051 26333 22060 26367
rect 22008 26324 22060 26333
rect 22836 26367 22888 26376
rect 22836 26333 22845 26367
rect 22845 26333 22879 26367
rect 22879 26333 22888 26367
rect 22836 26324 22888 26333
rect 23388 26324 23440 26376
rect 23572 26324 23624 26376
rect 23664 26367 23716 26376
rect 23664 26333 23673 26367
rect 23673 26333 23707 26367
rect 23707 26333 23716 26367
rect 23664 26324 23716 26333
rect 9312 26231 9364 26240
rect 9312 26197 9339 26231
rect 9339 26197 9364 26231
rect 9312 26188 9364 26197
rect 9772 26188 9824 26240
rect 10968 26188 11020 26240
rect 12532 26188 12584 26240
rect 18052 26231 18104 26240
rect 18052 26197 18061 26231
rect 18061 26197 18095 26231
rect 18095 26197 18104 26231
rect 18052 26188 18104 26197
rect 18144 26188 18196 26240
rect 19708 26188 19760 26240
rect 20076 26188 20128 26240
rect 22008 26188 22060 26240
rect 22376 26188 22428 26240
rect 24676 26256 24728 26308
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 25044 26367 25096 26376
rect 25044 26333 25053 26367
rect 25053 26333 25087 26367
rect 25087 26333 25096 26367
rect 25044 26324 25096 26333
rect 25136 26367 25188 26376
rect 25136 26333 25145 26367
rect 25145 26333 25179 26367
rect 25179 26333 25188 26367
rect 25136 26324 25188 26333
rect 26332 26460 26384 26512
rect 27712 26460 27764 26512
rect 27988 26460 28040 26512
rect 26792 26256 26844 26308
rect 27896 26367 27948 26376
rect 27896 26333 27905 26367
rect 27905 26333 27939 26367
rect 27939 26333 27948 26367
rect 27896 26324 27948 26333
rect 27988 26367 28040 26376
rect 27988 26333 27997 26367
rect 27997 26333 28031 26367
rect 28031 26333 28040 26367
rect 27988 26324 28040 26333
rect 28264 26503 28316 26512
rect 28264 26469 28273 26503
rect 28273 26469 28307 26503
rect 28307 26469 28316 26503
rect 28264 26460 28316 26469
rect 29552 26528 29604 26580
rect 33876 26528 33928 26580
rect 29920 26460 29972 26512
rect 30196 26392 30248 26444
rect 28540 26324 28592 26376
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 32680 26460 32732 26512
rect 33600 26460 33652 26512
rect 34152 26460 34204 26512
rect 34244 26460 34296 26512
rect 35532 26571 35584 26580
rect 35532 26537 35541 26571
rect 35541 26537 35575 26571
rect 35575 26537 35584 26571
rect 35532 26528 35584 26537
rect 37832 26528 37884 26580
rect 33416 26435 33468 26444
rect 33416 26401 33425 26435
rect 33425 26401 33459 26435
rect 33459 26401 33468 26435
rect 33416 26392 33468 26401
rect 34520 26392 34572 26444
rect 33968 26324 34020 26376
rect 34060 26367 34112 26376
rect 34060 26333 34069 26367
rect 34069 26333 34103 26367
rect 34103 26333 34112 26367
rect 34060 26324 34112 26333
rect 34244 26367 34296 26376
rect 34244 26333 34253 26367
rect 34253 26333 34287 26367
rect 34287 26333 34296 26367
rect 34244 26324 34296 26333
rect 34980 26367 35032 26376
rect 34980 26333 34989 26367
rect 34989 26333 35023 26367
rect 35023 26333 35032 26367
rect 34980 26324 35032 26333
rect 36360 26392 36412 26444
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 36820 26367 36872 26376
rect 36820 26333 36854 26367
rect 36854 26333 36872 26367
rect 36820 26324 36872 26333
rect 29552 26256 29604 26308
rect 22928 26188 22980 26240
rect 30196 26231 30248 26240
rect 30196 26197 30205 26231
rect 30205 26197 30239 26231
rect 30239 26197 30248 26231
rect 30196 26188 30248 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4896 25984 4948 26036
rect 6920 25984 6972 26036
rect 10600 25984 10652 26036
rect 11152 26027 11204 26036
rect 11152 25993 11161 26027
rect 11161 25993 11195 26027
rect 11195 25993 11204 26027
rect 11152 25984 11204 25993
rect 5264 25916 5316 25968
rect 12256 25916 12308 25968
rect 12440 25916 12492 25968
rect 4804 25848 4856 25900
rect 5540 25848 5592 25900
rect 5816 25848 5868 25900
rect 6644 25891 6696 25900
rect 6644 25857 6653 25891
rect 6653 25857 6687 25891
rect 6687 25857 6696 25891
rect 6644 25848 6696 25857
rect 6828 25891 6880 25900
rect 6828 25857 6837 25891
rect 6837 25857 6871 25891
rect 6871 25857 6880 25891
rect 6828 25848 6880 25857
rect 7288 25848 7340 25900
rect 8116 25891 8168 25900
rect 8116 25857 8125 25891
rect 8125 25857 8159 25891
rect 8159 25857 8168 25891
rect 8116 25848 8168 25857
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 9496 25848 9548 25900
rect 5172 25780 5224 25832
rect 5908 25780 5960 25832
rect 9404 25780 9456 25832
rect 9772 25823 9824 25832
rect 9772 25789 9781 25823
rect 9781 25789 9815 25823
rect 9815 25789 9824 25823
rect 9772 25780 9824 25789
rect 5816 25712 5868 25764
rect 6644 25712 6696 25764
rect 8300 25712 8352 25764
rect 10232 25848 10284 25900
rect 10416 25848 10468 25900
rect 10692 25848 10744 25900
rect 10968 25891 11020 25900
rect 10968 25857 10977 25891
rect 10977 25857 11011 25891
rect 11011 25857 11020 25891
rect 10968 25848 11020 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 12532 25780 12584 25832
rect 11980 25712 12032 25764
rect 4896 25644 4948 25696
rect 9956 25687 10008 25696
rect 9956 25653 9965 25687
rect 9965 25653 9999 25687
rect 9999 25653 10008 25687
rect 9956 25644 10008 25653
rect 10232 25644 10284 25696
rect 10324 25644 10376 25696
rect 14096 25984 14148 26036
rect 18052 25984 18104 26036
rect 19892 25984 19944 26036
rect 21364 25984 21416 26036
rect 16948 25916 17000 25968
rect 19340 25916 19392 25968
rect 20260 25916 20312 25968
rect 20720 25916 20772 25968
rect 21732 25916 21784 25968
rect 12992 25891 13044 25900
rect 12992 25857 13001 25891
rect 13001 25857 13035 25891
rect 13035 25857 13044 25891
rect 12992 25848 13044 25857
rect 13636 25848 13688 25900
rect 15200 25848 15252 25900
rect 17684 25848 17736 25900
rect 18144 25891 18196 25900
rect 18144 25857 18153 25891
rect 18153 25857 18187 25891
rect 18187 25857 18196 25891
rect 18144 25848 18196 25857
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 22100 25848 22152 25900
rect 17316 25780 17368 25832
rect 17776 25780 17828 25832
rect 20076 25823 20128 25832
rect 20076 25789 20085 25823
rect 20085 25789 20119 25823
rect 20119 25789 20128 25823
rect 20076 25780 20128 25789
rect 17500 25712 17552 25764
rect 13176 25687 13228 25696
rect 13176 25653 13185 25687
rect 13185 25653 13219 25687
rect 13219 25653 13228 25687
rect 13176 25644 13228 25653
rect 17776 25644 17828 25696
rect 18144 25712 18196 25764
rect 20812 25780 20864 25832
rect 26240 25984 26292 26036
rect 22744 25916 22796 25968
rect 27620 25916 27672 25968
rect 27896 25959 27948 25968
rect 27896 25925 27905 25959
rect 27905 25925 27939 25959
rect 27939 25925 27948 25959
rect 27896 25916 27948 25925
rect 23296 25891 23348 25900
rect 23296 25857 23305 25891
rect 23305 25857 23339 25891
rect 23339 25857 23348 25891
rect 23296 25848 23348 25857
rect 23756 25848 23808 25900
rect 25136 25848 25188 25900
rect 27712 25891 27764 25900
rect 27712 25857 27721 25891
rect 27721 25857 27755 25891
rect 27755 25857 27764 25891
rect 27712 25848 27764 25857
rect 24860 25780 24912 25832
rect 23296 25755 23348 25764
rect 23296 25721 23305 25755
rect 23305 25721 23339 25755
rect 23339 25721 23348 25755
rect 23296 25712 23348 25721
rect 20904 25644 20956 25696
rect 27528 25687 27580 25696
rect 27528 25653 27537 25687
rect 27537 25653 27571 25687
rect 27571 25653 27580 25687
rect 27528 25644 27580 25653
rect 32404 25984 32456 26036
rect 33692 25984 33744 26036
rect 29000 25959 29052 25968
rect 29000 25925 29009 25959
rect 29009 25925 29043 25959
rect 29043 25925 29052 25959
rect 29000 25916 29052 25925
rect 33140 25916 33192 25968
rect 29460 25848 29512 25900
rect 30196 25891 30248 25900
rect 30196 25857 30205 25891
rect 30205 25857 30239 25891
rect 30239 25857 30248 25891
rect 30196 25848 30248 25857
rect 30656 25891 30708 25900
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 30656 25848 30708 25857
rect 30748 25891 30800 25900
rect 30748 25857 30757 25891
rect 30757 25857 30791 25891
rect 30791 25857 30800 25891
rect 30748 25848 30800 25857
rect 30288 25780 30340 25832
rect 31024 25891 31076 25900
rect 31024 25857 31033 25891
rect 31033 25857 31067 25891
rect 31067 25857 31076 25891
rect 31024 25848 31076 25857
rect 33876 25848 33928 25900
rect 34980 25984 35032 26036
rect 36268 25916 36320 25968
rect 31668 25780 31720 25832
rect 33784 25780 33836 25832
rect 37924 25848 37976 25900
rect 36728 25780 36780 25832
rect 39028 25780 39080 25832
rect 32036 25712 32088 25764
rect 30748 25644 30800 25696
rect 33416 25644 33468 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5632 25440 5684 25492
rect 6920 25440 6972 25492
rect 9312 25440 9364 25492
rect 12992 25440 13044 25492
rect 17684 25440 17736 25492
rect 24308 25440 24360 25492
rect 25320 25440 25372 25492
rect 28080 25440 28132 25492
rect 5080 25372 5132 25424
rect 10324 25372 10376 25424
rect 4620 25304 4672 25356
rect 4896 25347 4948 25356
rect 4896 25313 4905 25347
rect 4905 25313 4939 25347
rect 4939 25313 4948 25347
rect 4896 25304 4948 25313
rect 5264 25347 5316 25356
rect 5264 25313 5273 25347
rect 5273 25313 5307 25347
rect 5307 25313 5316 25347
rect 5264 25304 5316 25313
rect 5356 25347 5408 25356
rect 5356 25313 5365 25347
rect 5365 25313 5399 25347
rect 5399 25313 5408 25347
rect 5356 25304 5408 25313
rect 8208 25304 8260 25356
rect 10140 25304 10192 25356
rect 4620 25168 4672 25220
rect 6736 25279 6788 25288
rect 6736 25245 6745 25279
rect 6745 25245 6779 25279
rect 6779 25245 6788 25279
rect 6736 25236 6788 25245
rect 9680 25236 9732 25288
rect 10600 25236 10652 25288
rect 12348 25279 12400 25288
rect 12348 25245 12357 25279
rect 12357 25245 12391 25279
rect 12391 25245 12400 25279
rect 12348 25236 12400 25245
rect 13176 25236 13228 25288
rect 7840 25168 7892 25220
rect 8208 25168 8260 25220
rect 8300 25168 8352 25220
rect 9956 25168 10008 25220
rect 12532 25168 12584 25220
rect 19892 25372 19944 25424
rect 20076 25372 20128 25424
rect 24860 25372 24912 25424
rect 25504 25372 25556 25424
rect 13636 25304 13688 25356
rect 13452 25236 13504 25288
rect 18052 25304 18104 25356
rect 18328 25304 18380 25356
rect 19064 25304 19116 25356
rect 15752 25236 15804 25288
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 3976 25143 4028 25152
rect 3976 25109 3985 25143
rect 3985 25109 4019 25143
rect 4019 25109 4028 25143
rect 3976 25100 4028 25109
rect 5540 25143 5592 25152
rect 5540 25109 5549 25143
rect 5549 25109 5583 25143
rect 5583 25109 5592 25143
rect 5540 25100 5592 25109
rect 7104 25100 7156 25152
rect 8484 25100 8536 25152
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 18144 25236 18196 25288
rect 16764 25168 16816 25220
rect 14004 25100 14056 25152
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 18696 25279 18748 25288
rect 18696 25245 18705 25279
rect 18705 25245 18739 25279
rect 18739 25245 18748 25279
rect 18696 25236 18748 25245
rect 20260 25304 20312 25356
rect 19984 25279 20036 25288
rect 19984 25245 19993 25279
rect 19993 25245 20027 25279
rect 20027 25245 20036 25279
rect 24492 25304 24544 25356
rect 27712 25372 27764 25424
rect 28540 25372 28592 25424
rect 19984 25236 20036 25245
rect 20536 25279 20588 25288
rect 20536 25245 20545 25279
rect 20545 25245 20579 25279
rect 20579 25245 20588 25279
rect 20536 25236 20588 25245
rect 21180 25236 21232 25288
rect 23112 25279 23164 25288
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 25136 25279 25188 25288
rect 25136 25245 25145 25279
rect 25145 25245 25179 25279
rect 25179 25245 25188 25279
rect 25136 25236 25188 25245
rect 26240 25279 26292 25288
rect 26240 25245 26249 25279
rect 26249 25245 26283 25279
rect 26283 25245 26292 25279
rect 26240 25236 26292 25245
rect 26516 25279 26568 25288
rect 26516 25245 26525 25279
rect 26525 25245 26559 25279
rect 26559 25245 26568 25279
rect 26516 25236 26568 25245
rect 26884 25236 26936 25288
rect 27252 25279 27304 25288
rect 27252 25245 27261 25279
rect 27261 25245 27295 25279
rect 27295 25245 27304 25279
rect 27252 25236 27304 25245
rect 28080 25236 28132 25288
rect 30564 25304 30616 25356
rect 31024 25304 31076 25356
rect 20904 25168 20956 25220
rect 24952 25211 25004 25220
rect 24952 25177 24961 25211
rect 24961 25177 24995 25211
rect 24995 25177 25004 25211
rect 24952 25168 25004 25177
rect 19432 25100 19484 25152
rect 20628 25100 20680 25152
rect 22100 25100 22152 25152
rect 24124 25100 24176 25152
rect 28632 25168 28684 25220
rect 31852 25236 31904 25288
rect 32036 25279 32088 25288
rect 32036 25245 32046 25279
rect 32046 25245 32080 25279
rect 32080 25245 32088 25279
rect 32312 25304 32364 25356
rect 32036 25236 32088 25245
rect 33416 25279 33468 25288
rect 33416 25245 33425 25279
rect 33425 25245 33459 25279
rect 33459 25245 33468 25279
rect 33416 25236 33468 25245
rect 33600 25279 33652 25288
rect 33600 25245 33609 25279
rect 33609 25245 33643 25279
rect 33643 25245 33652 25279
rect 33600 25236 33652 25245
rect 34796 25236 34848 25288
rect 36728 25236 36780 25288
rect 30104 25168 30156 25220
rect 30288 25211 30340 25220
rect 30288 25177 30297 25211
rect 30297 25177 30331 25211
rect 30331 25177 30340 25211
rect 30288 25168 30340 25177
rect 32220 25211 32272 25220
rect 32220 25177 32229 25211
rect 32229 25177 32263 25211
rect 32263 25177 32272 25211
rect 32220 25168 32272 25177
rect 32496 25168 32548 25220
rect 37464 25168 37516 25220
rect 25964 25143 26016 25152
rect 25964 25109 25973 25143
rect 25973 25109 26007 25143
rect 26007 25109 26016 25143
rect 25964 25100 26016 25109
rect 29000 25143 29052 25152
rect 29000 25109 29009 25143
rect 29009 25109 29043 25143
rect 29043 25109 29052 25143
rect 29000 25100 29052 25109
rect 31944 25100 31996 25152
rect 34060 25100 34112 25152
rect 38016 25143 38068 25152
rect 38016 25109 38025 25143
rect 38025 25109 38059 25143
rect 38059 25109 38068 25143
rect 38016 25100 38068 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7656 24896 7708 24948
rect 3976 24828 4028 24880
rect 5540 24828 5592 24880
rect 7840 24828 7892 24880
rect 19248 24939 19300 24948
rect 19248 24905 19257 24939
rect 19257 24905 19291 24939
rect 19291 24905 19300 24939
rect 19248 24896 19300 24905
rect 24308 24939 24360 24948
rect 24308 24905 24317 24939
rect 24317 24905 24351 24939
rect 24351 24905 24360 24939
rect 24308 24896 24360 24905
rect 37464 24939 37516 24948
rect 37464 24905 37473 24939
rect 37473 24905 37507 24939
rect 37507 24905 37516 24939
rect 37464 24896 37516 24905
rect 8484 24828 8536 24880
rect 2780 24803 2832 24812
rect 2780 24769 2789 24803
rect 2789 24769 2823 24803
rect 2823 24769 2832 24803
rect 2780 24760 2832 24769
rect 5632 24760 5684 24812
rect 6920 24760 6972 24812
rect 9772 24828 9824 24880
rect 9680 24760 9732 24812
rect 10416 24871 10468 24880
rect 10416 24837 10425 24871
rect 10425 24837 10459 24871
rect 10459 24837 10468 24871
rect 10416 24828 10468 24837
rect 13452 24871 13504 24880
rect 13452 24837 13461 24871
rect 13461 24837 13495 24871
rect 13495 24837 13504 24871
rect 13452 24828 13504 24837
rect 10508 24803 10560 24812
rect 10508 24769 10517 24803
rect 10517 24769 10551 24803
rect 10551 24769 10560 24803
rect 10508 24760 10560 24769
rect 5172 24735 5224 24744
rect 5172 24701 5181 24735
rect 5181 24701 5215 24735
rect 5215 24701 5224 24735
rect 5172 24692 5224 24701
rect 4988 24624 5040 24676
rect 5448 24692 5500 24744
rect 4620 24556 4672 24608
rect 6736 24624 6788 24676
rect 9772 24692 9824 24744
rect 10416 24692 10468 24744
rect 12440 24760 12492 24812
rect 12716 24624 12768 24676
rect 9496 24556 9548 24608
rect 9588 24599 9640 24608
rect 9588 24565 9597 24599
rect 9597 24565 9631 24599
rect 9631 24565 9640 24599
rect 9588 24556 9640 24565
rect 10876 24556 10928 24608
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 18052 24803 18104 24812
rect 18052 24769 18061 24803
rect 18061 24769 18095 24803
rect 18095 24769 18104 24803
rect 18052 24760 18104 24769
rect 19340 24828 19392 24880
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 20536 24828 20588 24880
rect 21272 24871 21324 24880
rect 21272 24837 21281 24871
rect 21281 24837 21315 24871
rect 21315 24837 21324 24871
rect 21272 24828 21324 24837
rect 22744 24828 22796 24880
rect 20444 24760 20496 24812
rect 21916 24760 21968 24812
rect 13912 24692 13964 24744
rect 14464 24692 14516 24744
rect 16580 24692 16632 24744
rect 23112 24803 23164 24812
rect 23112 24769 23121 24803
rect 23121 24769 23155 24803
rect 23155 24769 23164 24803
rect 23112 24760 23164 24769
rect 23296 24803 23348 24812
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 23388 24760 23440 24812
rect 25688 24828 25740 24880
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 24584 24803 24636 24812
rect 24584 24769 24593 24803
rect 24593 24769 24627 24803
rect 24627 24769 24636 24803
rect 24584 24760 24636 24769
rect 24952 24760 25004 24812
rect 24768 24692 24820 24744
rect 25136 24692 25188 24744
rect 27712 24760 27764 24812
rect 27896 24803 27948 24812
rect 27896 24769 27905 24803
rect 27905 24769 27939 24803
rect 27939 24769 27948 24803
rect 27896 24760 27948 24769
rect 29000 24803 29052 24812
rect 29000 24769 29009 24803
rect 29009 24769 29043 24803
rect 29043 24769 29052 24803
rect 29000 24760 29052 24769
rect 29460 24803 29512 24812
rect 29460 24769 29469 24803
rect 29469 24769 29503 24803
rect 29503 24769 29512 24803
rect 29460 24760 29512 24769
rect 29920 24760 29972 24812
rect 30932 24828 30984 24880
rect 32036 24828 32088 24880
rect 38016 24828 38068 24880
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 30380 24760 30432 24769
rect 33692 24760 33744 24812
rect 26148 24692 26200 24744
rect 28540 24692 28592 24744
rect 28816 24735 28868 24744
rect 28816 24701 28825 24735
rect 28825 24701 28859 24735
rect 28859 24701 28868 24735
rect 28816 24692 28868 24701
rect 31300 24692 31352 24744
rect 33876 24735 33928 24744
rect 33876 24701 33885 24735
rect 33885 24701 33919 24735
rect 33919 24701 33928 24735
rect 33876 24692 33928 24701
rect 26240 24624 26292 24676
rect 26424 24624 26476 24676
rect 18420 24599 18472 24608
rect 18420 24565 18429 24599
rect 18429 24565 18463 24599
rect 18463 24565 18472 24599
rect 18420 24556 18472 24565
rect 27620 24556 27672 24608
rect 28632 24624 28684 24676
rect 29552 24624 29604 24676
rect 29920 24624 29972 24676
rect 32680 24624 32732 24676
rect 37924 24735 37976 24744
rect 37924 24701 37933 24735
rect 37933 24701 37967 24735
rect 37967 24701 37976 24735
rect 37924 24692 37976 24701
rect 38108 24735 38160 24744
rect 38108 24701 38117 24735
rect 38117 24701 38151 24735
rect 38151 24701 38160 24735
rect 38108 24692 38160 24701
rect 30012 24556 30064 24608
rect 35992 24556 36044 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 5172 24352 5224 24404
rect 6000 24352 6052 24404
rect 10508 24352 10560 24404
rect 5724 24284 5776 24336
rect 12072 24352 12124 24404
rect 16856 24352 16908 24404
rect 23204 24395 23256 24404
rect 23204 24361 23213 24395
rect 23213 24361 23247 24395
rect 23247 24361 23256 24395
rect 23204 24352 23256 24361
rect 5356 24216 5408 24268
rect 5632 24216 5684 24268
rect 18696 24284 18748 24336
rect 5724 24191 5776 24200
rect 5724 24157 5733 24191
rect 5733 24157 5767 24191
rect 5767 24157 5776 24191
rect 5724 24148 5776 24157
rect 5816 24191 5868 24200
rect 5816 24157 5825 24191
rect 5825 24157 5859 24191
rect 5859 24157 5868 24191
rect 5816 24148 5868 24157
rect 6552 24148 6604 24200
rect 8024 24216 8076 24268
rect 9404 24259 9456 24268
rect 9404 24225 9413 24259
rect 9413 24225 9447 24259
rect 9447 24225 9456 24259
rect 9404 24216 9456 24225
rect 9588 24259 9640 24268
rect 9588 24225 9597 24259
rect 9597 24225 9631 24259
rect 9631 24225 9640 24259
rect 9588 24216 9640 24225
rect 16856 24216 16908 24268
rect 8116 24148 8168 24200
rect 10324 24148 10376 24200
rect 12348 24148 12400 24200
rect 17316 24148 17368 24200
rect 17408 24191 17460 24200
rect 17408 24157 17417 24191
rect 17417 24157 17451 24191
rect 17451 24157 17460 24191
rect 17408 24148 17460 24157
rect 17776 24191 17828 24200
rect 17776 24157 17785 24191
rect 17785 24157 17819 24191
rect 17819 24157 17828 24191
rect 17776 24148 17828 24157
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 18788 24148 18840 24200
rect 20812 24259 20864 24268
rect 20812 24225 20821 24259
rect 20821 24225 20855 24259
rect 20855 24225 20864 24259
rect 20812 24216 20864 24225
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 21732 24148 21784 24200
rect 22652 24216 22704 24268
rect 4620 24080 4672 24132
rect 10876 24123 10928 24132
rect 6184 24055 6236 24064
rect 6184 24021 6193 24055
rect 6193 24021 6227 24055
rect 6227 24021 6236 24055
rect 6184 24012 6236 24021
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 7012 24055 7064 24064
rect 7012 24021 7021 24055
rect 7021 24021 7055 24055
rect 7055 24021 7064 24055
rect 7012 24012 7064 24021
rect 7656 24012 7708 24064
rect 7840 24012 7892 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 10876 24089 10910 24123
rect 10910 24089 10928 24123
rect 10876 24080 10928 24089
rect 15292 24080 15344 24132
rect 19340 24080 19392 24132
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 23204 24216 23256 24268
rect 24124 24352 24176 24404
rect 24308 24352 24360 24404
rect 23388 24216 23440 24268
rect 25228 24284 25280 24336
rect 26148 24284 26200 24336
rect 27620 24352 27672 24404
rect 23848 24191 23900 24200
rect 23848 24157 23857 24191
rect 23857 24157 23891 24191
rect 23891 24157 23900 24191
rect 23848 24148 23900 24157
rect 24400 24216 24452 24268
rect 25780 24216 25832 24268
rect 24676 24148 24728 24200
rect 26884 24148 26936 24200
rect 29368 24284 29420 24336
rect 27896 24148 27948 24200
rect 28724 24216 28776 24268
rect 28632 24148 28684 24200
rect 29552 24148 29604 24200
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 30380 24352 30432 24404
rect 33784 24352 33836 24404
rect 34244 24352 34296 24404
rect 34704 24352 34756 24404
rect 31852 24284 31904 24336
rect 31208 24191 31260 24200
rect 31208 24157 31217 24191
rect 31217 24157 31251 24191
rect 31251 24157 31260 24191
rect 31208 24148 31260 24157
rect 31484 24216 31536 24268
rect 32036 24216 32088 24268
rect 32404 24259 32456 24268
rect 32404 24225 32413 24259
rect 32413 24225 32447 24259
rect 32447 24225 32456 24259
rect 32404 24216 32456 24225
rect 23388 24080 23440 24132
rect 12072 24012 12124 24064
rect 20260 24055 20312 24064
rect 20260 24021 20269 24055
rect 20269 24021 20303 24055
rect 20303 24021 20312 24055
rect 20260 24012 20312 24021
rect 21088 24012 21140 24064
rect 22836 24055 22888 24064
rect 22836 24021 22845 24055
rect 22845 24021 22879 24055
rect 22879 24021 22888 24055
rect 22836 24012 22888 24021
rect 23296 24012 23348 24064
rect 27160 24080 27212 24132
rect 27712 24080 27764 24132
rect 24768 24055 24820 24064
rect 24768 24021 24777 24055
rect 24777 24021 24811 24055
rect 24811 24021 24820 24055
rect 24768 24012 24820 24021
rect 27988 24012 28040 24064
rect 28172 24123 28224 24132
rect 28172 24089 28181 24123
rect 28181 24089 28215 24123
rect 28215 24089 28224 24123
rect 28172 24080 28224 24089
rect 28816 24080 28868 24132
rect 29736 24080 29788 24132
rect 30012 24080 30064 24132
rect 29276 24012 29328 24064
rect 30840 24012 30892 24064
rect 31300 24012 31352 24064
rect 32312 24191 32364 24200
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 32312 24148 32364 24157
rect 33692 24216 33744 24268
rect 33876 24148 33928 24200
rect 34060 24148 34112 24200
rect 37832 24191 37884 24200
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 39028 24080 39080 24132
rect 32036 24012 32088 24064
rect 32496 24012 32548 24064
rect 37924 24012 37976 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4896 23808 4948 23860
rect 17960 23808 18012 23860
rect 21456 23808 21508 23860
rect 29920 23808 29972 23860
rect 32864 23808 32916 23860
rect 4068 23740 4120 23792
rect 2780 23715 2832 23724
rect 2780 23681 2789 23715
rect 2789 23681 2823 23715
rect 2823 23681 2832 23715
rect 2780 23672 2832 23681
rect 3976 23672 4028 23724
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 4988 23672 5040 23724
rect 5540 23740 5592 23792
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5908 23740 5960 23792
rect 6000 23740 6052 23792
rect 7012 23740 7064 23792
rect 7840 23740 7892 23792
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 9128 23740 9180 23792
rect 12348 23740 12400 23792
rect 13912 23740 13964 23792
rect 18236 23740 18288 23792
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 17224 23672 17276 23724
rect 19432 23672 19484 23724
rect 21272 23740 21324 23792
rect 22192 23740 22244 23792
rect 20812 23672 20864 23724
rect 23112 23672 23164 23724
rect 23388 23715 23440 23724
rect 23388 23681 23397 23715
rect 23397 23681 23431 23715
rect 23431 23681 23440 23715
rect 23388 23672 23440 23681
rect 17132 23604 17184 23656
rect 21640 23604 21692 23656
rect 24768 23715 24820 23724
rect 24768 23681 24777 23715
rect 24777 23681 24811 23715
rect 24811 23681 24820 23715
rect 24768 23672 24820 23681
rect 26240 23740 26292 23792
rect 27988 23783 28040 23792
rect 27988 23749 27997 23783
rect 27997 23749 28031 23783
rect 28031 23749 28040 23783
rect 27988 23740 28040 23749
rect 27712 23715 27764 23724
rect 27712 23681 27721 23715
rect 27721 23681 27755 23715
rect 27755 23681 27764 23715
rect 27712 23672 27764 23681
rect 28632 23715 28684 23724
rect 28632 23681 28641 23715
rect 28641 23681 28675 23715
rect 28675 23681 28684 23715
rect 28632 23672 28684 23681
rect 24584 23604 24636 23656
rect 4620 23511 4672 23520
rect 4620 23477 4629 23511
rect 4629 23477 4663 23511
rect 4663 23477 4672 23511
rect 4620 23468 4672 23477
rect 8576 23468 8628 23520
rect 9772 23511 9824 23520
rect 9772 23477 9781 23511
rect 9781 23477 9815 23511
rect 9815 23477 9824 23511
rect 16304 23536 16356 23588
rect 20352 23579 20404 23588
rect 20352 23545 20361 23579
rect 20361 23545 20395 23579
rect 20395 23545 20404 23579
rect 20352 23536 20404 23545
rect 20628 23536 20680 23588
rect 23480 23579 23532 23588
rect 23480 23545 23489 23579
rect 23489 23545 23523 23579
rect 23523 23545 23532 23579
rect 23480 23536 23532 23545
rect 9772 23468 9824 23477
rect 16948 23468 17000 23520
rect 20720 23511 20772 23520
rect 20720 23477 20729 23511
rect 20729 23477 20763 23511
rect 20763 23477 20772 23511
rect 20720 23468 20772 23477
rect 25136 23536 25188 23588
rect 26148 23647 26200 23656
rect 26148 23613 26157 23647
rect 26157 23613 26191 23647
rect 26191 23613 26200 23647
rect 26148 23604 26200 23613
rect 27344 23604 27396 23656
rect 29276 23672 29328 23724
rect 29368 23672 29420 23724
rect 29736 23715 29788 23724
rect 29736 23681 29745 23715
rect 29745 23681 29779 23715
rect 29779 23681 29788 23715
rect 29736 23672 29788 23681
rect 30656 23740 30708 23792
rect 32220 23740 32272 23792
rect 33876 23851 33928 23860
rect 33876 23817 33891 23851
rect 33891 23817 33925 23851
rect 33925 23817 33928 23851
rect 33876 23808 33928 23817
rect 34152 23740 34204 23792
rect 34612 23740 34664 23792
rect 30564 23672 30616 23724
rect 31024 23715 31076 23724
rect 31024 23681 31033 23715
rect 31033 23681 31067 23715
rect 31067 23681 31076 23715
rect 31024 23672 31076 23681
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 31576 23672 31628 23681
rect 31760 23672 31812 23724
rect 27896 23536 27948 23588
rect 28080 23536 28132 23588
rect 28908 23604 28960 23656
rect 29552 23647 29604 23656
rect 29552 23613 29561 23647
rect 29561 23613 29595 23647
rect 29595 23613 29604 23647
rect 29552 23604 29604 23613
rect 31116 23604 31168 23656
rect 32312 23604 32364 23656
rect 33048 23715 33100 23724
rect 33048 23681 33057 23715
rect 33057 23681 33091 23715
rect 33091 23681 33100 23715
rect 33048 23672 33100 23681
rect 33508 23672 33560 23724
rect 33600 23672 33652 23724
rect 34520 23672 34572 23724
rect 34796 23672 34848 23724
rect 34704 23604 34756 23656
rect 35348 23715 35400 23724
rect 35348 23681 35362 23715
rect 35362 23681 35396 23715
rect 35396 23681 35400 23715
rect 35348 23672 35400 23681
rect 37832 23808 37884 23860
rect 35992 23715 36044 23724
rect 35992 23681 36001 23715
rect 36001 23681 36035 23715
rect 36035 23681 36044 23715
rect 35992 23672 36044 23681
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 38200 23672 38252 23724
rect 38108 23647 38160 23656
rect 38108 23613 38117 23647
rect 38117 23613 38151 23647
rect 38151 23613 38160 23647
rect 38108 23604 38160 23613
rect 25504 23468 25556 23520
rect 28448 23511 28500 23520
rect 28448 23477 28457 23511
rect 28457 23477 28491 23511
rect 28491 23477 28500 23511
rect 28448 23468 28500 23477
rect 28540 23468 28592 23520
rect 28908 23468 28960 23520
rect 29368 23468 29420 23520
rect 31484 23468 31536 23520
rect 35808 23536 35860 23588
rect 32772 23468 32824 23520
rect 33600 23468 33652 23520
rect 35624 23468 35676 23520
rect 35900 23468 35952 23520
rect 37096 23468 37148 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3976 23307 4028 23316
rect 3976 23273 3985 23307
rect 3985 23273 4019 23307
rect 4019 23273 4028 23307
rect 3976 23264 4028 23273
rect 5172 23307 5224 23316
rect 5172 23273 5181 23307
rect 5181 23273 5215 23307
rect 5215 23273 5224 23307
rect 5172 23264 5224 23273
rect 5632 23264 5684 23316
rect 3884 23196 3936 23248
rect 5080 23128 5132 23180
rect 4620 23060 4672 23112
rect 6644 23196 6696 23248
rect 5724 23060 5776 23112
rect 6460 23060 6512 23112
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 9956 23060 10008 23112
rect 4896 22992 4948 23044
rect 6276 22992 6328 23044
rect 7472 22924 7524 22976
rect 10324 23035 10376 23044
rect 10324 23001 10333 23035
rect 10333 23001 10367 23035
rect 10367 23001 10376 23035
rect 10324 22992 10376 23001
rect 22284 23264 22336 23316
rect 22836 23264 22888 23316
rect 26240 23307 26292 23316
rect 26240 23273 26249 23307
rect 26249 23273 26283 23307
rect 26283 23273 26292 23307
rect 26240 23264 26292 23273
rect 36268 23264 36320 23316
rect 38200 23307 38252 23316
rect 38200 23273 38209 23307
rect 38209 23273 38243 23307
rect 38243 23273 38252 23307
rect 38200 23264 38252 23273
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 12348 23060 12400 23112
rect 14648 23196 14700 23248
rect 24676 23196 24728 23248
rect 26884 23196 26936 23248
rect 30104 23196 30156 23248
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 19984 23128 20036 23180
rect 20260 23128 20312 23180
rect 20444 23171 20496 23180
rect 20444 23137 20453 23171
rect 20453 23137 20487 23171
rect 20487 23137 20496 23171
rect 20444 23128 20496 23137
rect 20628 23128 20680 23180
rect 14556 23060 14608 23112
rect 14832 22992 14884 23044
rect 15200 23103 15252 23112
rect 15200 23069 15209 23103
rect 15209 23069 15243 23103
rect 15243 23069 15252 23103
rect 15200 23060 15252 23069
rect 15936 23060 15988 23112
rect 20904 23060 20956 23112
rect 29000 23128 29052 23180
rect 29184 23128 29236 23180
rect 24308 23060 24360 23112
rect 24952 23060 25004 23112
rect 25412 23060 25464 23112
rect 26976 23060 27028 23112
rect 27620 23060 27672 23112
rect 28816 23060 28868 23112
rect 29552 23128 29604 23180
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 34704 23128 34756 23180
rect 30564 23103 30616 23112
rect 30564 23069 30573 23103
rect 30573 23069 30607 23103
rect 30607 23069 30616 23103
rect 30564 23060 30616 23069
rect 33048 23060 33100 23112
rect 15292 22924 15344 22976
rect 18512 22924 18564 22976
rect 20076 22924 20128 22976
rect 20536 22992 20588 23044
rect 21364 22924 21416 22976
rect 21456 22967 21508 22976
rect 21456 22933 21465 22967
rect 21465 22933 21499 22967
rect 21499 22933 21508 22967
rect 21456 22924 21508 22933
rect 22192 22992 22244 23044
rect 25228 22992 25280 23044
rect 28632 22992 28684 23044
rect 30288 22992 30340 23044
rect 34520 22992 34572 23044
rect 36728 23060 36780 23112
rect 37096 23103 37148 23112
rect 37096 23069 37130 23103
rect 37130 23069 37148 23103
rect 37096 23060 37148 23069
rect 22652 22924 22704 22976
rect 25320 22924 25372 22976
rect 25596 22924 25648 22976
rect 27896 22924 27948 22976
rect 29092 22924 29144 22976
rect 30564 22924 30616 22976
rect 35624 22924 35676 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 5816 22763 5868 22772
rect 5816 22729 5825 22763
rect 5825 22729 5859 22763
rect 5859 22729 5868 22763
rect 5816 22720 5868 22729
rect 8300 22720 8352 22772
rect 10140 22720 10192 22772
rect 10324 22720 10376 22772
rect 11060 22720 11112 22772
rect 19984 22720 20036 22772
rect 20076 22763 20128 22772
rect 20076 22729 20085 22763
rect 20085 22729 20119 22763
rect 20119 22729 20128 22763
rect 20076 22720 20128 22729
rect 20168 22720 20220 22772
rect 20444 22720 20496 22772
rect 20536 22763 20588 22772
rect 20536 22729 20545 22763
rect 20545 22729 20579 22763
rect 20579 22729 20588 22763
rect 20536 22720 20588 22729
rect 4988 22652 5040 22704
rect 5632 22584 5684 22636
rect 6000 22584 6052 22636
rect 7196 22584 7248 22636
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 7564 22584 7616 22593
rect 7748 22695 7800 22704
rect 7748 22661 7757 22695
rect 7757 22661 7791 22695
rect 7791 22661 7800 22695
rect 7748 22652 7800 22661
rect 8760 22652 8812 22704
rect 11980 22695 12032 22704
rect 11980 22661 12014 22695
rect 12014 22661 12032 22695
rect 11980 22652 12032 22661
rect 14832 22652 14884 22704
rect 22284 22720 22336 22772
rect 24584 22763 24636 22772
rect 24584 22729 24593 22763
rect 24593 22729 24627 22763
rect 24627 22729 24636 22763
rect 24584 22720 24636 22729
rect 24768 22720 24820 22772
rect 27344 22720 27396 22772
rect 27436 22720 27488 22772
rect 32588 22720 32640 22772
rect 8208 22584 8260 22636
rect 12348 22584 12400 22636
rect 14464 22627 14516 22636
rect 14464 22593 14473 22627
rect 14473 22593 14507 22627
rect 14507 22593 14516 22627
rect 14464 22584 14516 22593
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 15200 22627 15252 22636
rect 15200 22593 15209 22627
rect 15209 22593 15243 22627
rect 15243 22593 15252 22627
rect 15200 22584 15252 22593
rect 14188 22516 14240 22568
rect 8300 22491 8352 22500
rect 8300 22457 8309 22491
rect 8309 22457 8343 22491
rect 8343 22457 8352 22491
rect 8300 22448 8352 22457
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 15568 22627 15620 22636
rect 15568 22593 15577 22627
rect 15577 22593 15611 22627
rect 15611 22593 15620 22627
rect 15568 22584 15620 22593
rect 15660 22584 15712 22636
rect 17224 22584 17276 22636
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 16672 22516 16724 22568
rect 16856 22448 16908 22500
rect 7012 22380 7064 22432
rect 7472 22423 7524 22432
rect 7472 22389 7481 22423
rect 7481 22389 7515 22423
rect 7515 22389 7524 22423
rect 7472 22380 7524 22389
rect 15384 22380 15436 22432
rect 15936 22380 15988 22432
rect 20168 22627 20220 22636
rect 20168 22593 20177 22627
rect 20177 22593 20211 22627
rect 20211 22593 20220 22627
rect 20168 22584 20220 22593
rect 22100 22584 22152 22636
rect 22468 22627 22520 22636
rect 22468 22593 22477 22627
rect 22477 22593 22511 22627
rect 22511 22593 22520 22627
rect 22468 22584 22520 22593
rect 22744 22584 22796 22636
rect 24492 22627 24544 22636
rect 24492 22593 24501 22627
rect 24501 22593 24535 22627
rect 24535 22593 24544 22627
rect 24492 22584 24544 22593
rect 24676 22627 24728 22636
rect 24676 22593 24685 22627
rect 24685 22593 24719 22627
rect 24719 22593 24728 22627
rect 24676 22584 24728 22593
rect 25688 22627 25740 22636
rect 25688 22593 25697 22627
rect 25697 22593 25731 22627
rect 25731 22593 25740 22627
rect 25688 22584 25740 22593
rect 26240 22652 26292 22704
rect 27988 22695 28040 22704
rect 27988 22661 27997 22695
rect 27997 22661 28031 22695
rect 28031 22661 28040 22695
rect 27988 22652 28040 22661
rect 26148 22627 26200 22636
rect 26148 22593 26157 22627
rect 26157 22593 26191 22627
rect 26191 22593 26200 22627
rect 26148 22584 26200 22593
rect 26516 22584 26568 22636
rect 20720 22516 20772 22568
rect 24768 22516 24820 22568
rect 26240 22516 26292 22568
rect 21824 22380 21876 22432
rect 22008 22380 22060 22432
rect 26424 22448 26476 22500
rect 27620 22584 27672 22636
rect 30012 22652 30064 22704
rect 27712 22516 27764 22568
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 31116 22652 31168 22704
rect 33600 22652 33652 22704
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 31116 22559 31168 22568
rect 31116 22525 31125 22559
rect 31125 22525 31159 22559
rect 31159 22525 31168 22559
rect 31116 22516 31168 22525
rect 31576 22627 31628 22636
rect 31576 22593 31585 22627
rect 31585 22593 31619 22627
rect 31619 22593 31628 22627
rect 31576 22584 31628 22593
rect 33508 22584 33560 22636
rect 37740 22584 37792 22636
rect 32496 22516 32548 22568
rect 33692 22516 33744 22568
rect 39028 22516 39080 22568
rect 31760 22448 31812 22500
rect 32312 22448 32364 22500
rect 33048 22448 33100 22500
rect 25044 22380 25096 22432
rect 25872 22380 25924 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 7196 22219 7248 22228
rect 7196 22185 7205 22219
rect 7205 22185 7239 22219
rect 7239 22185 7248 22219
rect 7196 22176 7248 22185
rect 6828 22108 6880 22160
rect 15476 22176 15528 22228
rect 20444 22176 20496 22228
rect 20628 22176 20680 22228
rect 25136 22176 25188 22228
rect 27712 22176 27764 22228
rect 28356 22176 28408 22228
rect 31852 22176 31904 22228
rect 32588 22176 32640 22228
rect 35716 22176 35768 22228
rect 14004 22108 14056 22160
rect 14556 22108 14608 22160
rect 15568 22108 15620 22160
rect 23940 22108 23992 22160
rect 27160 22108 27212 22160
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 4804 21972 4856 22024
rect 6644 22040 6696 22092
rect 6736 22040 6788 22092
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 5632 21904 5684 21956
rect 7656 22015 7708 22024
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 8300 22040 8352 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 9128 21972 9180 22024
rect 16856 22040 16908 22092
rect 17132 22040 17184 22092
rect 23020 22083 23072 22092
rect 23020 22049 23029 22083
rect 23029 22049 23063 22083
rect 23063 22049 23072 22083
rect 23020 22040 23072 22049
rect 25320 22040 25372 22092
rect 15016 22015 15068 22024
rect 15016 21981 15025 22015
rect 15025 21981 15059 22015
rect 15059 21981 15068 22015
rect 15016 21972 15068 21981
rect 15660 21972 15712 22024
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 19432 21972 19484 22024
rect 21456 21972 21508 22024
rect 22560 21972 22612 22024
rect 26792 22040 26844 22092
rect 23572 21972 23624 22024
rect 25228 22015 25280 22024
rect 25228 21981 25237 22015
rect 25237 21981 25271 22015
rect 25271 21981 25280 22015
rect 25228 21972 25280 21981
rect 25872 22015 25924 22024
rect 25872 21981 25881 22015
rect 25881 21981 25915 22015
rect 25915 21981 25924 22015
rect 25872 21972 25924 21981
rect 26148 21972 26200 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 28724 22108 28776 22160
rect 29276 22108 29328 22160
rect 29920 22108 29972 22160
rect 27988 22015 28040 22024
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 27988 21972 28040 21981
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 3976 21879 4028 21888
rect 3976 21845 3985 21879
rect 3985 21845 4019 21879
rect 4019 21845 4028 21879
rect 3976 21836 4028 21845
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 4344 21836 4396 21845
rect 6552 21836 6604 21888
rect 8116 21904 8168 21956
rect 9956 21904 10008 21956
rect 15568 21904 15620 21956
rect 23296 21904 23348 21956
rect 27620 21904 27672 21956
rect 28080 21904 28132 21956
rect 28724 21972 28776 22024
rect 29092 21972 29144 22024
rect 29184 21972 29236 22024
rect 30472 22040 30524 22092
rect 30380 21972 30432 22024
rect 10876 21836 10928 21888
rect 10968 21879 11020 21888
rect 10968 21845 10977 21879
rect 10977 21845 11011 21879
rect 11011 21845 11020 21879
rect 10968 21836 11020 21845
rect 14648 21836 14700 21888
rect 15752 21836 15804 21888
rect 16396 21836 16448 21888
rect 20168 21836 20220 21888
rect 25044 21836 25096 21888
rect 25688 21836 25740 21888
rect 26792 21879 26844 21888
rect 26792 21845 26801 21879
rect 26801 21845 26835 21879
rect 26835 21845 26844 21879
rect 26792 21836 26844 21845
rect 27068 21836 27120 21888
rect 29368 21836 29420 21888
rect 29644 21836 29696 21888
rect 30196 21904 30248 21956
rect 33232 22040 33284 22092
rect 33600 22083 33652 22092
rect 33600 22049 33609 22083
rect 33609 22049 33643 22083
rect 33643 22049 33652 22083
rect 33600 22040 33652 22049
rect 34060 22083 34112 22092
rect 34060 22049 34069 22083
rect 34069 22049 34103 22083
rect 34103 22049 34112 22083
rect 34060 22040 34112 22049
rect 35716 22040 35768 22092
rect 30932 21972 30984 22024
rect 31208 21972 31260 22024
rect 31484 22015 31536 22024
rect 31484 21981 31493 22015
rect 31493 21981 31527 22015
rect 31527 21981 31536 22015
rect 31484 21972 31536 21981
rect 32496 21972 32548 22024
rect 32864 21972 32916 22024
rect 32680 21947 32732 21956
rect 32680 21913 32689 21947
rect 32689 21913 32723 21947
rect 32723 21913 32732 21947
rect 32680 21904 32732 21913
rect 33048 22015 33100 22024
rect 33048 21981 33057 22015
rect 33057 21981 33091 22015
rect 33091 21981 33100 22015
rect 33048 21972 33100 21981
rect 33508 21972 33560 22024
rect 35532 22015 35584 22024
rect 35532 21981 35541 22015
rect 35541 21981 35575 22015
rect 35575 21981 35584 22015
rect 35532 21972 35584 21981
rect 35808 22015 35860 22024
rect 35808 21981 35817 22015
rect 35817 21981 35851 22015
rect 35851 21981 35860 22015
rect 35808 21972 35860 21981
rect 36268 21972 36320 22024
rect 36728 21972 36780 22024
rect 35992 21904 36044 21956
rect 37464 21904 37516 21956
rect 31392 21836 31444 21888
rect 32404 21879 32456 21888
rect 32404 21845 32413 21879
rect 32413 21845 32447 21879
rect 32447 21845 32456 21879
rect 32404 21836 32456 21845
rect 35900 21836 35952 21888
rect 37740 21836 37792 21888
rect 37924 21836 37976 21888
rect 38200 21879 38252 21888
rect 38200 21845 38209 21879
rect 38209 21845 38243 21879
rect 38243 21845 38252 21879
rect 38200 21836 38252 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4344 21632 4396 21684
rect 3976 21564 4028 21616
rect 6644 21564 6696 21616
rect 7656 21564 7708 21616
rect 5724 21496 5776 21548
rect 6184 21496 6236 21548
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 6828 21539 6880 21548
rect 6828 21505 6837 21539
rect 6837 21505 6871 21539
rect 6871 21505 6880 21539
rect 6828 21496 6880 21505
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7012 21496 7064 21548
rect 8300 21564 8352 21616
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 4620 21428 4672 21480
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 9496 21496 9548 21548
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 15384 21632 15436 21684
rect 10968 21564 11020 21616
rect 10140 21539 10192 21548
rect 10140 21505 10149 21539
rect 10149 21505 10183 21539
rect 10183 21505 10192 21539
rect 10140 21496 10192 21505
rect 10508 21496 10560 21548
rect 8116 21428 8168 21437
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 11060 21496 11112 21548
rect 14464 21539 14516 21548
rect 14464 21505 14473 21539
rect 14473 21505 14507 21539
rect 14507 21505 14516 21539
rect 14464 21496 14516 21505
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 16304 21564 16356 21616
rect 17592 21607 17644 21616
rect 17592 21573 17601 21607
rect 17601 21573 17635 21607
rect 17635 21573 17644 21607
rect 17592 21564 17644 21573
rect 18880 21675 18932 21684
rect 18880 21641 18889 21675
rect 18889 21641 18923 21675
rect 18923 21641 18932 21675
rect 18880 21632 18932 21641
rect 22744 21632 22796 21684
rect 19984 21564 20036 21616
rect 24860 21632 24912 21684
rect 26424 21632 26476 21684
rect 27252 21632 27304 21684
rect 16396 21496 16448 21548
rect 18052 21496 18104 21548
rect 19156 21496 19208 21548
rect 27528 21564 27580 21616
rect 25596 21496 25648 21548
rect 26608 21496 26660 21548
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 28540 21632 28592 21684
rect 28816 21632 28868 21684
rect 29644 21632 29696 21684
rect 29828 21632 29880 21684
rect 29920 21632 29972 21684
rect 35532 21632 35584 21684
rect 36268 21675 36320 21684
rect 36268 21641 36277 21675
rect 36277 21641 36311 21675
rect 36311 21641 36320 21675
rect 36268 21632 36320 21641
rect 37464 21675 37516 21684
rect 37464 21641 37473 21675
rect 37473 21641 37507 21675
rect 37507 21641 37516 21675
rect 37464 21632 37516 21641
rect 37924 21675 37976 21684
rect 37924 21641 37933 21675
rect 37933 21641 37967 21675
rect 37967 21641 37976 21675
rect 37924 21632 37976 21641
rect 28448 21564 28500 21616
rect 30104 21564 30156 21616
rect 30564 21564 30616 21616
rect 31208 21564 31260 21616
rect 32404 21564 32456 21616
rect 34060 21564 34112 21616
rect 34612 21564 34664 21616
rect 35992 21607 36044 21616
rect 35992 21573 36001 21607
rect 36001 21573 36035 21607
rect 36035 21573 36044 21607
rect 35992 21564 36044 21573
rect 38200 21564 38252 21616
rect 16028 21428 16080 21480
rect 15936 21360 15988 21412
rect 16304 21471 16356 21480
rect 16304 21437 16313 21471
rect 16313 21437 16347 21471
rect 16347 21437 16356 21471
rect 16304 21428 16356 21437
rect 16948 21428 17000 21480
rect 24492 21471 24544 21480
rect 24492 21437 24501 21471
rect 24501 21437 24535 21471
rect 24535 21437 24544 21471
rect 24492 21428 24544 21437
rect 16580 21360 16632 21412
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 10324 21292 10376 21344
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 23572 21292 23624 21344
rect 24860 21428 24912 21480
rect 27068 21428 27120 21480
rect 27528 21428 27580 21480
rect 27896 21428 27948 21480
rect 25044 21360 25096 21412
rect 24676 21292 24728 21344
rect 24768 21292 24820 21344
rect 25780 21292 25832 21344
rect 27620 21292 27672 21344
rect 27988 21360 28040 21412
rect 29368 21360 29420 21412
rect 29828 21539 29880 21548
rect 29828 21505 29837 21539
rect 29837 21505 29871 21539
rect 29871 21505 29880 21539
rect 29828 21496 29880 21505
rect 31484 21496 31536 21548
rect 32772 21496 32824 21548
rect 34796 21496 34848 21548
rect 30012 21428 30064 21480
rect 30196 21471 30248 21480
rect 30196 21437 30205 21471
rect 30205 21437 30239 21471
rect 30239 21437 30248 21471
rect 30196 21428 30248 21437
rect 30932 21360 30984 21412
rect 32036 21428 32088 21480
rect 33692 21471 33744 21480
rect 33692 21437 33701 21471
rect 33701 21437 33735 21471
rect 33735 21437 33744 21471
rect 33692 21428 33744 21437
rect 33600 21360 33652 21412
rect 28448 21292 28500 21344
rect 28540 21335 28592 21344
rect 28540 21301 28549 21335
rect 28549 21301 28583 21335
rect 28583 21301 28592 21335
rect 28540 21292 28592 21301
rect 30748 21292 30800 21344
rect 35440 21428 35492 21480
rect 35348 21360 35400 21412
rect 38016 21471 38068 21480
rect 38016 21437 38025 21471
rect 38025 21437 38059 21471
rect 38059 21437 38068 21471
rect 38016 21428 38068 21437
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6828 21088 6880 21140
rect 7656 21088 7708 21140
rect 3056 20884 3108 20936
rect 5448 20884 5500 20936
rect 10324 20927 10376 20936
rect 10324 20893 10333 20927
rect 10333 20893 10367 20927
rect 10367 20893 10376 20927
rect 10324 20884 10376 20893
rect 15200 21088 15252 21140
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 11060 20952 11112 21004
rect 7104 20816 7156 20868
rect 9496 20859 9548 20868
rect 9496 20825 9505 20859
rect 9505 20825 9539 20859
rect 9539 20825 9548 20859
rect 9496 20816 9548 20825
rect 11152 20884 11204 20936
rect 11428 20884 11480 20936
rect 14280 21020 14332 21072
rect 26700 21088 26752 21140
rect 27436 21088 27488 21140
rect 21548 21020 21600 21072
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 15844 20884 15896 20936
rect 14464 20816 14516 20868
rect 14648 20859 14700 20868
rect 14648 20825 14657 20859
rect 14657 20825 14691 20859
rect 14691 20825 14700 20859
rect 14648 20816 14700 20825
rect 11060 20748 11112 20800
rect 12072 20748 12124 20800
rect 13820 20748 13872 20800
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 16580 20952 16632 21004
rect 22008 20952 22060 21004
rect 22192 20952 22244 21004
rect 22284 20952 22336 21004
rect 22468 20952 22520 21004
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 17040 20816 17092 20868
rect 22100 20816 22152 20868
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 26148 20995 26200 21004
rect 26148 20961 26157 20995
rect 26157 20961 26191 20995
rect 26191 20961 26200 20995
rect 26148 20952 26200 20961
rect 22928 20859 22980 20868
rect 22928 20825 22954 20859
rect 22954 20825 22980 20859
rect 22928 20816 22980 20825
rect 24492 20884 24544 20936
rect 24952 20884 25004 20936
rect 25044 20927 25096 20936
rect 25044 20893 25053 20927
rect 25053 20893 25087 20927
rect 25087 20893 25096 20927
rect 25044 20884 25096 20893
rect 26424 20927 26476 20936
rect 26424 20893 26433 20927
rect 26433 20893 26467 20927
rect 26467 20893 26476 20927
rect 26424 20884 26476 20893
rect 29644 21088 29696 21140
rect 31300 21131 31352 21140
rect 27712 21020 27764 21072
rect 31300 21097 31324 21131
rect 31324 21097 31352 21131
rect 31300 21088 31352 21097
rect 31392 21063 31444 21072
rect 31392 21029 31401 21063
rect 31401 21029 31435 21063
rect 31435 21029 31444 21063
rect 31392 21020 31444 21029
rect 32588 21088 32640 21140
rect 35808 21088 35860 21140
rect 31852 21020 31904 21072
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 27712 20927 27764 20936
rect 27712 20893 27722 20927
rect 27722 20893 27756 20927
rect 27756 20893 27764 20927
rect 29368 20952 29420 21004
rect 29552 20952 29604 21004
rect 27712 20884 27764 20893
rect 27988 20927 28040 20936
rect 27988 20893 27997 20927
rect 27997 20893 28031 20927
rect 28031 20893 28040 20927
rect 27988 20884 28040 20893
rect 28080 20927 28132 20936
rect 28080 20893 28094 20927
rect 28094 20893 28128 20927
rect 28128 20893 28132 20927
rect 28080 20884 28132 20893
rect 28356 20884 28408 20936
rect 29460 20884 29512 20936
rect 30656 20952 30708 21004
rect 30840 20952 30892 21004
rect 31576 20952 31628 21004
rect 34520 20952 34572 21004
rect 35900 21020 35952 21072
rect 34704 20884 34756 20936
rect 35624 20884 35676 20936
rect 16028 20748 16080 20800
rect 17592 20748 17644 20800
rect 23112 20748 23164 20800
rect 24860 20748 24912 20800
rect 26884 20748 26936 20800
rect 31484 20816 31536 20868
rect 35716 20816 35768 20868
rect 37740 20884 37792 20936
rect 39028 20816 39080 20868
rect 29368 20748 29420 20800
rect 29828 20748 29880 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6828 20544 6880 20596
rect 5540 20476 5592 20528
rect 9128 20476 9180 20528
rect 13820 20476 13872 20528
rect 14464 20544 14516 20596
rect 14740 20544 14792 20596
rect 15568 20544 15620 20596
rect 19708 20544 19760 20596
rect 19984 20544 20036 20596
rect 16672 20476 16724 20528
rect 7104 20408 7156 20460
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 17592 20408 17644 20460
rect 19248 20476 19300 20528
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 19524 20408 19576 20460
rect 20076 20476 20128 20528
rect 22560 20476 22612 20528
rect 23112 20476 23164 20528
rect 11520 20340 11572 20392
rect 15384 20383 15436 20392
rect 15384 20349 15393 20383
rect 15393 20349 15427 20383
rect 15427 20349 15436 20383
rect 15384 20340 15436 20349
rect 15568 20383 15620 20392
rect 15568 20349 15577 20383
rect 15577 20349 15611 20383
rect 15611 20349 15620 20383
rect 15568 20340 15620 20349
rect 16304 20340 16356 20392
rect 18328 20383 18380 20392
rect 18328 20349 18337 20383
rect 18337 20349 18371 20383
rect 18371 20349 18380 20383
rect 18328 20340 18380 20349
rect 15936 20272 15988 20324
rect 19248 20272 19300 20324
rect 16948 20204 17000 20256
rect 19708 20204 19760 20256
rect 19800 20204 19852 20256
rect 20352 20204 20404 20256
rect 22744 20408 22796 20460
rect 24584 20451 24636 20460
rect 24584 20417 24593 20451
rect 24593 20417 24627 20451
rect 24627 20417 24636 20451
rect 24584 20408 24636 20417
rect 25044 20408 25096 20460
rect 25596 20451 25648 20460
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 20996 20340 21048 20392
rect 20720 20272 20772 20324
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 24860 20340 24912 20392
rect 27344 20544 27396 20596
rect 27712 20544 27764 20596
rect 29000 20544 29052 20596
rect 33508 20587 33560 20596
rect 33508 20553 33517 20587
rect 33517 20553 33551 20587
rect 33551 20553 33560 20587
rect 33508 20544 33560 20553
rect 28172 20476 28224 20528
rect 31668 20476 31720 20528
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27620 20408 27672 20460
rect 28724 20408 28776 20460
rect 29000 20408 29052 20460
rect 27896 20340 27948 20392
rect 29736 20340 29788 20392
rect 30656 20451 30708 20460
rect 30656 20417 30665 20451
rect 30665 20417 30699 20451
rect 30699 20417 30708 20451
rect 30656 20408 30708 20417
rect 30748 20451 30800 20460
rect 30748 20417 30757 20451
rect 30757 20417 30791 20451
rect 30791 20417 30800 20451
rect 30748 20408 30800 20417
rect 30932 20408 30984 20460
rect 32680 20340 32732 20392
rect 33232 20408 33284 20460
rect 37740 20476 37792 20528
rect 35440 20408 35492 20460
rect 33508 20340 33560 20392
rect 33968 20340 34020 20392
rect 35624 20451 35676 20460
rect 35624 20417 35633 20451
rect 35633 20417 35667 20451
rect 35667 20417 35676 20451
rect 35624 20408 35676 20417
rect 37832 20451 37884 20460
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 38016 20383 38068 20392
rect 38016 20349 38025 20383
rect 38025 20349 38059 20383
rect 38059 20349 38068 20383
rect 38016 20340 38068 20349
rect 24952 20272 25004 20324
rect 31392 20272 31444 20324
rect 27436 20204 27488 20256
rect 29828 20204 29880 20256
rect 30748 20204 30800 20256
rect 31576 20204 31628 20256
rect 35808 20204 35860 20256
rect 37464 20247 37516 20256
rect 37464 20213 37473 20247
rect 37473 20213 37507 20247
rect 37507 20213 37516 20247
rect 37464 20204 37516 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7104 20043 7156 20052
rect 7104 20009 7113 20043
rect 7113 20009 7147 20043
rect 7147 20009 7156 20043
rect 7104 20000 7156 20009
rect 5632 19932 5684 19984
rect 15384 20000 15436 20052
rect 16672 20000 16724 20052
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 19524 20000 19576 20052
rect 17408 19932 17460 19984
rect 4620 19907 4672 19916
rect 4620 19873 4629 19907
rect 4629 19873 4663 19907
rect 4663 19873 4672 19907
rect 4620 19864 4672 19873
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 16028 19864 16080 19916
rect 16396 19864 16448 19916
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 4712 19796 4764 19848
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 6920 19839 6972 19848
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 8944 19796 8996 19848
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 14556 19796 14608 19848
rect 15660 19796 15712 19848
rect 6736 19771 6788 19780
rect 6736 19737 6745 19771
rect 6745 19737 6779 19771
rect 6779 19737 6788 19771
rect 6736 19728 6788 19737
rect 9220 19728 9272 19780
rect 10968 19728 11020 19780
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 4436 19703 4488 19712
rect 4436 19669 4445 19703
rect 4445 19669 4479 19703
rect 4479 19669 4488 19703
rect 4436 19660 4488 19669
rect 6828 19660 6880 19712
rect 7932 19660 7984 19712
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 14832 19728 14884 19780
rect 17500 19796 17552 19848
rect 20996 19932 21048 19984
rect 21456 19975 21508 19984
rect 21456 19941 21465 19975
rect 21465 19941 21499 19975
rect 21499 19941 21508 19975
rect 21456 19932 21508 19941
rect 17684 19864 17736 19916
rect 19708 19864 19760 19916
rect 22008 20000 22060 20052
rect 22468 20000 22520 20052
rect 24768 20000 24820 20052
rect 25044 20043 25096 20052
rect 25044 20009 25053 20043
rect 25053 20009 25087 20043
rect 25087 20009 25096 20043
rect 25044 20000 25096 20009
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 28632 20000 28684 20052
rect 29828 20043 29880 20052
rect 29828 20009 29837 20043
rect 29837 20009 29871 20043
rect 29871 20009 29880 20043
rect 29828 20000 29880 20009
rect 34612 20000 34664 20052
rect 35164 20000 35216 20052
rect 35624 20000 35676 20052
rect 15936 19728 15988 19780
rect 17132 19771 17184 19780
rect 17132 19737 17141 19771
rect 17141 19737 17175 19771
rect 17175 19737 17184 19771
rect 17132 19728 17184 19737
rect 20720 19796 20772 19848
rect 21640 19839 21692 19848
rect 21640 19805 21644 19839
rect 21644 19805 21678 19839
rect 21678 19805 21692 19839
rect 21640 19796 21692 19805
rect 23204 19907 23256 19916
rect 23204 19873 23213 19907
rect 23213 19873 23247 19907
rect 23247 19873 23256 19907
rect 23204 19864 23256 19873
rect 24676 19907 24728 19916
rect 24676 19873 24685 19907
rect 24685 19873 24719 19907
rect 24719 19873 24728 19907
rect 24676 19864 24728 19873
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 10508 19660 10560 19669
rect 14740 19660 14792 19712
rect 15568 19660 15620 19712
rect 16396 19660 16448 19712
rect 17316 19660 17368 19712
rect 17408 19660 17460 19712
rect 18696 19660 18748 19712
rect 19984 19728 20036 19780
rect 21916 19728 21968 19780
rect 22284 19728 22336 19780
rect 20260 19660 20312 19712
rect 20628 19660 20680 19712
rect 22652 19796 22704 19848
rect 23388 19839 23440 19848
rect 23388 19805 23397 19839
rect 23397 19805 23431 19839
rect 23431 19805 23440 19839
rect 23388 19796 23440 19805
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 26240 19932 26292 19984
rect 26516 19864 26568 19916
rect 27620 19932 27672 19984
rect 27896 19932 27948 19984
rect 27068 19796 27120 19848
rect 23112 19660 23164 19712
rect 27160 19660 27212 19712
rect 28172 19796 28224 19848
rect 27988 19728 28040 19780
rect 31576 19932 31628 19984
rect 29092 19864 29144 19916
rect 30656 19864 30708 19916
rect 28724 19796 28776 19848
rect 28908 19839 28960 19848
rect 28908 19805 28917 19839
rect 28917 19805 28951 19839
rect 28951 19805 28960 19839
rect 28908 19796 28960 19805
rect 29000 19839 29052 19848
rect 29000 19805 29014 19839
rect 29014 19805 29048 19839
rect 29048 19805 29052 19839
rect 29000 19796 29052 19805
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 29828 19839 29880 19848
rect 29828 19805 29837 19839
rect 29837 19805 29871 19839
rect 29871 19805 29880 19839
rect 29828 19796 29880 19805
rect 29920 19796 29972 19848
rect 32496 19864 32548 19916
rect 32220 19796 32272 19848
rect 32404 19839 32456 19848
rect 32404 19805 32414 19839
rect 32414 19805 32448 19839
rect 32448 19805 32456 19839
rect 32404 19796 32456 19805
rect 33508 19907 33560 19916
rect 33508 19873 33517 19907
rect 33517 19873 33551 19907
rect 33551 19873 33560 19907
rect 33508 19864 33560 19873
rect 34428 19864 34480 19916
rect 28540 19660 28592 19712
rect 28632 19660 28684 19712
rect 29184 19703 29236 19712
rect 29184 19669 29193 19703
rect 29193 19669 29227 19703
rect 29227 19669 29236 19703
rect 29184 19660 29236 19669
rect 29460 19660 29512 19712
rect 31024 19771 31076 19780
rect 31024 19737 31033 19771
rect 31033 19737 31067 19771
rect 31067 19737 31076 19771
rect 31024 19728 31076 19737
rect 32036 19728 32088 19780
rect 33232 19796 33284 19848
rect 34796 19796 34848 19848
rect 35072 19864 35124 19916
rect 35256 19839 35308 19848
rect 35256 19805 35265 19839
rect 35265 19805 35299 19839
rect 35299 19805 35308 19839
rect 35256 19796 35308 19805
rect 35348 19839 35400 19848
rect 35348 19805 35362 19839
rect 35362 19805 35396 19839
rect 35396 19805 35400 19839
rect 35348 19796 35400 19805
rect 36728 19839 36780 19848
rect 36728 19805 36737 19839
rect 36737 19805 36771 19839
rect 36771 19805 36780 19839
rect 36728 19796 36780 19805
rect 37464 19796 37516 19848
rect 29920 19660 29972 19712
rect 35164 19771 35216 19780
rect 35164 19737 35173 19771
rect 35173 19737 35207 19771
rect 35207 19737 35216 19771
rect 35164 19728 35216 19737
rect 32864 19660 32916 19712
rect 32956 19703 33008 19712
rect 32956 19669 32965 19703
rect 32965 19669 32999 19703
rect 32999 19669 33008 19703
rect 32956 19660 33008 19669
rect 37832 19660 37884 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5632 19499 5684 19508
rect 5632 19465 5641 19499
rect 5641 19465 5675 19499
rect 5675 19465 5684 19499
rect 5632 19456 5684 19465
rect 7564 19456 7616 19508
rect 9220 19456 9272 19508
rect 4068 19388 4120 19440
rect 7932 19388 7984 19440
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 4620 19320 4672 19372
rect 6644 19320 6696 19372
rect 8484 19320 8536 19372
rect 10508 19388 10560 19440
rect 9312 19363 9364 19372
rect 9312 19329 9321 19363
rect 9321 19329 9355 19363
rect 9355 19329 9364 19363
rect 9312 19320 9364 19329
rect 9680 19363 9732 19372
rect 9680 19329 9689 19363
rect 9689 19329 9723 19363
rect 9723 19329 9732 19363
rect 9680 19320 9732 19329
rect 10600 19363 10652 19372
rect 10600 19329 10609 19363
rect 10609 19329 10643 19363
rect 10643 19329 10652 19363
rect 10600 19320 10652 19329
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 4436 19184 4488 19236
rect 5448 19184 5500 19236
rect 15200 19456 15252 19508
rect 15568 19499 15620 19508
rect 15568 19465 15577 19499
rect 15577 19465 15611 19499
rect 15611 19465 15620 19499
rect 15568 19456 15620 19465
rect 17500 19456 17552 19508
rect 19248 19456 19300 19508
rect 15476 19388 15528 19440
rect 11520 19320 11572 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 14832 19184 14884 19236
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 17408 19363 17460 19372
rect 17408 19329 17417 19363
rect 17417 19329 17451 19363
rect 17451 19329 17460 19363
rect 17408 19320 17460 19329
rect 18236 19388 18288 19440
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 20168 19456 20220 19508
rect 21732 19388 21784 19440
rect 30932 19456 30984 19508
rect 33508 19456 33560 19508
rect 35440 19456 35492 19508
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 19340 19252 19392 19304
rect 20260 19320 20312 19372
rect 20536 19320 20588 19372
rect 21180 19320 21232 19372
rect 22284 19363 22336 19372
rect 22284 19329 22293 19363
rect 22293 19329 22327 19363
rect 22327 19329 22336 19363
rect 22284 19320 22336 19329
rect 27068 19388 27120 19440
rect 23020 19363 23072 19372
rect 23020 19329 23029 19363
rect 23029 19329 23063 19363
rect 23063 19329 23072 19363
rect 23020 19320 23072 19329
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 23296 19320 23348 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 24584 19363 24636 19372
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 28080 19388 28132 19440
rect 27988 19320 28040 19372
rect 29092 19388 29144 19440
rect 30196 19388 30248 19440
rect 31668 19388 31720 19440
rect 32956 19388 33008 19440
rect 33692 19388 33744 19440
rect 20996 19252 21048 19304
rect 25504 19252 25556 19304
rect 28356 19252 28408 19304
rect 28540 19252 28592 19304
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 6736 19116 6788 19168
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15200 19116 15252 19168
rect 15384 19116 15436 19168
rect 15844 19116 15896 19168
rect 16948 19116 17000 19168
rect 19064 19116 19116 19168
rect 24400 19184 24452 19236
rect 24492 19184 24544 19236
rect 27712 19184 27764 19236
rect 19984 19159 20036 19168
rect 19984 19125 19993 19159
rect 19993 19125 20027 19159
rect 20027 19125 20036 19159
rect 19984 19116 20036 19125
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 29460 19363 29512 19372
rect 29460 19329 29467 19363
rect 29467 19329 29512 19363
rect 29460 19320 29512 19329
rect 29644 19363 29696 19372
rect 29644 19329 29653 19363
rect 29653 19329 29687 19363
rect 29687 19329 29696 19363
rect 29644 19320 29696 19329
rect 29736 19363 29788 19372
rect 29736 19329 29750 19363
rect 29750 19329 29784 19363
rect 29784 19329 29788 19363
rect 29736 19320 29788 19329
rect 32680 19320 32732 19372
rect 33324 19363 33376 19372
rect 33324 19329 33333 19363
rect 33333 19329 33367 19363
rect 33367 19329 33376 19363
rect 33324 19320 33376 19329
rect 33508 19363 33560 19372
rect 33508 19329 33517 19363
rect 33517 19329 33551 19363
rect 33551 19329 33560 19363
rect 33508 19320 33560 19329
rect 36728 19388 36780 19440
rect 34428 19320 34480 19372
rect 37556 19320 37608 19372
rect 39028 19320 39080 19372
rect 29092 19252 29144 19304
rect 31852 19252 31904 19304
rect 29828 19184 29880 19236
rect 30104 19184 30156 19236
rect 34152 19184 34204 19236
rect 29184 19116 29236 19168
rect 29276 19116 29328 19168
rect 33600 19116 33652 19168
rect 35072 19116 35124 19168
rect 35440 19116 35492 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5632 18912 5684 18964
rect 13268 18912 13320 18964
rect 5448 18844 5500 18896
rect 15936 18912 15988 18964
rect 17132 18912 17184 18964
rect 19892 18912 19944 18964
rect 20076 18912 20128 18964
rect 20536 18912 20588 18964
rect 24584 18955 24636 18964
rect 24584 18921 24593 18955
rect 24593 18921 24627 18955
rect 24627 18921 24636 18955
rect 24584 18912 24636 18921
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 6920 18776 6972 18828
rect 3424 18708 3476 18760
rect 5632 18708 5684 18760
rect 6092 18708 6144 18760
rect 7380 18776 7432 18828
rect 13360 18776 13412 18828
rect 8668 18708 8720 18760
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 15200 18708 15252 18760
rect 5264 18640 5316 18692
rect 6552 18615 6604 18624
rect 6552 18581 6561 18615
rect 6561 18581 6595 18615
rect 6595 18581 6604 18615
rect 6552 18572 6604 18581
rect 6828 18572 6880 18624
rect 8576 18572 8628 18624
rect 9404 18683 9456 18692
rect 9404 18649 9413 18683
rect 9413 18649 9447 18683
rect 9447 18649 9456 18683
rect 9404 18640 9456 18649
rect 10324 18640 10376 18692
rect 19064 18844 19116 18896
rect 19156 18844 19208 18896
rect 19616 18844 19668 18896
rect 23296 18844 23348 18896
rect 32680 18912 32732 18964
rect 33508 18912 33560 18964
rect 36084 18844 36136 18896
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 30104 18776 30156 18828
rect 31024 18776 31076 18828
rect 31484 18776 31536 18828
rect 18328 18708 18380 18760
rect 16488 18640 16540 18692
rect 19892 18708 19944 18760
rect 20996 18708 21048 18760
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 22008 18708 22060 18760
rect 23572 18708 23624 18760
rect 24492 18708 24544 18760
rect 18972 18640 19024 18692
rect 24676 18640 24728 18692
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 26424 18751 26476 18760
rect 26424 18717 26433 18751
rect 26433 18717 26467 18751
rect 26467 18717 26476 18751
rect 26424 18708 26476 18717
rect 26516 18751 26568 18760
rect 26516 18717 26525 18751
rect 26525 18717 26559 18751
rect 26559 18717 26568 18751
rect 26516 18708 26568 18717
rect 27252 18640 27304 18692
rect 12716 18572 12768 18624
rect 13268 18572 13320 18624
rect 16764 18572 16816 18624
rect 20628 18572 20680 18624
rect 27896 18572 27948 18624
rect 27988 18615 28040 18624
rect 27988 18581 27997 18615
rect 27997 18581 28031 18615
rect 28031 18581 28040 18615
rect 27988 18572 28040 18581
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 31300 18751 31352 18760
rect 31300 18717 31309 18751
rect 31309 18717 31343 18751
rect 31343 18717 31352 18751
rect 31300 18708 31352 18717
rect 31852 18751 31904 18760
rect 31852 18717 31861 18751
rect 31861 18717 31895 18751
rect 31895 18717 31904 18751
rect 31852 18708 31904 18717
rect 32496 18776 32548 18828
rect 32220 18708 32272 18760
rect 28264 18683 28316 18692
rect 28264 18649 28273 18683
rect 28273 18649 28307 18683
rect 28307 18649 28316 18683
rect 28264 18640 28316 18649
rect 28724 18640 28776 18692
rect 29736 18640 29788 18692
rect 29000 18572 29052 18624
rect 32220 18572 32272 18624
rect 32680 18640 32732 18692
rect 33048 18751 33100 18760
rect 33048 18717 33057 18751
rect 33057 18717 33091 18751
rect 33091 18717 33100 18751
rect 33048 18708 33100 18717
rect 38016 18776 38068 18828
rect 33140 18683 33192 18692
rect 33140 18649 33149 18683
rect 33149 18649 33183 18683
rect 33183 18649 33192 18683
rect 35532 18708 35584 18760
rect 33140 18640 33192 18649
rect 38108 18640 38160 18692
rect 35348 18572 35400 18624
rect 37004 18572 37056 18624
rect 37556 18615 37608 18624
rect 37556 18581 37565 18615
rect 37565 18581 37599 18615
rect 37599 18581 37608 18615
rect 37556 18572 37608 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9312 18368 9364 18420
rect 9128 18300 9180 18352
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 8576 18275 8628 18284
rect 8576 18241 8610 18275
rect 8610 18241 8628 18275
rect 8576 18232 8628 18241
rect 10600 18300 10652 18352
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 10968 18368 11020 18420
rect 11704 18300 11756 18352
rect 12256 18300 12308 18352
rect 10600 18164 10652 18216
rect 9404 18096 9456 18148
rect 11244 18028 11296 18080
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 15844 18368 15896 18420
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 13452 18300 13504 18352
rect 16212 18300 16264 18352
rect 13360 18232 13412 18284
rect 13452 18207 13504 18216
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 14832 18232 14884 18284
rect 16764 18232 16816 18284
rect 20628 18300 20680 18352
rect 21272 18368 21324 18420
rect 22008 18411 22060 18420
rect 22008 18377 22017 18411
rect 22017 18377 22051 18411
rect 22051 18377 22060 18411
rect 22008 18368 22060 18377
rect 24860 18411 24912 18420
rect 24860 18377 24869 18411
rect 24869 18377 24903 18411
rect 24903 18377 24912 18411
rect 24860 18368 24912 18377
rect 28264 18368 28316 18420
rect 22836 18300 22888 18352
rect 20444 18232 20496 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 22100 18232 22152 18284
rect 22376 18232 22428 18284
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 23112 18232 23164 18284
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 23664 18300 23716 18352
rect 24676 18300 24728 18352
rect 27896 18300 27948 18352
rect 29552 18368 29604 18420
rect 33232 18411 33284 18420
rect 33232 18377 33241 18411
rect 33241 18377 33275 18411
rect 33275 18377 33284 18411
rect 33232 18368 33284 18377
rect 37556 18368 37608 18420
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 24768 18232 24820 18284
rect 17132 18164 17184 18216
rect 17592 18207 17644 18216
rect 17592 18173 17601 18207
rect 17601 18173 17635 18207
rect 17635 18173 17644 18207
rect 17592 18164 17644 18173
rect 19984 18164 20036 18216
rect 20260 18164 20312 18216
rect 21088 18207 21140 18216
rect 21088 18173 21097 18207
rect 21097 18173 21131 18207
rect 21131 18173 21140 18207
rect 21088 18164 21140 18173
rect 12900 18028 12952 18080
rect 14832 18096 14884 18148
rect 16028 18096 16080 18148
rect 24216 18207 24268 18216
rect 24216 18173 24225 18207
rect 24225 18173 24259 18207
rect 24259 18173 24268 18207
rect 24216 18164 24268 18173
rect 24860 18164 24912 18216
rect 25596 18275 25648 18284
rect 25596 18241 25605 18275
rect 25605 18241 25639 18275
rect 25639 18241 25648 18275
rect 25596 18232 25648 18241
rect 28908 18232 28960 18284
rect 27804 18164 27856 18216
rect 28356 18164 28408 18216
rect 29092 18164 29144 18216
rect 14648 18028 14700 18080
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 20444 18028 20496 18080
rect 21272 18028 21324 18080
rect 22836 18096 22888 18148
rect 28448 18096 28500 18148
rect 29276 18139 29328 18148
rect 29276 18105 29285 18139
rect 29285 18105 29319 18139
rect 29319 18105 29328 18139
rect 29276 18096 29328 18105
rect 33600 18343 33652 18352
rect 33600 18309 33609 18343
rect 33609 18309 33643 18343
rect 33643 18309 33652 18343
rect 33600 18300 33652 18309
rect 35256 18343 35308 18352
rect 35256 18309 35265 18343
rect 35265 18309 35299 18343
rect 35299 18309 35308 18343
rect 35256 18300 35308 18309
rect 35348 18343 35400 18352
rect 35348 18309 35357 18343
rect 35357 18309 35391 18343
rect 35391 18309 35400 18343
rect 35348 18300 35400 18309
rect 33508 18232 33560 18284
rect 34796 18232 34848 18284
rect 35072 18275 35124 18284
rect 35072 18241 35082 18275
rect 35082 18241 35116 18275
rect 35116 18241 35124 18275
rect 35072 18232 35124 18241
rect 35440 18275 35492 18284
rect 35440 18241 35454 18275
rect 35454 18241 35488 18275
rect 35488 18241 35492 18275
rect 35440 18232 35492 18241
rect 35900 18232 35952 18284
rect 36360 18275 36412 18284
rect 36360 18241 36369 18275
rect 36369 18241 36403 18275
rect 36403 18241 36412 18275
rect 36360 18232 36412 18241
rect 37832 18275 37884 18284
rect 37832 18241 37841 18275
rect 37841 18241 37875 18275
rect 37875 18241 37884 18275
rect 37832 18232 37884 18241
rect 35440 18096 35492 18148
rect 39028 18164 39080 18216
rect 24584 18028 24636 18080
rect 24952 18028 25004 18080
rect 25320 18071 25372 18080
rect 25320 18037 25329 18071
rect 25329 18037 25363 18071
rect 25363 18037 25372 18071
rect 25320 18028 25372 18037
rect 27620 18028 27672 18080
rect 30196 18028 30248 18080
rect 31668 18028 31720 18080
rect 33324 18028 33376 18080
rect 35808 18028 35860 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 7380 17867 7432 17876
rect 7380 17833 7389 17867
rect 7389 17833 7423 17867
rect 7423 17833 7432 17867
rect 7380 17824 7432 17833
rect 10600 17824 10652 17876
rect 17132 17867 17184 17876
rect 17132 17833 17141 17867
rect 17141 17833 17175 17867
rect 17175 17833 17184 17867
rect 17132 17824 17184 17833
rect 12256 17756 12308 17808
rect 12716 17731 12768 17740
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 5632 17620 5684 17672
rect 8300 17620 8352 17672
rect 11244 17663 11296 17672
rect 11244 17629 11262 17663
rect 11262 17629 11296 17663
rect 11244 17620 11296 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 17224 17756 17276 17808
rect 20076 17756 20128 17808
rect 24216 17824 24268 17876
rect 24308 17824 24360 17876
rect 22376 17756 22428 17808
rect 6552 17552 6604 17604
rect 13820 17552 13872 17604
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 14832 17620 14884 17672
rect 18604 17731 18656 17740
rect 18604 17697 18613 17731
rect 18613 17697 18647 17731
rect 18647 17697 18656 17731
rect 18604 17688 18656 17697
rect 18696 17731 18748 17740
rect 18696 17697 18705 17731
rect 18705 17697 18739 17731
rect 18739 17697 18748 17731
rect 18696 17688 18748 17697
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 17040 17620 17092 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 17500 17620 17552 17672
rect 17868 17620 17920 17672
rect 21640 17663 21692 17672
rect 21640 17629 21689 17663
rect 21689 17629 21692 17663
rect 21640 17620 21692 17629
rect 17132 17552 17184 17604
rect 18052 17552 18104 17604
rect 19248 17552 19300 17604
rect 21916 17595 21968 17604
rect 21916 17561 21925 17595
rect 21925 17561 21959 17595
rect 21959 17561 21968 17595
rect 21916 17552 21968 17561
rect 23112 17620 23164 17672
rect 23296 17620 23348 17672
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 25596 17756 25648 17808
rect 32956 17824 33008 17876
rect 38108 17867 38160 17876
rect 38108 17833 38117 17867
rect 38117 17833 38151 17867
rect 38151 17833 38160 17867
rect 38108 17824 38160 17833
rect 29460 17688 29512 17740
rect 31116 17688 31168 17740
rect 32496 17688 32548 17740
rect 24308 17620 24360 17672
rect 24584 17620 24636 17672
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 27620 17620 27672 17672
rect 27712 17663 27764 17672
rect 27712 17629 27721 17663
rect 27721 17629 27755 17663
rect 27755 17629 27764 17663
rect 27712 17620 27764 17629
rect 27804 17620 27856 17672
rect 30472 17620 30524 17672
rect 31852 17663 31904 17672
rect 31852 17629 31861 17663
rect 31861 17629 31895 17663
rect 31895 17629 31904 17663
rect 31852 17620 31904 17629
rect 32588 17620 32640 17672
rect 36728 17663 36780 17672
rect 36728 17629 36737 17663
rect 36737 17629 36771 17663
rect 36771 17629 36780 17663
rect 36728 17620 36780 17629
rect 37004 17663 37056 17672
rect 37004 17629 37038 17663
rect 37038 17629 37056 17663
rect 37004 17620 37056 17629
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 13084 17484 13136 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 16120 17484 16172 17536
rect 18236 17484 18288 17536
rect 23756 17552 23808 17604
rect 26424 17552 26476 17604
rect 28908 17595 28960 17604
rect 28908 17561 28917 17595
rect 28917 17561 28951 17595
rect 28951 17561 28960 17595
rect 28908 17552 28960 17561
rect 30748 17552 30800 17604
rect 32312 17552 32364 17604
rect 32864 17552 32916 17604
rect 33048 17552 33100 17604
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 26240 17484 26292 17536
rect 30932 17484 30984 17536
rect 34888 17484 34940 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8392 17212 8444 17264
rect 10508 17212 10560 17264
rect 11152 17212 11204 17264
rect 15752 17280 15804 17332
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 8944 17076 8996 17128
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 13084 17212 13136 17264
rect 12348 17076 12400 17128
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 13084 16940 13136 16992
rect 15016 17144 15068 17196
rect 15936 17144 15988 17196
rect 19432 17212 19484 17264
rect 18236 17187 18288 17196
rect 18236 17153 18270 17187
rect 18270 17153 18288 17187
rect 18236 17144 18288 17153
rect 17868 17076 17920 17128
rect 15660 17051 15712 17060
rect 15660 17017 15669 17051
rect 15669 17017 15703 17051
rect 15703 17017 15712 17051
rect 15660 17008 15712 17017
rect 17592 17008 17644 17060
rect 16212 16940 16264 16992
rect 17224 16940 17276 16992
rect 22560 17255 22612 17264
rect 22560 17221 22569 17255
rect 22569 17221 22603 17255
rect 22603 17221 22612 17255
rect 22560 17212 22612 17221
rect 23296 17212 23348 17264
rect 23664 17212 23716 17264
rect 23848 17212 23900 17264
rect 23296 17076 23348 17128
rect 24032 17144 24084 17196
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 24584 17144 24636 17153
rect 25228 17212 25280 17264
rect 28080 17212 28132 17264
rect 28632 17255 28684 17264
rect 28632 17221 28641 17255
rect 28641 17221 28675 17255
rect 28675 17221 28684 17255
rect 28632 17212 28684 17221
rect 30932 17280 30984 17332
rect 29828 17212 29880 17264
rect 30380 17212 30432 17264
rect 30656 17212 30708 17264
rect 31116 17212 31168 17264
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 25320 17187 25372 17196
rect 25320 17153 25329 17187
rect 25329 17153 25363 17187
rect 25363 17153 25372 17187
rect 25320 17144 25372 17153
rect 27988 17144 28040 17196
rect 28448 17187 28500 17196
rect 28448 17153 28458 17187
rect 28458 17153 28492 17187
rect 28492 17153 28500 17187
rect 28448 17144 28500 17153
rect 26332 17076 26384 17128
rect 27252 17076 27304 17128
rect 28264 17076 28316 17128
rect 29000 17144 29052 17196
rect 29644 17144 29696 17196
rect 30840 17144 30892 17196
rect 30380 17076 30432 17128
rect 19248 17008 19300 17060
rect 23112 17008 23164 17060
rect 28448 17008 28500 17060
rect 31852 17144 31904 17196
rect 33692 17280 33744 17332
rect 37740 17212 37792 17264
rect 33048 17144 33100 17196
rect 34520 17144 34572 17196
rect 34704 17144 34756 17196
rect 34888 17187 34940 17196
rect 34888 17153 34897 17187
rect 34897 17153 34931 17187
rect 34931 17153 34940 17187
rect 34888 17144 34940 17153
rect 32128 17076 32180 17128
rect 34796 17076 34848 17128
rect 35716 17187 35768 17196
rect 35716 17153 35725 17187
rect 35725 17153 35759 17187
rect 35759 17153 35768 17187
rect 35716 17144 35768 17153
rect 35992 17187 36044 17196
rect 35992 17153 36001 17187
rect 36001 17153 36035 17187
rect 36035 17153 36044 17187
rect 35992 17144 36044 17153
rect 36084 17187 36136 17196
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 39028 17076 39080 17128
rect 19984 16940 20036 16992
rect 22744 16983 22796 16992
rect 22744 16949 22753 16983
rect 22753 16949 22787 16983
rect 22787 16949 22796 16983
rect 22744 16940 22796 16949
rect 26148 16940 26200 16992
rect 29460 16940 29512 16992
rect 35808 17051 35860 17060
rect 35808 17017 35817 17051
rect 35817 17017 35851 17051
rect 35851 17017 35860 17051
rect 35808 17008 35860 17017
rect 37832 17008 37884 17060
rect 35716 16940 35768 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8760 16736 8812 16788
rect 9496 16736 9548 16788
rect 15660 16736 15712 16788
rect 16212 16736 16264 16788
rect 22744 16736 22796 16788
rect 27528 16736 27580 16788
rect 30472 16736 30524 16788
rect 34796 16736 34848 16788
rect 13084 16668 13136 16720
rect 17132 16668 17184 16720
rect 19156 16668 19208 16720
rect 19248 16668 19300 16720
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 8300 16600 8352 16652
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 8852 16532 8904 16584
rect 11060 16532 11112 16584
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 19432 16600 19484 16652
rect 21640 16600 21692 16652
rect 12348 16532 12400 16584
rect 16120 16575 16172 16584
rect 16120 16541 16154 16575
rect 16154 16541 16172 16575
rect 16120 16532 16172 16541
rect 6552 16464 6604 16516
rect 8392 16507 8444 16516
rect 8392 16473 8401 16507
rect 8401 16473 8435 16507
rect 8435 16473 8444 16507
rect 8392 16464 8444 16473
rect 6920 16396 6972 16448
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 12256 16464 12308 16516
rect 15292 16464 15344 16516
rect 21548 16532 21600 16584
rect 21916 16575 21968 16584
rect 21916 16541 21925 16575
rect 21925 16541 21959 16575
rect 21959 16541 21968 16575
rect 21916 16532 21968 16541
rect 23388 16600 23440 16652
rect 22744 16532 22796 16584
rect 26240 16600 26292 16652
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 27528 16600 27580 16652
rect 26516 16532 26568 16541
rect 12164 16396 12216 16448
rect 23296 16464 23348 16516
rect 26240 16464 26292 16516
rect 26424 16507 26476 16516
rect 23848 16396 23900 16448
rect 26424 16473 26433 16507
rect 26433 16473 26467 16507
rect 26467 16473 26476 16507
rect 26424 16464 26476 16473
rect 27620 16532 27672 16584
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 28172 16532 28224 16541
rect 28264 16532 28316 16584
rect 27344 16396 27396 16448
rect 28080 16464 28132 16516
rect 28448 16507 28500 16516
rect 28448 16473 28457 16507
rect 28457 16473 28491 16507
rect 28491 16473 28500 16507
rect 28448 16464 28500 16473
rect 29276 16600 29328 16652
rect 29828 16643 29880 16652
rect 29828 16609 29837 16643
rect 29837 16609 29871 16643
rect 29871 16609 29880 16643
rect 29828 16600 29880 16609
rect 29184 16532 29236 16584
rect 29736 16575 29788 16584
rect 29736 16541 29745 16575
rect 29745 16541 29779 16575
rect 29779 16541 29788 16575
rect 29736 16532 29788 16541
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 30288 16643 30340 16652
rect 30288 16609 30297 16643
rect 30297 16609 30331 16643
rect 30331 16609 30340 16643
rect 30288 16600 30340 16609
rect 30380 16600 30432 16652
rect 30932 16575 30984 16584
rect 30932 16541 30941 16575
rect 30941 16541 30975 16575
rect 30975 16541 30984 16575
rect 30932 16532 30984 16541
rect 31024 16532 31076 16584
rect 31300 16575 31352 16584
rect 31300 16541 31309 16575
rect 31309 16541 31343 16575
rect 31343 16541 31352 16575
rect 31300 16532 31352 16541
rect 31944 16532 31996 16584
rect 30748 16464 30800 16516
rect 29000 16396 29052 16448
rect 32036 16396 32088 16448
rect 32312 16575 32364 16584
rect 32312 16541 32321 16575
rect 32321 16541 32355 16575
rect 32355 16541 32364 16575
rect 32312 16532 32364 16541
rect 32496 16575 32548 16584
rect 32496 16541 32510 16575
rect 32510 16541 32544 16575
rect 32544 16541 32548 16575
rect 33600 16643 33652 16652
rect 33600 16609 33609 16643
rect 33609 16609 33643 16643
rect 33643 16609 33652 16643
rect 33600 16600 33652 16609
rect 32496 16532 32548 16541
rect 33508 16575 33560 16584
rect 33508 16541 33517 16575
rect 33517 16541 33551 16575
rect 33551 16541 33560 16575
rect 33508 16532 33560 16541
rect 33876 16643 33928 16652
rect 33876 16609 33885 16643
rect 33885 16609 33919 16643
rect 33919 16609 33928 16643
rect 33876 16600 33928 16609
rect 34704 16532 34756 16584
rect 35072 16575 35124 16584
rect 35072 16541 35076 16575
rect 35076 16541 35110 16575
rect 35110 16541 35124 16575
rect 35072 16532 35124 16541
rect 36728 16643 36780 16652
rect 36728 16609 36737 16643
rect 36737 16609 36771 16643
rect 36771 16609 36780 16643
rect 36728 16600 36780 16609
rect 35256 16507 35308 16516
rect 35256 16473 35265 16507
rect 35265 16473 35299 16507
rect 35299 16473 35308 16507
rect 35256 16464 35308 16473
rect 33048 16396 33100 16448
rect 34612 16396 34664 16448
rect 37556 16532 37608 16584
rect 37464 16464 37516 16516
rect 35440 16396 35492 16448
rect 38108 16439 38160 16448
rect 38108 16405 38117 16439
rect 38117 16405 38151 16439
rect 38151 16405 38160 16439
rect 38108 16396 38160 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 7012 16235 7064 16244
rect 7012 16201 7021 16235
rect 7021 16201 7055 16235
rect 7055 16201 7064 16235
rect 7012 16192 7064 16201
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 8944 16235 8996 16244
rect 8944 16201 8953 16235
rect 8953 16201 8987 16235
rect 8987 16201 8996 16235
rect 8944 16192 8996 16201
rect 6644 15988 6696 16040
rect 8668 16056 8720 16108
rect 10692 16192 10744 16244
rect 21548 16192 21600 16244
rect 11060 16124 11112 16176
rect 16028 16124 16080 16176
rect 10416 16056 10468 16108
rect 11520 16056 11572 16108
rect 12992 16056 13044 16108
rect 15844 16056 15896 16108
rect 16856 16056 16908 16108
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 9496 15988 9548 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 22560 16124 22612 16176
rect 22744 16124 22796 16176
rect 22928 16124 22980 16176
rect 23112 16192 23164 16244
rect 25688 16192 25740 16244
rect 24400 16124 24452 16176
rect 25964 16167 26016 16176
rect 25964 16133 25973 16167
rect 25973 16133 26007 16167
rect 26007 16133 26016 16167
rect 25964 16124 26016 16133
rect 19984 16099 20036 16108
rect 19984 16065 20018 16099
rect 20018 16065 20036 16099
rect 19984 16056 20036 16065
rect 21272 16056 21324 16108
rect 8484 15852 8536 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 17868 15988 17920 16040
rect 20720 15920 20772 15972
rect 23020 15988 23072 16040
rect 25044 16056 25096 16108
rect 25688 16099 25740 16108
rect 25688 16065 25697 16099
rect 25697 16065 25731 16099
rect 25731 16065 25740 16099
rect 25688 16056 25740 16065
rect 27620 16124 27672 16176
rect 30472 16167 30524 16176
rect 30472 16133 30481 16167
rect 30481 16133 30515 16167
rect 30515 16133 30524 16167
rect 30472 16124 30524 16133
rect 27160 16056 27212 16108
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 27436 16099 27488 16108
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 28816 16099 28868 16108
rect 28816 16065 28825 16099
rect 28825 16065 28859 16099
rect 28859 16065 28868 16099
rect 28816 16056 28868 16065
rect 28908 16099 28960 16108
rect 28908 16065 28917 16099
rect 28917 16065 28951 16099
rect 28951 16065 28960 16099
rect 28908 16056 28960 16065
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 29092 16099 29144 16108
rect 29092 16065 29101 16099
rect 29101 16065 29135 16099
rect 29135 16065 29144 16099
rect 29092 16056 29144 16065
rect 30380 16099 30432 16108
rect 30380 16065 30389 16099
rect 30389 16065 30423 16099
rect 30423 16065 30432 16099
rect 30380 16056 30432 16065
rect 30932 16056 30984 16108
rect 31116 16192 31168 16244
rect 32496 16192 32548 16244
rect 33508 16235 33560 16244
rect 33508 16201 33517 16235
rect 33517 16201 33551 16235
rect 33551 16201 33560 16235
rect 33508 16192 33560 16201
rect 32036 16124 32088 16176
rect 35072 16192 35124 16244
rect 32588 16099 32640 16108
rect 32588 16065 32597 16099
rect 32597 16065 32631 16099
rect 32631 16065 32640 16099
rect 32588 16056 32640 16065
rect 34520 16124 34572 16176
rect 17684 15895 17736 15904
rect 17684 15861 17693 15895
rect 17693 15861 17727 15895
rect 17727 15861 17736 15895
rect 17684 15852 17736 15861
rect 23388 15920 23440 15972
rect 24032 15920 24084 15972
rect 30840 16031 30892 16040
rect 30840 15997 30849 16031
rect 30849 15997 30883 16031
rect 30883 15997 30892 16031
rect 30840 15988 30892 15997
rect 31760 15988 31812 16040
rect 33048 16056 33100 16108
rect 33692 16099 33744 16108
rect 33692 16065 33701 16099
rect 33701 16065 33735 16099
rect 33735 16065 33744 16099
rect 33692 16056 33744 16065
rect 34980 15988 35032 16040
rect 35348 16056 35400 16108
rect 36084 16192 36136 16244
rect 37464 16235 37516 16244
rect 37464 16201 37473 16235
rect 37473 16201 37507 16235
rect 37507 16201 37516 16235
rect 37464 16192 37516 16201
rect 37832 16192 37884 16244
rect 38108 16056 38160 16108
rect 25044 15920 25096 15972
rect 24400 15852 24452 15904
rect 25228 15852 25280 15904
rect 25964 15895 26016 15904
rect 25964 15861 25973 15895
rect 25973 15861 26007 15895
rect 26007 15861 26016 15895
rect 25964 15852 26016 15861
rect 28080 15852 28132 15904
rect 29552 15852 29604 15904
rect 31484 15852 31536 15904
rect 32864 15895 32916 15904
rect 32864 15861 32873 15895
rect 32873 15861 32907 15895
rect 32907 15861 32916 15895
rect 32864 15852 32916 15861
rect 32956 15852 33008 15904
rect 33784 15852 33836 15904
rect 38016 16031 38068 16040
rect 38016 15997 38025 16031
rect 38025 15997 38059 16031
rect 38059 15997 38068 16031
rect 38016 15988 38068 15997
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8484 15648 8536 15700
rect 10416 15691 10468 15700
rect 10416 15657 10425 15691
rect 10425 15657 10459 15691
rect 10459 15657 10468 15691
rect 10416 15648 10468 15657
rect 13452 15648 13504 15700
rect 27160 15691 27212 15700
rect 27160 15657 27169 15691
rect 27169 15657 27203 15691
rect 27203 15657 27212 15691
rect 27160 15648 27212 15657
rect 28816 15648 28868 15700
rect 11704 15580 11756 15632
rect 11152 15512 11204 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 7748 15444 7800 15496
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 10232 15444 10284 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 14280 15444 14332 15496
rect 18420 15580 18472 15632
rect 18512 15623 18564 15632
rect 18512 15589 18521 15623
rect 18521 15589 18555 15623
rect 18555 15589 18564 15623
rect 18512 15580 18564 15589
rect 20260 15580 20312 15632
rect 26424 15580 26476 15632
rect 34704 15648 34756 15700
rect 35992 15648 36044 15700
rect 8392 15376 8444 15428
rect 11980 15376 12032 15428
rect 30840 15580 30892 15632
rect 11796 15308 11848 15360
rect 16856 15376 16908 15428
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 17500 15376 17552 15428
rect 20352 15444 20404 15496
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 21640 15487 21692 15496
rect 21640 15453 21644 15487
rect 21644 15453 21678 15487
rect 21678 15453 21692 15487
rect 21640 15444 21692 15453
rect 21824 15419 21876 15428
rect 21824 15385 21833 15419
rect 21833 15385 21867 15419
rect 21867 15385 21876 15419
rect 21824 15376 21876 15385
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22928 15444 22980 15496
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 24860 15487 24912 15496
rect 24860 15453 24869 15487
rect 24869 15453 24903 15487
rect 24903 15453 24912 15487
rect 24860 15444 24912 15453
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 25872 15444 25924 15496
rect 30380 15555 30432 15564
rect 30380 15521 30389 15555
rect 30389 15521 30423 15555
rect 30423 15521 30432 15555
rect 30380 15512 30432 15521
rect 31484 15555 31536 15564
rect 31484 15521 31493 15555
rect 31493 15521 31527 15555
rect 31527 15521 31536 15555
rect 31484 15512 31536 15521
rect 35440 15555 35492 15564
rect 35440 15521 35449 15555
rect 35449 15521 35483 15555
rect 35483 15521 35492 15555
rect 35440 15512 35492 15521
rect 37740 15512 37792 15564
rect 38016 15580 38068 15632
rect 27528 15444 27580 15496
rect 29092 15444 29144 15496
rect 29184 15487 29236 15496
rect 29184 15453 29193 15487
rect 29193 15453 29227 15487
rect 29227 15453 29236 15487
rect 29184 15444 29236 15453
rect 32220 15444 32272 15496
rect 35348 15487 35400 15496
rect 35348 15453 35357 15487
rect 35357 15453 35391 15487
rect 35391 15453 35400 15487
rect 35348 15444 35400 15453
rect 12164 15308 12216 15360
rect 20720 15308 20772 15360
rect 24492 15376 24544 15428
rect 28448 15376 28500 15428
rect 34980 15419 35032 15428
rect 34980 15385 34989 15419
rect 34989 15385 35023 15419
rect 35023 15385 35032 15419
rect 34980 15376 35032 15385
rect 35072 15419 35124 15428
rect 35072 15385 35081 15419
rect 35081 15385 35115 15419
rect 35115 15385 35124 15419
rect 35072 15376 35124 15385
rect 37556 15376 37608 15428
rect 25412 15308 25464 15360
rect 31024 15351 31076 15360
rect 31024 15317 31033 15351
rect 31033 15317 31067 15351
rect 31067 15317 31076 15351
rect 31024 15308 31076 15317
rect 31760 15308 31812 15360
rect 32588 15308 32640 15360
rect 32864 15308 32916 15360
rect 35716 15308 35768 15360
rect 37188 15308 37240 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9864 15104 9916 15156
rect 14556 15104 14608 15156
rect 18052 15104 18104 15156
rect 7840 15036 7892 15088
rect 9128 15036 9180 15088
rect 11980 15079 12032 15088
rect 11980 15045 11989 15079
rect 11989 15045 12023 15079
rect 12023 15045 12032 15079
rect 11980 15036 12032 15045
rect 15292 15036 15344 15088
rect 16488 15036 16540 15088
rect 8392 14968 8444 15020
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 13268 14968 13320 15020
rect 16396 14968 16448 15020
rect 9496 14900 9548 14952
rect 12072 14900 12124 14952
rect 12348 14900 12400 14952
rect 12900 14900 12952 14952
rect 16212 14900 16264 14952
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 17316 15011 17368 15020
rect 17316 14977 17325 15011
rect 17325 14977 17359 15011
rect 17359 14977 17368 15011
rect 17316 14968 17368 14977
rect 18420 15036 18472 15088
rect 18788 15036 18840 15088
rect 21916 15036 21968 15088
rect 17776 14968 17828 15020
rect 21640 14968 21692 15020
rect 23848 15104 23900 15156
rect 24860 15104 24912 15156
rect 27436 15104 27488 15156
rect 18236 14900 18288 14952
rect 17500 14832 17552 14884
rect 18052 14875 18104 14884
rect 18052 14841 18061 14875
rect 18061 14841 18095 14875
rect 18095 14841 18104 14875
rect 18052 14832 18104 14841
rect 18144 14832 18196 14884
rect 19984 14875 20036 14884
rect 19984 14841 19993 14875
rect 19993 14841 20027 14875
rect 20027 14841 20036 14875
rect 19984 14832 20036 14841
rect 20352 14943 20404 14952
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 20628 14900 20680 14952
rect 23204 14968 23256 15020
rect 23572 14968 23624 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24400 15011 24452 15020
rect 24400 14977 24409 15011
rect 24409 14977 24443 15011
rect 24443 14977 24452 15011
rect 24400 14968 24452 14977
rect 25412 15011 25464 15020
rect 25412 14977 25421 15011
rect 25421 14977 25455 15011
rect 25455 14977 25464 15011
rect 25412 14968 25464 14977
rect 25596 15011 25648 15020
rect 25596 14977 25605 15011
rect 25605 14977 25639 15011
rect 25639 14977 25648 15011
rect 25596 14968 25648 14977
rect 24952 14900 25004 14952
rect 25044 14900 25096 14952
rect 26240 14968 26292 15020
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 27528 14900 27580 14952
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 16212 14764 16264 14816
rect 16948 14764 17000 14816
rect 17868 14764 17920 14816
rect 20168 14764 20220 14816
rect 20352 14764 20404 14816
rect 23112 14764 23164 14816
rect 24492 14764 24544 14816
rect 28172 14764 28224 14816
rect 28356 15011 28408 15020
rect 28356 14977 28365 15011
rect 28365 14977 28399 15011
rect 28399 14977 28408 15011
rect 28356 14968 28408 14977
rect 31760 15147 31812 15156
rect 31760 15113 31769 15147
rect 31769 15113 31803 15147
rect 31803 15113 31812 15147
rect 31760 15104 31812 15113
rect 31024 15036 31076 15088
rect 31300 15036 31352 15088
rect 34980 15104 35032 15156
rect 35440 15104 35492 15156
rect 33876 15036 33928 15088
rect 38108 15079 38160 15088
rect 38108 15045 38117 15079
rect 38117 15045 38151 15079
rect 38151 15045 38160 15079
rect 38108 15036 38160 15045
rect 30932 14968 30984 15020
rect 35348 14968 35400 15020
rect 35716 14968 35768 15020
rect 29000 14900 29052 14952
rect 29644 14900 29696 14952
rect 30380 14943 30432 14952
rect 30380 14909 30389 14943
rect 30389 14909 30423 14943
rect 30423 14909 30432 14943
rect 30380 14900 30432 14909
rect 32220 14900 32272 14952
rect 33416 14900 33468 14952
rect 33968 14832 34020 14884
rect 34520 14764 34572 14816
rect 35716 14764 35768 14816
rect 35992 14807 36044 14816
rect 35992 14773 36001 14807
rect 36001 14773 36035 14807
rect 36035 14773 36044 14807
rect 35992 14764 36044 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 12900 14560 12952 14612
rect 13268 14603 13320 14612
rect 13268 14569 13277 14603
rect 13277 14569 13311 14603
rect 13311 14569 13320 14603
rect 13268 14560 13320 14569
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 18236 14560 18288 14612
rect 24400 14560 24452 14612
rect 25596 14560 25648 14612
rect 27344 14560 27396 14612
rect 27528 14560 27580 14612
rect 29276 14560 29328 14612
rect 31668 14560 31720 14612
rect 35992 14560 36044 14612
rect 36360 14560 36412 14612
rect 37556 14560 37608 14612
rect 13360 14535 13412 14544
rect 13360 14501 13369 14535
rect 13369 14501 13403 14535
rect 13403 14501 13412 14535
rect 13360 14492 13412 14501
rect 21364 14492 21416 14544
rect 26240 14492 26292 14544
rect 31300 14492 31352 14544
rect 10508 14424 10560 14476
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 24952 14467 25004 14476
rect 24952 14433 24961 14467
rect 24961 14433 24995 14467
rect 24995 14433 25004 14467
rect 24952 14424 25004 14433
rect 25320 14424 25372 14476
rect 32956 14535 33008 14544
rect 32956 14501 32965 14535
rect 32965 14501 32999 14535
rect 32999 14501 33008 14535
rect 32956 14492 33008 14501
rect 34520 14492 34572 14544
rect 35624 14492 35676 14544
rect 33048 14424 33100 14476
rect 35440 14467 35492 14476
rect 35440 14433 35449 14467
rect 35449 14433 35483 14467
rect 35483 14433 35492 14467
rect 35440 14424 35492 14433
rect 35716 14424 35768 14476
rect 11796 14356 11848 14408
rect 12256 14288 12308 14340
rect 14188 14356 14240 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 17592 14356 17644 14408
rect 12900 14288 12952 14340
rect 14004 14288 14056 14340
rect 15108 14331 15160 14340
rect 15108 14297 15117 14331
rect 15117 14297 15151 14331
rect 15151 14297 15160 14331
rect 15108 14288 15160 14297
rect 15476 14331 15528 14340
rect 15476 14297 15485 14331
rect 15485 14297 15519 14331
rect 15519 14297 15528 14331
rect 15476 14288 15528 14297
rect 18512 14288 18564 14340
rect 18788 14356 18840 14408
rect 18972 14356 19024 14408
rect 21640 14399 21692 14408
rect 21640 14365 21644 14399
rect 21644 14365 21678 14399
rect 21678 14365 21692 14399
rect 21640 14356 21692 14365
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 21916 14356 21968 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 23940 14399 23992 14408
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 24400 14356 24452 14408
rect 24492 14356 24544 14408
rect 15200 14220 15252 14272
rect 17224 14220 17276 14272
rect 17776 14220 17828 14272
rect 18880 14220 18932 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 20996 14288 21048 14340
rect 26608 14356 26660 14408
rect 27160 14356 27212 14408
rect 30656 14356 30708 14408
rect 35348 14356 35400 14408
rect 37188 14399 37240 14408
rect 37188 14365 37222 14399
rect 37222 14365 37240 14399
rect 29828 14288 29880 14340
rect 35532 14331 35584 14340
rect 20812 14220 20864 14272
rect 21088 14220 21140 14272
rect 23480 14220 23532 14272
rect 24216 14220 24268 14272
rect 24952 14220 25004 14272
rect 29000 14220 29052 14272
rect 29092 14220 29144 14272
rect 35532 14297 35541 14331
rect 35541 14297 35575 14331
rect 35575 14297 35584 14331
rect 35532 14288 35584 14297
rect 35624 14288 35676 14340
rect 37188 14356 37240 14365
rect 33692 14220 33744 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9864 14016 9916 14068
rect 13176 14016 13228 14068
rect 17316 14016 17368 14068
rect 9496 13948 9548 14000
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 11796 13948 11848 14000
rect 14188 13948 14240 14000
rect 15476 13948 15528 14000
rect 18144 13948 18196 14000
rect 18236 13948 18288 14000
rect 11888 13812 11940 13864
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 14004 13880 14056 13932
rect 14556 13880 14608 13932
rect 15108 13880 15160 13932
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 17040 13880 17092 13932
rect 17500 13880 17552 13932
rect 17776 13880 17828 13932
rect 18880 14016 18932 14068
rect 24124 14016 24176 14068
rect 30932 14016 30984 14068
rect 13360 13812 13412 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 17408 13812 17460 13864
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 19984 13948 20036 14000
rect 25596 13948 25648 14000
rect 19432 13812 19484 13864
rect 20076 13880 20128 13932
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 20352 13812 20404 13864
rect 13820 13744 13872 13796
rect 15844 13744 15896 13796
rect 10232 13676 10284 13728
rect 10968 13676 11020 13728
rect 15568 13676 15620 13728
rect 23480 13880 23532 13932
rect 23756 13923 23808 13932
rect 23756 13889 23765 13923
rect 23765 13889 23799 13923
rect 23799 13889 23808 13923
rect 23756 13880 23808 13889
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 24216 13880 24268 13932
rect 25688 13880 25740 13932
rect 26056 13991 26108 14000
rect 26056 13957 26065 13991
rect 26065 13957 26099 13991
rect 26099 13957 26108 13991
rect 26056 13948 26108 13957
rect 27988 13991 28040 14000
rect 27988 13957 27997 13991
rect 27997 13957 28031 13991
rect 28031 13957 28040 13991
rect 27988 13948 28040 13957
rect 28448 13991 28500 14000
rect 28448 13957 28457 13991
rect 28457 13957 28491 13991
rect 28491 13957 28500 13991
rect 28448 13948 28500 13957
rect 28540 13948 28592 14000
rect 29092 13948 29144 14000
rect 29644 13948 29696 14000
rect 24308 13812 24360 13864
rect 23296 13744 23348 13796
rect 24492 13744 24544 13796
rect 23664 13676 23716 13728
rect 24860 13812 24912 13864
rect 27160 13880 27212 13932
rect 27436 13812 27488 13864
rect 27896 13880 27948 13932
rect 28540 13812 28592 13864
rect 29000 13923 29052 13932
rect 29000 13889 29009 13923
rect 29009 13889 29043 13923
rect 29043 13889 29052 13923
rect 29000 13880 29052 13889
rect 29460 13923 29512 13932
rect 29460 13889 29469 13923
rect 29469 13889 29503 13923
rect 29503 13889 29512 13923
rect 29460 13880 29512 13889
rect 35624 13948 35676 14000
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 31300 13923 31352 13932
rect 31300 13889 31309 13923
rect 31309 13889 31343 13923
rect 31343 13889 31352 13923
rect 31300 13880 31352 13889
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 29736 13812 29788 13864
rect 31024 13855 31076 13864
rect 31024 13821 31033 13855
rect 31033 13821 31067 13855
rect 31067 13821 31076 13855
rect 31024 13812 31076 13821
rect 32312 13812 32364 13864
rect 33600 13812 33652 13864
rect 38292 13855 38344 13864
rect 38292 13821 38301 13855
rect 38301 13821 38335 13855
rect 38335 13821 38344 13855
rect 38292 13812 38344 13821
rect 28908 13744 28960 13796
rect 25596 13676 25648 13728
rect 27988 13719 28040 13728
rect 27988 13685 27997 13719
rect 27997 13685 28031 13719
rect 28031 13685 28040 13719
rect 27988 13676 28040 13685
rect 30012 13676 30064 13728
rect 34796 13676 34848 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 15016 13472 15068 13524
rect 10508 13447 10560 13456
rect 10508 13413 10517 13447
rect 10517 13413 10551 13447
rect 10551 13413 10560 13447
rect 10508 13404 10560 13413
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 15292 13336 15344 13388
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 22468 13472 22520 13524
rect 23296 13472 23348 13524
rect 23756 13472 23808 13524
rect 26332 13472 26384 13524
rect 29184 13472 29236 13524
rect 31024 13472 31076 13524
rect 33232 13472 33284 13524
rect 15752 13336 15804 13388
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 16580 13336 16632 13388
rect 14004 13132 14056 13184
rect 15660 13132 15712 13184
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 20812 13311 20864 13320
rect 20812 13277 20821 13311
rect 20821 13277 20855 13311
rect 20855 13277 20864 13311
rect 20812 13268 20864 13277
rect 21364 13336 21416 13388
rect 21272 13268 21324 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 21732 13379 21784 13388
rect 21732 13345 21741 13379
rect 21741 13345 21775 13379
rect 21775 13345 21784 13379
rect 21732 13336 21784 13345
rect 23664 13379 23716 13388
rect 23664 13345 23673 13379
rect 23673 13345 23707 13379
rect 23707 13345 23716 13379
rect 23664 13336 23716 13345
rect 24216 13336 24268 13388
rect 29644 13404 29696 13456
rect 25964 13336 26016 13388
rect 26608 13336 26660 13388
rect 22008 13268 22060 13320
rect 23480 13268 23532 13320
rect 19524 13200 19576 13252
rect 22376 13200 22428 13252
rect 24032 13268 24084 13320
rect 24492 13268 24544 13320
rect 24768 13200 24820 13252
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 26516 13243 26568 13252
rect 26516 13209 26525 13243
rect 26525 13209 26559 13243
rect 26559 13209 26568 13243
rect 26516 13200 26568 13209
rect 26792 13268 26844 13320
rect 27252 13311 27304 13320
rect 27252 13277 27261 13311
rect 27261 13277 27295 13311
rect 27295 13277 27304 13311
rect 27252 13268 27304 13277
rect 27988 13336 28040 13388
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 32956 13447 33008 13456
rect 32956 13413 32965 13447
rect 32965 13413 32999 13447
rect 32999 13413 33008 13447
rect 32956 13404 33008 13413
rect 32864 13336 32916 13388
rect 34612 13336 34664 13388
rect 35716 13379 35768 13388
rect 35716 13345 35725 13379
rect 35725 13345 35759 13379
rect 35759 13345 35768 13379
rect 35716 13336 35768 13345
rect 27436 13200 27488 13252
rect 29092 13268 29144 13320
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 33232 13268 33284 13320
rect 33692 13311 33744 13320
rect 33692 13277 33701 13311
rect 33701 13277 33735 13311
rect 33735 13277 33744 13311
rect 33692 13268 33744 13277
rect 34796 13268 34848 13320
rect 22192 13132 22244 13184
rect 22468 13132 22520 13184
rect 33784 13132 33836 13184
rect 35808 13132 35860 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12900 12928 12952 12980
rect 21272 12928 21324 12980
rect 22468 12928 22520 12980
rect 23664 12928 23716 12980
rect 27252 12928 27304 12980
rect 34704 12928 34756 12980
rect 7840 12860 7892 12912
rect 13268 12860 13320 12912
rect 15476 12903 15528 12912
rect 15476 12869 15485 12903
rect 15485 12869 15519 12903
rect 15519 12869 15528 12903
rect 15476 12860 15528 12869
rect 15568 12903 15620 12912
rect 15568 12869 15577 12903
rect 15577 12869 15611 12903
rect 15611 12869 15620 12903
rect 15568 12860 15620 12869
rect 16120 12860 16172 12912
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 10416 12724 10468 12776
rect 12716 12792 12768 12844
rect 12900 12724 12952 12776
rect 13176 12724 13228 12776
rect 13636 12792 13688 12844
rect 15200 12792 15252 12844
rect 16580 12792 16632 12844
rect 17316 12792 17368 12844
rect 17684 12792 17736 12844
rect 21180 12835 21232 12844
rect 21180 12801 21189 12835
rect 21189 12801 21223 12835
rect 21223 12801 21232 12835
rect 21180 12792 21232 12801
rect 21364 12792 21416 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 17500 12724 17552 12776
rect 26516 12860 26568 12912
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 23480 12835 23532 12844
rect 23480 12801 23489 12835
rect 23489 12801 23523 12835
rect 23523 12801 23532 12835
rect 23480 12792 23532 12801
rect 23940 12792 23992 12844
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 26608 12792 26660 12844
rect 27896 12835 27948 12844
rect 27896 12801 27905 12835
rect 27905 12801 27939 12835
rect 27939 12801 27948 12835
rect 27896 12792 27948 12801
rect 29368 12792 29420 12844
rect 33140 12792 33192 12844
rect 34612 12860 34664 12912
rect 33784 12792 33836 12844
rect 26332 12724 26384 12776
rect 27804 12724 27856 12776
rect 15292 12656 15344 12708
rect 17684 12656 17736 12708
rect 21916 12656 21968 12708
rect 11060 12588 11112 12640
rect 17224 12588 17276 12640
rect 17868 12588 17920 12640
rect 20996 12588 21048 12640
rect 21640 12588 21692 12640
rect 38292 12631 38344 12640
rect 38292 12597 38301 12631
rect 38301 12597 38335 12631
rect 38335 12597 38344 12631
rect 38292 12588 38344 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10968 12427 11020 12436
rect 10968 12393 10977 12427
rect 10977 12393 11011 12427
rect 11011 12393 11020 12427
rect 10968 12384 11020 12393
rect 13544 12359 13596 12368
rect 13544 12325 13553 12359
rect 13553 12325 13587 12359
rect 13587 12325 13596 12359
rect 13544 12316 13596 12325
rect 7840 12248 7892 12300
rect 8760 12248 8812 12300
rect 11704 12248 11756 12300
rect 10324 12180 10376 12232
rect 12164 12180 12216 12232
rect 12716 12248 12768 12300
rect 16764 12316 16816 12368
rect 17868 12384 17920 12436
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 15568 12248 15620 12300
rect 16672 12248 16724 12300
rect 18236 12316 18288 12368
rect 11152 12112 11204 12164
rect 12348 12112 12400 12164
rect 12900 12112 12952 12164
rect 13176 12112 13228 12164
rect 15752 12180 15804 12232
rect 15936 12180 15988 12232
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17500 12248 17552 12300
rect 17960 12248 18012 12300
rect 18880 12248 18932 12300
rect 19340 12316 19392 12368
rect 21180 12384 21232 12436
rect 25872 12384 25924 12436
rect 27804 12384 27856 12436
rect 29092 12384 29144 12436
rect 22100 12316 22152 12368
rect 31392 12316 31444 12368
rect 20628 12248 20680 12300
rect 24584 12248 24636 12300
rect 25320 12248 25372 12300
rect 31484 12248 31536 12300
rect 32772 12248 32824 12300
rect 38016 12384 38068 12436
rect 35808 12248 35860 12300
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 11980 12044 12032 12096
rect 14188 12044 14240 12096
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 16120 12155 16172 12164
rect 16120 12121 16129 12155
rect 16129 12121 16163 12155
rect 16163 12121 16172 12155
rect 16120 12112 16172 12121
rect 17408 12112 17460 12164
rect 16672 12044 16724 12096
rect 17684 12044 17736 12096
rect 17776 12044 17828 12096
rect 18696 12180 18748 12232
rect 20260 12180 20312 12232
rect 20536 12180 20588 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 21548 12180 21600 12232
rect 20168 12112 20220 12164
rect 18972 12044 19024 12096
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 27436 12223 27488 12232
rect 27436 12189 27445 12223
rect 27445 12189 27479 12223
rect 27479 12189 27488 12223
rect 27436 12180 27488 12189
rect 27620 12180 27672 12232
rect 31576 12180 31628 12232
rect 25964 12112 26016 12164
rect 25596 12044 25648 12096
rect 27528 12087 27580 12096
rect 27528 12053 27537 12087
rect 27537 12053 27571 12087
rect 27571 12053 27580 12087
rect 27528 12044 27580 12053
rect 30564 12044 30616 12096
rect 31668 12112 31720 12164
rect 34612 12180 34664 12232
rect 32864 12112 32916 12164
rect 37924 12180 37976 12232
rect 37464 12112 37516 12164
rect 32220 12044 32272 12096
rect 32312 12087 32364 12096
rect 32312 12053 32321 12087
rect 32321 12053 32355 12087
rect 32355 12053 32364 12087
rect 32312 12044 32364 12053
rect 32680 12087 32732 12096
rect 32680 12053 32689 12087
rect 32689 12053 32723 12087
rect 32723 12053 32732 12087
rect 32680 12044 32732 12053
rect 32772 12087 32824 12096
rect 32772 12053 32781 12087
rect 32781 12053 32815 12087
rect 32815 12053 32824 12087
rect 32772 12044 32824 12053
rect 35348 12044 35400 12096
rect 35440 12087 35492 12096
rect 35440 12053 35449 12087
rect 35449 12053 35483 12087
rect 35483 12053 35492 12087
rect 35440 12044 35492 12053
rect 37832 12044 37884 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 7840 11840 7892 11892
rect 9404 11840 9456 11892
rect 12256 11840 12308 11892
rect 10784 11772 10836 11824
rect 11060 11704 11112 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12348 11772 12400 11824
rect 15200 11840 15252 11892
rect 16488 11840 16540 11892
rect 13268 11772 13320 11824
rect 16120 11772 16172 11824
rect 17132 11772 17184 11824
rect 17776 11772 17828 11824
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 14004 11704 14056 11756
rect 15476 11704 15528 11756
rect 15660 11704 15712 11756
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 12900 11611 12952 11620
rect 12900 11577 12909 11611
rect 12909 11577 12943 11611
rect 12943 11577 12952 11611
rect 12900 11568 12952 11577
rect 15936 11636 15988 11688
rect 16028 11636 16080 11688
rect 15752 11568 15804 11620
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 21364 11840 21416 11892
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 25228 11883 25280 11892
rect 25228 11849 25237 11883
rect 25237 11849 25271 11883
rect 25271 11849 25280 11883
rect 25228 11840 25280 11849
rect 32680 11840 32732 11892
rect 33508 11840 33560 11892
rect 34520 11840 34572 11892
rect 37464 11883 37516 11892
rect 37464 11849 37473 11883
rect 37473 11849 37507 11883
rect 37507 11849 37516 11883
rect 37464 11840 37516 11849
rect 37832 11883 37884 11892
rect 37832 11849 37841 11883
rect 37841 11849 37875 11883
rect 37875 11849 37884 11883
rect 37832 11840 37884 11849
rect 37924 11883 37976 11892
rect 37924 11849 37933 11883
rect 37933 11849 37967 11883
rect 37967 11849 37976 11883
rect 37924 11840 37976 11849
rect 21732 11704 21784 11756
rect 22560 11704 22612 11756
rect 19984 11636 20036 11688
rect 21640 11636 21692 11688
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 11980 11500 12032 11552
rect 17316 11500 17368 11552
rect 18512 11500 18564 11552
rect 19156 11543 19208 11552
rect 19156 11509 19165 11543
rect 19165 11509 19199 11543
rect 19199 11509 19208 11543
rect 19156 11500 19208 11509
rect 19432 11568 19484 11620
rect 21272 11568 21324 11620
rect 25872 11704 25924 11756
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26240 11704 26292 11713
rect 30380 11704 30432 11756
rect 30564 11747 30616 11756
rect 30564 11713 30598 11747
rect 30598 11713 30616 11747
rect 30564 11704 30616 11713
rect 29092 11636 29144 11688
rect 32312 11772 32364 11824
rect 35716 11704 35768 11756
rect 35992 11747 36044 11756
rect 35992 11713 36001 11747
rect 36001 11713 36035 11747
rect 36035 11713 36044 11747
rect 35992 11704 36044 11713
rect 25964 11611 26016 11620
rect 25964 11577 25973 11611
rect 25973 11577 26007 11611
rect 26007 11577 26016 11611
rect 25964 11568 26016 11577
rect 19800 11500 19852 11552
rect 20444 11500 20496 11552
rect 20628 11500 20680 11552
rect 26240 11500 26292 11552
rect 31668 11543 31720 11552
rect 31668 11509 31677 11543
rect 31677 11509 31711 11543
rect 31711 11509 31720 11543
rect 31668 11500 31720 11509
rect 35440 11636 35492 11688
rect 36268 11679 36320 11688
rect 36268 11645 36277 11679
rect 36277 11645 36311 11679
rect 36311 11645 36320 11679
rect 36268 11636 36320 11645
rect 38016 11679 38068 11688
rect 38016 11645 38025 11679
rect 38025 11645 38059 11679
rect 38059 11645 38068 11679
rect 38016 11636 38068 11645
rect 33048 11500 33100 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 10324 11339 10376 11348
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 12164 11296 12216 11348
rect 17960 11296 18012 11348
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 19892 11296 19944 11348
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 21916 11339 21968 11348
rect 21916 11305 21925 11339
rect 21925 11305 21959 11339
rect 21959 11305 21968 11339
rect 21916 11296 21968 11305
rect 25688 11339 25740 11348
rect 25688 11305 25697 11339
rect 25697 11305 25731 11339
rect 25731 11305 25740 11339
rect 25688 11296 25740 11305
rect 25872 11339 25924 11348
rect 25872 11305 25881 11339
rect 25881 11305 25915 11339
rect 25915 11305 25924 11339
rect 25872 11296 25924 11305
rect 12348 11228 12400 11280
rect 10416 11092 10468 11144
rect 11704 11160 11756 11212
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 11888 11092 11940 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 16488 11228 16540 11280
rect 18512 11228 18564 11280
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 14096 11024 14148 11076
rect 11336 10956 11388 11008
rect 16304 11024 16356 11076
rect 16580 11092 16632 11144
rect 17224 11092 17276 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 18972 11160 19024 11212
rect 19524 11092 19576 11144
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 21456 11092 21508 11144
rect 22284 11228 22336 11280
rect 21732 11160 21784 11212
rect 22192 11092 22244 11144
rect 25780 11228 25832 11280
rect 27620 11296 27672 11348
rect 27896 11271 27948 11280
rect 27896 11237 27905 11271
rect 27905 11237 27939 11271
rect 27939 11237 27948 11271
rect 33140 11296 33192 11348
rect 35532 11296 35584 11348
rect 27896 11228 27948 11237
rect 27620 11160 27672 11212
rect 29092 11203 29144 11212
rect 29092 11169 29101 11203
rect 29101 11169 29135 11203
rect 29135 11169 29144 11203
rect 29092 11160 29144 11169
rect 29368 11160 29420 11212
rect 21088 11024 21140 11076
rect 17684 10956 17736 11008
rect 17868 10956 17920 11008
rect 24860 11024 24912 11076
rect 25504 11067 25556 11076
rect 25504 11033 25513 11067
rect 25513 11033 25547 11067
rect 25547 11033 25556 11067
rect 25504 11024 25556 11033
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27712 11092 27764 11144
rect 29644 11092 29696 11144
rect 33416 11228 33468 11280
rect 31668 11160 31720 11212
rect 34612 11160 34664 11212
rect 27160 11024 27212 11076
rect 29920 11024 29972 11076
rect 31300 11024 31352 11076
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 33140 11135 33192 11144
rect 33140 11101 33149 11135
rect 33149 11101 33183 11135
rect 33183 11101 33192 11135
rect 33140 11092 33192 11101
rect 33508 11135 33560 11144
rect 33508 11101 33517 11135
rect 33517 11101 33551 11135
rect 33551 11101 33560 11135
rect 33508 11092 33560 11101
rect 22100 10999 22152 11008
rect 22100 10965 22109 10999
rect 22109 10965 22143 10999
rect 22143 10965 22152 10999
rect 22100 10956 22152 10965
rect 22376 10956 22428 11008
rect 28448 10999 28500 11008
rect 28448 10965 28457 10999
rect 28457 10965 28491 10999
rect 28491 10965 28500 10999
rect 28448 10956 28500 10965
rect 31484 10956 31536 11008
rect 34520 10956 34572 11008
rect 35348 11024 35400 11076
rect 36268 11024 36320 11076
rect 37464 11024 37516 11076
rect 38200 10999 38252 11008
rect 38200 10965 38209 10999
rect 38209 10965 38243 10999
rect 38243 10965 38252 10999
rect 38200 10956 38252 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 17316 10752 17368 10804
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 14740 10684 14792 10736
rect 17776 10684 17828 10736
rect 18144 10684 18196 10736
rect 26884 10752 26936 10804
rect 27160 10795 27212 10804
rect 27160 10761 27169 10795
rect 27169 10761 27203 10795
rect 27203 10761 27212 10795
rect 27160 10752 27212 10761
rect 27896 10752 27948 10804
rect 29920 10752 29972 10804
rect 37464 10795 37516 10804
rect 37464 10761 37473 10795
rect 37473 10761 37507 10795
rect 37507 10761 37516 10795
rect 37464 10752 37516 10761
rect 22284 10727 22336 10736
rect 22284 10693 22293 10727
rect 22293 10693 22327 10727
rect 22327 10693 22336 10727
rect 22284 10684 22336 10693
rect 22376 10727 22428 10736
rect 22376 10693 22385 10727
rect 22385 10693 22419 10727
rect 22419 10693 22428 10727
rect 22376 10684 22428 10693
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 14188 10616 14240 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 26516 10684 26568 10736
rect 27620 10727 27672 10736
rect 27620 10693 27629 10727
rect 27629 10693 27663 10727
rect 27663 10693 27672 10727
rect 27620 10684 27672 10693
rect 27712 10684 27764 10736
rect 28448 10684 28500 10736
rect 24676 10659 24728 10668
rect 24676 10625 24710 10659
rect 24710 10625 24728 10659
rect 10324 10548 10376 10600
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 22100 10548 22152 10600
rect 24676 10616 24728 10625
rect 26148 10616 26200 10668
rect 34152 10659 34204 10668
rect 34152 10625 34161 10659
rect 34161 10625 34195 10659
rect 34195 10625 34204 10659
rect 34152 10616 34204 10625
rect 17776 10480 17828 10532
rect 22652 10480 22704 10532
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 13544 10412 13596 10464
rect 20904 10412 20956 10464
rect 25136 10412 25188 10464
rect 25504 10412 25556 10464
rect 27804 10591 27856 10600
rect 27804 10557 27813 10591
rect 27813 10557 27847 10591
rect 27847 10557 27856 10591
rect 27804 10548 27856 10557
rect 33968 10548 34020 10600
rect 37648 10684 37700 10736
rect 37372 10616 37424 10668
rect 38200 10616 38252 10668
rect 34520 10548 34572 10600
rect 35808 10548 35860 10600
rect 38016 10591 38068 10600
rect 38016 10557 38025 10591
rect 38025 10557 38059 10591
rect 38059 10557 38068 10591
rect 38016 10548 38068 10557
rect 33784 10455 33836 10464
rect 33784 10421 33793 10455
rect 33793 10421 33827 10455
rect 33827 10421 33836 10455
rect 33784 10412 33836 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 10876 10208 10928 10260
rect 17408 10208 17460 10260
rect 17684 10208 17736 10260
rect 14188 10140 14240 10192
rect 11060 10072 11112 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 19432 10140 19484 10192
rect 22192 10208 22244 10260
rect 24676 10208 24728 10260
rect 32220 10208 32272 10260
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11796 10004 11848 10056
rect 11244 9936 11296 9988
rect 14832 10004 14884 10056
rect 15292 10004 15344 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 15200 9868 15252 9920
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 20076 10072 20128 10124
rect 20720 10072 20772 10124
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 21456 10004 21508 10056
rect 34152 10140 34204 10192
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 27804 10072 27856 10124
rect 34428 10140 34480 10192
rect 36268 10115 36320 10124
rect 36268 10081 36277 10115
rect 36277 10081 36311 10115
rect 36311 10081 36320 10115
rect 36268 10072 36320 10081
rect 25136 10047 25188 10056
rect 25136 10013 25145 10047
rect 25145 10013 25179 10047
rect 25179 10013 25188 10047
rect 25136 10004 25188 10013
rect 32036 10047 32088 10056
rect 32036 10013 32045 10047
rect 32045 10013 32079 10047
rect 32079 10013 32088 10047
rect 32036 10004 32088 10013
rect 32128 10047 32180 10056
rect 32128 10013 32137 10047
rect 32137 10013 32171 10047
rect 32171 10013 32180 10047
rect 32128 10004 32180 10013
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 20904 9868 20956 9920
rect 33048 10004 33100 10056
rect 33784 10004 33836 10056
rect 35440 10004 35492 10056
rect 35992 10047 36044 10056
rect 35992 10013 36001 10047
rect 36001 10013 36035 10047
rect 36035 10013 36044 10047
rect 35992 10004 36044 10013
rect 36360 10004 36412 10056
rect 37372 10072 37424 10124
rect 39028 10072 39080 10124
rect 37832 10047 37884 10056
rect 37832 10013 37841 10047
rect 37841 10013 37875 10047
rect 37875 10013 37884 10047
rect 37832 10004 37884 10013
rect 33876 9936 33928 9988
rect 32956 9868 33008 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 10876 9707 10928 9716
rect 10876 9673 10885 9707
rect 10885 9673 10919 9707
rect 10919 9673 10928 9707
rect 10876 9664 10928 9673
rect 10416 9639 10468 9648
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 11336 9596 11388 9648
rect 13452 9664 13504 9716
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 20720 9707 20772 9716
rect 20720 9673 20729 9707
rect 20729 9673 20763 9707
rect 20763 9673 20772 9707
rect 20720 9664 20772 9673
rect 22560 9664 22612 9716
rect 26516 9664 26568 9716
rect 27804 9664 27856 9716
rect 28448 9664 28500 9716
rect 10508 9528 10560 9580
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 11244 9528 11296 9580
rect 11520 9528 11572 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 14004 9639 14056 9648
rect 14004 9605 14013 9639
rect 14013 9605 14047 9639
rect 14047 9605 14056 9639
rect 14004 9596 14056 9605
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 15200 9596 15252 9648
rect 15476 9528 15528 9580
rect 16028 9528 16080 9580
rect 22468 9596 22520 9648
rect 25228 9596 25280 9648
rect 25596 9639 25648 9648
rect 25596 9605 25605 9639
rect 25605 9605 25639 9639
rect 25639 9605 25648 9639
rect 25596 9596 25648 9605
rect 17592 9528 17644 9580
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 17776 9460 17828 9512
rect 13544 9392 13596 9444
rect 21456 9460 21508 9512
rect 20536 9392 20588 9444
rect 11152 9324 11204 9376
rect 12808 9324 12860 9376
rect 14556 9324 14608 9376
rect 16488 9324 16540 9376
rect 19800 9324 19852 9376
rect 27252 9528 27304 9580
rect 27436 9571 27488 9580
rect 27436 9537 27470 9571
rect 27470 9537 27488 9571
rect 27436 9528 27488 9537
rect 29000 9571 29052 9580
rect 29000 9537 29009 9571
rect 29009 9537 29043 9571
rect 29043 9537 29052 9571
rect 29000 9528 29052 9537
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 25044 9503 25096 9512
rect 25044 9469 25053 9503
rect 25053 9469 25087 9503
rect 25087 9469 25096 9503
rect 25044 9460 25096 9469
rect 25320 9460 25372 9512
rect 26240 9324 26292 9376
rect 26884 9324 26936 9376
rect 28540 9367 28592 9376
rect 28540 9333 28549 9367
rect 28549 9333 28583 9367
rect 28583 9333 28592 9367
rect 28540 9324 28592 9333
rect 29644 9639 29696 9648
rect 29644 9605 29653 9639
rect 29653 9605 29687 9639
rect 29687 9605 29696 9639
rect 29644 9596 29696 9605
rect 32036 9664 32088 9716
rect 31484 9596 31536 9648
rect 33140 9596 33192 9648
rect 36360 9596 36412 9648
rect 39028 9596 39080 9648
rect 30196 9528 30248 9580
rect 30288 9460 30340 9512
rect 32772 9503 32824 9512
rect 32772 9469 32781 9503
rect 32781 9469 32815 9503
rect 32815 9469 32824 9503
rect 32772 9460 32824 9469
rect 32864 9503 32916 9512
rect 32864 9469 32873 9503
rect 32873 9469 32907 9503
rect 32907 9469 32916 9503
rect 32864 9460 32916 9469
rect 32956 9460 33008 9512
rect 34520 9571 34572 9580
rect 34520 9537 34529 9571
rect 34529 9537 34563 9571
rect 34563 9537 34572 9571
rect 34520 9528 34572 9537
rect 34704 9460 34756 9512
rect 30564 9324 30616 9376
rect 31208 9324 31260 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 10784 9120 10836 9172
rect 16212 9120 16264 9172
rect 17776 9120 17828 9172
rect 19340 9120 19392 9172
rect 15660 9052 15712 9104
rect 17592 9052 17644 9104
rect 20812 9095 20864 9104
rect 20812 9061 20821 9095
rect 20821 9061 20855 9095
rect 20855 9061 20864 9095
rect 20812 9052 20864 9061
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 25320 9120 25372 9129
rect 30656 9120 30708 9172
rect 32864 9120 32916 9172
rect 36268 9120 36320 9172
rect 30564 9052 30616 9104
rect 32036 9052 32088 9104
rect 35624 9095 35676 9104
rect 35624 9061 35633 9095
rect 35633 9061 35667 9095
rect 35667 9061 35676 9095
rect 35624 9052 35676 9061
rect 17040 8984 17092 9036
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 16488 8959 16540 8968
rect 14372 8891 14424 8900
rect 14372 8857 14381 8891
rect 14381 8857 14415 8891
rect 14415 8857 14424 8891
rect 14372 8848 14424 8857
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 20076 8984 20128 9036
rect 21088 8984 21140 9036
rect 22008 8984 22060 9036
rect 27252 9027 27304 9036
rect 27252 8993 27261 9027
rect 27261 8993 27295 9027
rect 27295 8993 27304 9027
rect 27252 8984 27304 8993
rect 16028 8848 16080 8900
rect 18420 8848 18472 8900
rect 19156 8916 19208 8968
rect 19800 8959 19852 8968
rect 19800 8925 19809 8959
rect 19809 8925 19843 8959
rect 19843 8925 19852 8959
rect 19800 8916 19852 8925
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 24952 8959 25004 8968
rect 24952 8925 24961 8959
rect 24961 8925 24995 8959
rect 24995 8925 25004 8959
rect 24952 8916 25004 8925
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 26700 8959 26752 8968
rect 26700 8925 26709 8959
rect 26709 8925 26743 8959
rect 26743 8925 26752 8959
rect 26700 8916 26752 8925
rect 30196 8959 30248 8968
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 30472 8959 30524 8968
rect 30472 8925 30481 8959
rect 30481 8925 30515 8959
rect 30515 8925 30524 8959
rect 30472 8916 30524 8925
rect 33048 9027 33100 9036
rect 33048 8993 33057 9027
rect 33057 8993 33091 9027
rect 33091 8993 33100 9027
rect 33048 8984 33100 8993
rect 36268 9027 36320 9036
rect 36268 8993 36277 9027
rect 36277 8993 36311 9027
rect 36311 8993 36320 9027
rect 36268 8984 36320 8993
rect 17132 8780 17184 8832
rect 18972 8780 19024 8832
rect 22468 8848 22520 8900
rect 24308 8848 24360 8900
rect 26424 8848 26476 8900
rect 25412 8780 25464 8832
rect 29368 8848 29420 8900
rect 30748 8848 30800 8900
rect 30932 8959 30984 8968
rect 30932 8925 30941 8959
rect 30941 8925 30975 8959
rect 30975 8925 30984 8959
rect 30932 8916 30984 8925
rect 33784 8916 33836 8968
rect 35532 8959 35584 8968
rect 35532 8925 35541 8959
rect 35541 8925 35575 8959
rect 35575 8925 35584 8959
rect 35532 8916 35584 8925
rect 36360 8959 36412 8968
rect 36360 8925 36369 8959
rect 36369 8925 36403 8959
rect 36403 8925 36412 8959
rect 36360 8916 36412 8925
rect 31208 8891 31260 8900
rect 31208 8857 31242 8891
rect 31242 8857 31260 8891
rect 31208 8848 31260 8857
rect 37740 8848 37792 8900
rect 26884 8780 26936 8832
rect 28816 8780 28868 8832
rect 32956 8780 33008 8832
rect 34796 8780 34848 8832
rect 38108 8891 38160 8900
rect 38108 8857 38117 8891
rect 38117 8857 38151 8891
rect 38151 8857 38160 8891
rect 38108 8848 38160 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 11244 8576 11296 8628
rect 14648 8576 14700 8628
rect 13084 8508 13136 8560
rect 20904 8576 20956 8628
rect 25136 8576 25188 8628
rect 27436 8576 27488 8628
rect 28540 8576 28592 8628
rect 29828 8576 29880 8628
rect 34796 8576 34848 8628
rect 36268 8576 36320 8628
rect 37740 8576 37792 8628
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 19984 8551 20036 8560
rect 19984 8517 19993 8551
rect 19993 8517 20027 8551
rect 20027 8517 20036 8551
rect 19984 8508 20036 8517
rect 20076 8508 20128 8560
rect 23388 8508 23440 8560
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18420 8440 18472 8492
rect 18972 8440 19024 8492
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 24860 8440 24912 8492
rect 25044 8440 25096 8492
rect 18236 8372 18288 8424
rect 21272 8372 21324 8424
rect 24308 8415 24360 8424
rect 13728 8304 13780 8356
rect 16488 8304 16540 8356
rect 20720 8304 20772 8356
rect 15660 8236 15712 8288
rect 21548 8236 21600 8288
rect 24308 8381 24317 8415
rect 24317 8381 24351 8415
rect 24351 8381 24360 8415
rect 24308 8372 24360 8381
rect 27620 8440 27672 8492
rect 30196 8508 30248 8560
rect 31300 8551 31352 8560
rect 31300 8517 31309 8551
rect 31309 8517 31343 8551
rect 31343 8517 31352 8551
rect 31300 8508 31352 8517
rect 33784 8551 33836 8560
rect 33784 8517 33793 8551
rect 33793 8517 33827 8551
rect 33827 8517 33836 8551
rect 33784 8508 33836 8517
rect 29368 8440 29420 8492
rect 30472 8483 30524 8492
rect 30472 8449 30481 8483
rect 30481 8449 30515 8483
rect 30515 8449 30524 8483
rect 30472 8440 30524 8449
rect 30748 8483 30800 8492
rect 30748 8449 30757 8483
rect 30757 8449 30791 8483
rect 30791 8449 30800 8483
rect 30748 8440 30800 8449
rect 32956 8440 33008 8492
rect 36820 8508 36872 8560
rect 35256 8483 35308 8492
rect 35256 8449 35290 8483
rect 35290 8449 35308 8483
rect 35256 8440 35308 8449
rect 28264 8372 28316 8424
rect 34244 8372 34296 8424
rect 35992 8372 36044 8424
rect 38016 8415 38068 8424
rect 38016 8381 38025 8415
rect 38025 8381 38059 8415
rect 38059 8381 38068 8415
rect 38016 8372 38068 8381
rect 29460 8347 29512 8356
rect 29460 8313 29469 8347
rect 29469 8313 29503 8347
rect 29503 8313 29512 8347
rect 29460 8304 29512 8313
rect 32128 8304 32180 8356
rect 37188 8304 37240 8356
rect 27804 8236 27856 8288
rect 33048 8236 33100 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 15476 8032 15528 8084
rect 16028 8032 16080 8084
rect 14096 7964 14148 8016
rect 11060 7896 11112 7948
rect 22928 8075 22980 8084
rect 22928 8041 22937 8075
rect 22937 8041 22971 8075
rect 22971 8041 22980 8075
rect 22928 8032 22980 8041
rect 24860 8075 24912 8084
rect 24860 8041 24869 8075
rect 24869 8041 24903 8075
rect 24903 8041 24912 8075
rect 24860 8032 24912 8041
rect 29000 8032 29052 8084
rect 23204 7964 23256 8016
rect 25228 7964 25280 8016
rect 11152 7828 11204 7880
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 14188 7828 14240 7880
rect 14372 7828 14424 7880
rect 15476 7828 15528 7880
rect 17960 7760 18012 7812
rect 18512 7828 18564 7880
rect 20996 7896 21048 7948
rect 25504 7939 25556 7948
rect 25504 7905 25513 7939
rect 25513 7905 25547 7939
rect 25547 7905 25556 7939
rect 25504 7896 25556 7905
rect 29092 7896 29144 7948
rect 31208 8032 31260 8084
rect 32404 8032 32456 8084
rect 33048 7964 33100 8016
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 21088 7828 21140 7880
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 25136 7828 25188 7880
rect 26424 7871 26476 7880
rect 26424 7837 26433 7871
rect 26433 7837 26467 7871
rect 26467 7837 26476 7871
rect 26424 7828 26476 7837
rect 28264 7871 28316 7880
rect 28264 7837 28273 7871
rect 28273 7837 28307 7871
rect 28307 7837 28316 7871
rect 28264 7828 28316 7837
rect 30196 7871 30248 7880
rect 30196 7837 30205 7871
rect 30205 7837 30239 7871
rect 30239 7837 30248 7871
rect 30196 7828 30248 7837
rect 30932 7828 30984 7880
rect 32956 7828 33008 7880
rect 33876 8075 33928 8084
rect 33876 8041 33885 8075
rect 33885 8041 33919 8075
rect 33919 8041 33928 8075
rect 33876 8032 33928 8041
rect 35348 8032 35400 8084
rect 37832 8032 37884 8084
rect 35992 7964 36044 8016
rect 35808 7939 35860 7948
rect 35808 7905 35817 7939
rect 35817 7905 35851 7939
rect 35851 7905 35860 7939
rect 35808 7896 35860 7905
rect 34244 7871 34296 7880
rect 34244 7837 34253 7871
rect 34253 7837 34287 7871
rect 34287 7837 34296 7871
rect 34244 7828 34296 7837
rect 36268 7828 36320 7880
rect 36820 7828 36872 7880
rect 37188 7871 37240 7880
rect 37188 7837 37222 7871
rect 37222 7837 37240 7871
rect 37188 7828 37240 7837
rect 18972 7760 19024 7812
rect 22008 7760 22060 7812
rect 27160 7760 27212 7812
rect 19432 7692 19484 7744
rect 27528 7692 27580 7744
rect 32772 7760 32824 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12808 7420 12860 7472
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 22008 7531 22060 7540
rect 22008 7497 22017 7531
rect 22017 7497 22051 7531
rect 22051 7497 22060 7531
rect 22008 7488 22060 7497
rect 23756 7488 23808 7540
rect 24768 7488 24820 7540
rect 26240 7488 26292 7540
rect 27160 7531 27212 7540
rect 27160 7497 27169 7531
rect 27169 7497 27203 7531
rect 27203 7497 27212 7531
rect 27160 7488 27212 7497
rect 27528 7531 27580 7540
rect 27528 7497 27537 7531
rect 27537 7497 27571 7531
rect 27571 7497 27580 7531
rect 27528 7488 27580 7497
rect 28908 7488 28960 7540
rect 18420 7420 18472 7472
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14740 7352 14792 7404
rect 15660 7395 15712 7404
rect 15660 7361 15668 7395
rect 15668 7361 15702 7395
rect 15702 7361 15712 7395
rect 15660 7352 15712 7361
rect 16488 7352 16540 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 18972 7420 19024 7472
rect 23940 7463 23992 7472
rect 23940 7429 23949 7463
rect 23949 7429 23983 7463
rect 23983 7429 23992 7463
rect 23940 7420 23992 7429
rect 27436 7420 27488 7472
rect 33140 7420 33192 7472
rect 35716 7420 35768 7472
rect 13084 7284 13136 7336
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 18328 7284 18380 7336
rect 20812 7352 20864 7404
rect 20904 7284 20956 7336
rect 19248 7259 19300 7268
rect 19248 7225 19257 7259
rect 19257 7225 19291 7259
rect 19291 7225 19300 7259
rect 19248 7216 19300 7225
rect 22100 7352 22152 7404
rect 32772 7352 32824 7404
rect 34704 7395 34756 7404
rect 34704 7361 34713 7395
rect 34713 7361 34747 7395
rect 34747 7361 34756 7395
rect 34704 7352 34756 7361
rect 34796 7352 34848 7404
rect 25504 7284 25556 7336
rect 25872 7284 25924 7336
rect 27804 7327 27856 7336
rect 27804 7293 27813 7327
rect 27813 7293 27847 7327
rect 27847 7293 27856 7327
rect 27804 7284 27856 7293
rect 34612 7284 34664 7336
rect 37740 7352 37792 7404
rect 38108 7327 38160 7336
rect 38108 7293 38117 7327
rect 38117 7293 38151 7327
rect 38151 7293 38160 7327
rect 38108 7284 38160 7293
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 20352 7148 20404 7200
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 24308 7191 24360 7200
rect 24308 7157 24317 7191
rect 24317 7157 24351 7191
rect 24351 7157 24360 7191
rect 24308 7148 24360 7157
rect 34060 7191 34112 7200
rect 34060 7157 34069 7191
rect 34069 7157 34103 7191
rect 34103 7157 34112 7191
rect 34060 7148 34112 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12900 6944 12952 6996
rect 18236 6987 18288 6996
rect 18236 6953 18245 6987
rect 18245 6953 18279 6987
rect 18279 6953 18288 6987
rect 18236 6944 18288 6953
rect 18512 6944 18564 6996
rect 20352 6944 20404 6996
rect 23940 6944 23992 6996
rect 26332 6944 26384 6996
rect 33140 6987 33192 6996
rect 33140 6953 33149 6987
rect 33149 6953 33183 6987
rect 33183 6953 33192 6987
rect 33140 6944 33192 6953
rect 37740 6944 37792 6996
rect 13728 6876 13780 6928
rect 14004 6740 14056 6792
rect 14648 6808 14700 6860
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 17960 6808 18012 6860
rect 15476 6740 15528 6792
rect 15936 6740 15988 6792
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 18420 6808 18472 6860
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 20628 6783 20680 6792
rect 20628 6749 20637 6783
rect 20637 6749 20671 6783
rect 20671 6749 20680 6783
rect 20628 6740 20680 6749
rect 21548 6740 21600 6792
rect 22192 6740 22244 6792
rect 24124 6808 24176 6860
rect 24952 6808 25004 6860
rect 25412 6808 25464 6860
rect 26056 6740 26108 6792
rect 28264 6808 28316 6860
rect 28816 6808 28868 6860
rect 29460 6808 29512 6860
rect 29552 6808 29604 6860
rect 21088 6672 21140 6724
rect 21272 6715 21324 6724
rect 21272 6681 21281 6715
rect 21281 6681 21315 6715
rect 21315 6681 21324 6715
rect 21272 6672 21324 6681
rect 21456 6647 21508 6656
rect 21456 6613 21481 6647
rect 21481 6613 21508 6647
rect 21456 6604 21508 6613
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 23204 6672 23256 6724
rect 25320 6672 25372 6724
rect 23756 6604 23808 6656
rect 25412 6604 25464 6656
rect 26148 6715 26200 6724
rect 26148 6681 26157 6715
rect 26157 6681 26191 6715
rect 26191 6681 26200 6715
rect 26148 6672 26200 6681
rect 26240 6672 26292 6724
rect 29276 6740 29328 6792
rect 30564 6808 30616 6860
rect 33140 6808 33192 6860
rect 30380 6783 30432 6792
rect 30380 6749 30389 6783
rect 30389 6749 30423 6783
rect 30423 6749 30432 6783
rect 30380 6740 30432 6749
rect 29920 6672 29972 6724
rect 36820 6740 36872 6792
rect 34060 6672 34112 6724
rect 37464 6672 37516 6724
rect 28816 6604 28868 6656
rect 37924 6604 37976 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 20628 6400 20680 6452
rect 19340 6332 19392 6384
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 18328 6264 18380 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 16212 6239 16264 6248
rect 16212 6205 16221 6239
rect 16221 6205 16255 6239
rect 16255 6205 16264 6239
rect 16212 6196 16264 6205
rect 19156 6196 19208 6248
rect 21456 6332 21508 6384
rect 22100 6332 22152 6384
rect 23204 6443 23256 6452
rect 23204 6409 23213 6443
rect 23213 6409 23247 6443
rect 23247 6409 23256 6443
rect 23204 6400 23256 6409
rect 23940 6400 23992 6452
rect 26148 6400 26200 6452
rect 28264 6400 28316 6452
rect 29920 6443 29972 6452
rect 29920 6409 29929 6443
rect 29929 6409 29963 6443
rect 29963 6409 29972 6443
rect 29920 6400 29972 6409
rect 30380 6443 30432 6452
rect 30380 6409 30389 6443
rect 30389 6409 30423 6443
rect 30423 6409 30432 6443
rect 30380 6400 30432 6409
rect 24124 6332 24176 6384
rect 24308 6332 24360 6384
rect 24952 6332 25004 6384
rect 20352 6307 20404 6316
rect 20352 6273 20361 6307
rect 20361 6273 20395 6307
rect 20395 6273 20404 6307
rect 20352 6264 20404 6273
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21640 6264 21692 6316
rect 24216 6264 24268 6316
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 25320 6264 25372 6316
rect 14740 6128 14792 6180
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 26148 6307 26200 6316
rect 26148 6273 26157 6307
rect 26157 6273 26191 6307
rect 26191 6273 26200 6307
rect 26148 6264 26200 6273
rect 26240 6307 26292 6316
rect 26240 6273 26249 6307
rect 26249 6273 26283 6307
rect 26283 6273 26292 6307
rect 26240 6264 26292 6273
rect 26424 6264 26476 6316
rect 27252 6264 27304 6316
rect 27896 6264 27948 6316
rect 28632 6264 28684 6316
rect 26056 6196 26108 6248
rect 29276 6196 29328 6248
rect 34060 6332 34112 6384
rect 34704 6400 34756 6452
rect 35440 6443 35492 6452
rect 35440 6409 35449 6443
rect 35449 6409 35483 6443
rect 35483 6409 35492 6443
rect 35440 6400 35492 6409
rect 37464 6443 37516 6452
rect 37464 6409 37473 6443
rect 37473 6409 37507 6443
rect 37507 6409 37516 6443
rect 37464 6400 37516 6409
rect 37740 6400 37792 6452
rect 37924 6443 37976 6452
rect 37924 6409 37933 6443
rect 37933 6409 37967 6443
rect 37967 6409 37976 6443
rect 37924 6400 37976 6409
rect 34520 6332 34572 6384
rect 30748 6307 30800 6316
rect 30748 6273 30757 6307
rect 30757 6273 30791 6307
rect 30791 6273 30800 6307
rect 30748 6264 30800 6273
rect 34244 6264 34296 6316
rect 34796 6307 34848 6316
rect 34796 6273 34805 6307
rect 34805 6273 34839 6307
rect 34839 6273 34848 6307
rect 34796 6264 34848 6273
rect 34888 6264 34940 6316
rect 30840 6239 30892 6248
rect 30840 6205 30849 6239
rect 30849 6205 30883 6239
rect 30883 6205 30892 6239
rect 30840 6196 30892 6205
rect 20996 6060 21048 6112
rect 25504 6060 25556 6112
rect 29460 6128 29512 6180
rect 34612 6196 34664 6248
rect 37740 6264 37792 6316
rect 38016 6239 38068 6248
rect 38016 6205 38025 6239
rect 38025 6205 38059 6239
rect 38059 6205 38068 6239
rect 38016 6196 38068 6205
rect 28448 6060 28500 6112
rect 30012 6060 30064 6112
rect 37832 6060 37884 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 18052 5856 18104 5908
rect 19248 5856 19300 5908
rect 16212 5720 16264 5772
rect 16488 5720 16540 5772
rect 19340 5788 19392 5840
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 25320 5899 25372 5908
rect 25320 5865 25329 5899
rect 25329 5865 25363 5899
rect 25363 5865 25372 5899
rect 25320 5856 25372 5865
rect 25412 5899 25464 5908
rect 25412 5865 25421 5899
rect 25421 5865 25455 5899
rect 25455 5865 25464 5899
rect 25412 5856 25464 5865
rect 27896 5899 27948 5908
rect 27896 5865 27905 5899
rect 27905 5865 27939 5899
rect 27939 5865 27948 5899
rect 27896 5856 27948 5865
rect 30564 5856 30616 5908
rect 18052 5720 18104 5772
rect 19156 5720 19208 5772
rect 19432 5720 19484 5772
rect 20720 5763 20772 5772
rect 20720 5729 20729 5763
rect 20729 5729 20763 5763
rect 20763 5729 20772 5763
rect 20720 5720 20772 5729
rect 22192 5720 22244 5772
rect 25504 5763 25556 5772
rect 25504 5729 25513 5763
rect 25513 5729 25547 5763
rect 25547 5729 25556 5763
rect 25504 5720 25556 5729
rect 28172 5720 28224 5772
rect 28448 5763 28500 5772
rect 28448 5729 28457 5763
rect 28457 5729 28491 5763
rect 28491 5729 28500 5763
rect 28448 5720 28500 5729
rect 32404 5720 32456 5772
rect 33140 5763 33192 5772
rect 33140 5729 33149 5763
rect 33149 5729 33183 5763
rect 33183 5729 33192 5763
rect 33140 5720 33192 5729
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 25228 5695 25280 5704
rect 25228 5661 25237 5695
rect 25237 5661 25271 5695
rect 25271 5661 25280 5695
rect 25228 5652 25280 5661
rect 28264 5695 28316 5704
rect 28264 5661 28273 5695
rect 28273 5661 28307 5695
rect 28307 5661 28316 5695
rect 28264 5652 28316 5661
rect 29736 5652 29788 5704
rect 31760 5652 31812 5704
rect 33692 5652 33744 5704
rect 35532 5899 35584 5908
rect 35532 5865 35541 5899
rect 35541 5865 35575 5899
rect 35575 5865 35584 5899
rect 35532 5856 35584 5865
rect 30472 5627 30524 5636
rect 30472 5593 30506 5627
rect 30506 5593 30524 5627
rect 30472 5584 30524 5593
rect 34244 5584 34296 5636
rect 34520 5584 34572 5636
rect 36452 5652 36504 5704
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 38108 5627 38160 5636
rect 38108 5593 38117 5627
rect 38117 5593 38151 5627
rect 38151 5593 38160 5627
rect 38108 5584 38160 5593
rect 19432 5559 19484 5568
rect 19432 5525 19441 5559
rect 19441 5525 19475 5559
rect 19475 5525 19484 5559
rect 19432 5516 19484 5525
rect 30748 5516 30800 5568
rect 32588 5559 32640 5568
rect 32588 5525 32597 5559
rect 32597 5525 32631 5559
rect 32631 5525 32640 5559
rect 32588 5516 32640 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 23572 5355 23624 5364
rect 23572 5321 23581 5355
rect 23581 5321 23615 5355
rect 23615 5321 23624 5355
rect 23572 5312 23624 5321
rect 24584 5312 24636 5364
rect 30472 5312 30524 5364
rect 30748 5355 30800 5364
rect 30748 5321 30757 5355
rect 30757 5321 30791 5355
rect 30791 5321 30800 5355
rect 30748 5312 30800 5321
rect 33692 5355 33744 5364
rect 33692 5321 33701 5355
rect 33701 5321 33735 5355
rect 33735 5321 33744 5355
rect 33692 5312 33744 5321
rect 34796 5312 34848 5364
rect 36452 5355 36504 5364
rect 36452 5321 36461 5355
rect 36461 5321 36495 5355
rect 36495 5321 36504 5355
rect 36452 5312 36504 5321
rect 37740 5312 37792 5364
rect 16672 5244 16724 5296
rect 23480 5244 23532 5296
rect 31760 5244 31812 5296
rect 20720 5176 20772 5228
rect 23020 5176 23072 5228
rect 25228 5176 25280 5228
rect 25964 5176 26016 5228
rect 28172 5176 28224 5228
rect 30564 5176 30616 5228
rect 32956 5244 33008 5296
rect 34244 5244 34296 5296
rect 32588 5219 32640 5228
rect 32588 5185 32622 5219
rect 32622 5185 32640 5219
rect 32588 5176 32640 5185
rect 34336 5219 34388 5228
rect 34336 5185 34345 5219
rect 34345 5185 34379 5219
rect 34379 5185 34388 5219
rect 34336 5176 34388 5185
rect 36820 5244 36872 5296
rect 37648 5244 37700 5296
rect 35348 5219 35400 5228
rect 35348 5185 35382 5219
rect 35382 5185 35400 5219
rect 35348 5176 35400 5185
rect 19432 5108 19484 5160
rect 19524 5151 19576 5160
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 19524 5108 19576 5117
rect 22192 5151 22244 5160
rect 22192 5117 22201 5151
rect 22201 5117 22235 5151
rect 22235 5117 22244 5151
rect 22192 5108 22244 5117
rect 24952 5151 25004 5160
rect 24952 5117 24961 5151
rect 24961 5117 24995 5151
rect 24995 5117 25004 5151
rect 24952 5108 25004 5117
rect 25044 5151 25096 5160
rect 25044 5117 25053 5151
rect 25053 5117 25087 5151
rect 25087 5117 25096 5151
rect 25044 5108 25096 5117
rect 30656 5108 30708 5160
rect 31208 5108 31260 5160
rect 38016 5151 38068 5160
rect 38016 5117 38025 5151
rect 38025 5117 38059 5151
rect 38059 5117 38068 5151
rect 38016 5108 38068 5117
rect 37556 5040 37608 5092
rect 24676 4972 24728 5024
rect 37464 5015 37516 5024
rect 37464 4981 37473 5015
rect 37473 4981 37507 5015
rect 37507 4981 37516 5015
rect 37464 4972 37516 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20076 4768 20128 4820
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 11060 4632 11112 4684
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 25964 4743 26016 4752
rect 25964 4709 25973 4743
rect 25973 4709 26007 4743
rect 26007 4709 26016 4743
rect 25964 4700 26016 4709
rect 26056 4700 26108 4752
rect 28172 4632 28224 4684
rect 30840 4768 30892 4820
rect 31208 4768 31260 4820
rect 29184 4632 29236 4684
rect 29736 4675 29788 4684
rect 29736 4641 29745 4675
rect 29745 4641 29779 4675
rect 29779 4641 29788 4675
rect 29736 4632 29788 4641
rect 32956 4675 33008 4684
rect 32956 4641 32965 4675
rect 32965 4641 32999 4675
rect 32999 4641 33008 4675
rect 32956 4632 33008 4641
rect 34336 4811 34388 4820
rect 34336 4777 34345 4811
rect 34345 4777 34379 4811
rect 34379 4777 34388 4811
rect 34336 4768 34388 4777
rect 35348 4768 35400 4820
rect 37556 4768 37608 4820
rect 37740 4768 37792 4820
rect 36820 4675 36872 4684
rect 36820 4641 36829 4675
rect 36829 4641 36863 4675
rect 36863 4641 36872 4675
rect 36820 4632 36872 4641
rect 22192 4564 22244 4616
rect 24676 4564 24728 4616
rect 27252 4564 27304 4616
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 36452 4564 36504 4616
rect 37464 4564 37516 4616
rect 23572 4496 23624 4548
rect 26516 4496 26568 4548
rect 30104 4496 30156 4548
rect 33416 4496 33468 4548
rect 35992 4539 36044 4548
rect 35992 4505 36001 4539
rect 36001 4505 36035 4539
rect 36035 4505 36044 4539
rect 35992 4496 36044 4505
rect 23664 4428 23716 4480
rect 24952 4428 25004 4480
rect 28264 4471 28316 4480
rect 28264 4437 28273 4471
rect 28273 4437 28307 4471
rect 28307 4437 28316 4471
rect 28264 4428 28316 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 26056 4224 26108 4276
rect 26516 4267 26568 4276
rect 26516 4233 26525 4267
rect 26525 4233 26559 4267
rect 26559 4233 26568 4267
rect 26516 4224 26568 4233
rect 28632 4224 28684 4276
rect 30104 4267 30156 4276
rect 30104 4233 30113 4267
rect 30113 4233 30147 4267
rect 30147 4233 30156 4267
rect 30104 4224 30156 4233
rect 30840 4224 30892 4276
rect 33416 4267 33468 4276
rect 33416 4233 33425 4267
rect 33425 4233 33459 4267
rect 33459 4233 33468 4267
rect 33416 4224 33468 4233
rect 34336 4224 34388 4276
rect 28264 4156 28316 4208
rect 30564 4199 30616 4208
rect 30564 4165 30573 4199
rect 30573 4165 30607 4199
rect 30607 4165 30616 4199
rect 30564 4156 30616 4165
rect 24952 4088 25004 4140
rect 27252 4088 27304 4140
rect 33876 4131 33928 4140
rect 33876 4097 33885 4131
rect 33885 4097 33919 4131
rect 33919 4097 33928 4131
rect 33876 4088 33928 4097
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 33140 3952 33192 4004
rect 29644 3884 29696 3936
rect 39028 4088 39080 4140
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 37832 3043 37884 3052
rect 37832 3009 37841 3043
rect 37841 3009 37875 3043
rect 37875 3009 37884 3043
rect 37832 3000 37884 3009
rect 38108 2975 38160 2984
rect 38108 2941 38117 2975
rect 38117 2941 38151 2975
rect 38151 2941 38160 2975
rect 38108 2932 38160 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 28080 2388 28132 2440
rect 38108 2363 38160 2372
rect 38108 2329 38117 2363
rect 38117 2329 38151 2363
rect 38151 2329 38160 2363
rect 38108 2320 38160 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1766 39200 1822 40000
rect 5078 39200 5134 40000
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 38198 39200 38254 40000
rect 1780 37262 1808 39200
rect 5092 39166 5120 39200
rect 5080 39160 5132 39166
rect 5080 39102 5132 39108
rect 6644 39160 6696 39166
rect 6644 39102 6696 39108
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5816 37324 5868 37330
rect 5816 37266 5868 37272
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5172 37120 5224 37126
rect 5172 37062 5224 37068
rect 5184 36854 5212 37062
rect 5172 36848 5224 36854
rect 5172 36790 5224 36796
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 36654
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 34746 4660 36110
rect 5552 36106 5580 37130
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5644 36922 5672 37062
rect 5632 36916 5684 36922
rect 5632 36858 5684 36864
rect 5644 36242 5672 36858
rect 5632 36236 5684 36242
rect 5632 36178 5684 36184
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5264 36032 5316 36038
rect 5552 36009 5580 36042
rect 5264 35974 5316 35980
rect 5538 36000 5594 36009
rect 5172 34944 5224 34950
rect 5172 34886 5224 34892
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 5184 34610 5212 34886
rect 5172 34604 5224 34610
rect 5172 34546 5224 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4988 33108 5040 33114
rect 4988 33050 5040 33056
rect 4528 32904 4580 32910
rect 4528 32846 4580 32852
rect 4540 32434 4568 32846
rect 5000 32434 5028 33050
rect 5276 32910 5304 35974
rect 5538 35935 5594 35944
rect 5828 35630 5856 37266
rect 6656 37262 6684 39102
rect 8404 37262 8432 39200
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 6644 37256 6696 37262
rect 6644 37198 6696 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 7380 37188 7432 37194
rect 7380 37130 7432 37136
rect 5908 36236 5960 36242
rect 5908 36178 5960 36184
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5828 35154 5856 35566
rect 5816 35148 5868 35154
rect 5816 35090 5868 35096
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5644 34746 5672 34886
rect 5632 34740 5684 34746
rect 5632 34682 5684 34688
rect 5540 34672 5592 34678
rect 5540 34614 5592 34620
rect 5552 34066 5580 34614
rect 5644 34066 5672 34682
rect 5920 34678 5948 36178
rect 7024 35018 7052 37130
rect 7104 36100 7156 36106
rect 7104 36042 7156 36048
rect 7116 35834 7144 36042
rect 7392 35894 7420 37130
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9140 36854 9168 37062
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 9140 36174 9168 36518
rect 9220 36304 9272 36310
rect 9220 36246 9272 36252
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 7840 36032 7892 36038
rect 7840 35974 7892 35980
rect 7392 35866 7512 35894
rect 7104 35828 7156 35834
rect 7104 35770 7156 35776
rect 7484 35698 7512 35866
rect 7852 35834 7880 35974
rect 7564 35828 7616 35834
rect 7564 35770 7616 35776
rect 7840 35828 7892 35834
rect 7840 35770 7892 35776
rect 7472 35692 7524 35698
rect 7472 35634 7524 35640
rect 6368 35012 6420 35018
rect 6368 34954 6420 34960
rect 7012 35012 7064 35018
rect 7012 34954 7064 34960
rect 5908 34672 5960 34678
rect 5908 34614 5960 34620
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5632 34060 5684 34066
rect 5632 34002 5684 34008
rect 6380 33930 6408 34954
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 6368 33924 6420 33930
rect 6368 33866 6420 33872
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 6000 33448 6052 33454
rect 6000 33390 6052 33396
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 4528 32428 4580 32434
rect 4528 32370 4580 32376
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3424 31952 3476 31958
rect 3424 31894 3476 31900
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2792 26994 2820 30194
rect 3436 29714 3464 31894
rect 4068 31680 4120 31686
rect 4068 31622 4120 31628
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 3988 29850 4016 30194
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 3424 29708 3476 29714
rect 3424 29650 3476 29656
rect 3148 29640 3200 29646
rect 3148 29582 3200 29588
rect 3332 29640 3384 29646
rect 3332 29582 3384 29588
rect 3160 29170 3188 29582
rect 3344 29238 3372 29582
rect 3332 29232 3384 29238
rect 3332 29174 3384 29180
rect 3976 29232 4028 29238
rect 3976 29174 4028 29180
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3988 28762 4016 29174
rect 3976 28756 4028 28762
rect 3976 28698 4028 28704
rect 3884 28008 3936 28014
rect 3884 27950 3936 27956
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 2792 24818 2820 26930
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2792 23730 2820 24754
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 3896 23254 3924 27950
rect 3976 27328 4028 27334
rect 3976 27270 4028 27276
rect 3988 27062 4016 27270
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3988 24886 4016 25094
rect 3976 24880 4028 24886
rect 3976 24822 4028 24828
rect 4080 23798 4108 31622
rect 4908 31346 4936 32166
rect 5000 31754 5028 32370
rect 5644 32298 5672 33254
rect 6012 32978 6040 33390
rect 6000 32972 6052 32978
rect 6000 32914 6052 32920
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5632 32292 5684 32298
rect 5632 32234 5684 32240
rect 4988 31748 5040 31754
rect 4988 31690 5040 31696
rect 5000 31346 5028 31690
rect 5644 31482 5672 32234
rect 5724 32224 5776 32230
rect 5724 32166 5776 32172
rect 5736 32026 5764 32166
rect 5724 32020 5776 32026
rect 5724 31962 5776 31968
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4804 30864 4856 30870
rect 4804 30806 4856 30812
rect 4816 30258 4844 30806
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4908 30190 4936 31282
rect 5264 30932 5316 30938
rect 5264 30874 5316 30880
rect 5276 30666 5304 30874
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 4988 30592 5040 30598
rect 4988 30534 5040 30540
rect 4896 30184 4948 30190
rect 4896 30126 4948 30132
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29510 4660 29990
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4816 29238 4844 29990
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27606 4660 28970
rect 4908 28778 4936 29106
rect 5000 28937 5028 30534
rect 5080 30252 5132 30258
rect 5080 30194 5132 30200
rect 5092 29510 5120 30194
rect 5080 29504 5132 29510
rect 5080 29446 5132 29452
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5080 29028 5132 29034
rect 5080 28970 5132 28976
rect 4986 28928 5042 28937
rect 4986 28863 5042 28872
rect 4816 28750 4936 28778
rect 4988 28756 5040 28762
rect 4816 28218 4844 28750
rect 4988 28698 5040 28704
rect 4894 28656 4950 28665
rect 4894 28591 4950 28600
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 4804 27872 4856 27878
rect 4710 27840 4766 27849
rect 4804 27814 4856 27820
rect 4710 27775 4766 27784
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4448 27130 4476 27406
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4724 26874 4752 27775
rect 4816 27402 4844 27814
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 4816 26994 4844 27338
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4724 26846 4844 26874
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25362 4660 26182
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4632 24614 4660 25162
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24138 4660 24550
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 3988 23322 4016 23666
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3884 23248 3936 23254
rect 3884 23190 3936 23196
rect 4632 23118 4660 23462
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 3988 21622 4016 21830
rect 4356 21690 4384 21830
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4632 21486 4660 22034
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 3068 20942 3096 21422
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19922 4660 21422
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4080 19446 4108 19654
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3436 18766 3464 19314
rect 4448 19242 4476 19654
rect 4632 19378 4660 19858
rect 4724 19854 4752 26726
rect 4816 25906 4844 26846
rect 4908 26382 4936 28591
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4908 26042 4936 26318
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25362 4936 25638
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 5000 24682 5028 28698
rect 5092 27470 5120 28970
rect 5184 28082 5212 29038
rect 5172 28076 5224 28082
rect 5172 28018 5224 28024
rect 5276 27962 5304 29106
rect 5460 29102 5488 31282
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5552 30258 5580 31214
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30598 5672 31078
rect 5632 30592 5684 30598
rect 5632 30534 5684 30540
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 5368 28762 5396 28902
rect 5356 28756 5408 28762
rect 5356 28698 5408 28704
rect 5460 28558 5488 29038
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5184 27934 5304 27962
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 5080 27328 5132 27334
rect 5080 27270 5132 27276
rect 5092 25430 5120 27270
rect 5184 25838 5212 27934
rect 5368 27538 5396 28358
rect 5552 28082 5580 30194
rect 5644 29646 5672 30534
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5644 27849 5672 29446
rect 5630 27840 5686 27849
rect 5630 27775 5686 27784
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5460 27112 5488 27406
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5276 27084 5488 27112
rect 5276 25974 5304 27084
rect 5552 27062 5580 27270
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5356 26988 5408 26994
rect 5356 26930 5408 26936
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 4988 24676 5040 24682
rect 4988 24618 5040 24624
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4816 22030 4844 23666
rect 4908 23050 4936 23802
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 5000 22710 5028 23666
rect 5092 23186 5120 25366
rect 5276 25362 5304 25910
rect 5368 25362 5396 26930
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5172 24744 5224 24750
rect 5172 24686 5224 24692
rect 5184 24410 5212 24686
rect 5172 24404 5224 24410
rect 5172 24346 5224 24352
rect 5368 24274 5396 25298
rect 5460 24750 5488 26386
rect 5644 26382 5672 27542
rect 5736 27470 5764 31962
rect 5828 31822 5856 32370
rect 6104 32366 6132 33798
rect 6184 32836 6236 32842
rect 6184 32778 6236 32784
rect 6092 32360 6144 32366
rect 6092 32302 6144 32308
rect 6196 31906 6224 32778
rect 6104 31890 6224 31906
rect 6092 31884 6224 31890
rect 6144 31878 6224 31884
rect 6092 31826 6144 31832
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 6196 31754 6224 31878
rect 6196 31726 6316 31754
rect 6000 31476 6052 31482
rect 6000 31418 6052 31424
rect 5816 31340 5868 31346
rect 5816 31282 5868 31288
rect 5828 30870 5856 31282
rect 5816 30864 5868 30870
rect 5816 30806 5868 30812
rect 5828 30734 5856 30806
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 5908 30660 5960 30666
rect 5908 30602 5960 30608
rect 5920 30394 5948 30602
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 6012 30274 6040 31418
rect 6092 31340 6144 31346
rect 6092 31282 6144 31288
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 5920 30246 6040 30274
rect 5828 29306 5856 30194
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 5920 28966 5948 30246
rect 6104 30054 6132 31282
rect 6000 30048 6052 30054
rect 6000 29990 6052 29996
rect 6092 30048 6144 30054
rect 6092 29990 6144 29996
rect 6012 29782 6040 29990
rect 6000 29776 6052 29782
rect 6000 29718 6052 29724
rect 6000 29164 6052 29170
rect 6000 29106 6052 29112
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 5816 28416 5868 28422
rect 5816 28358 5868 28364
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5552 25242 5580 25842
rect 5644 25498 5672 26318
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5736 25786 5764 26250
rect 5828 25906 5856 28358
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 5920 26994 5948 27270
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 6012 26874 6040 29106
rect 6288 27402 6316 31726
rect 6184 27396 6236 27402
rect 6184 27338 6236 27344
rect 6276 27396 6328 27402
rect 6276 27338 6328 27344
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5920 26846 6040 26874
rect 5920 26382 5948 26846
rect 6104 26382 6132 26930
rect 6196 26926 6224 27338
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5920 25838 5948 26318
rect 6196 26314 6224 26862
rect 6184 26308 6236 26314
rect 6184 26250 6236 26256
rect 6196 26194 6224 26250
rect 6104 26166 6224 26194
rect 5908 25832 5960 25838
rect 5736 25770 5856 25786
rect 5908 25774 5960 25780
rect 5736 25764 5868 25770
rect 5736 25758 5816 25764
rect 5816 25706 5868 25712
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5552 25214 5672 25242
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5552 24886 5580 25094
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5552 23798 5580 24822
rect 5644 24818 5672 25214
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5724 24336 5776 24342
rect 5724 24278 5776 24284
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5540 23792 5592 23798
rect 5540 23734 5592 23740
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5184 23322 5212 23666
rect 5644 23322 5672 24210
rect 5736 24206 5764 24278
rect 5828 24206 5856 25706
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 4988 22704 5040 22710
rect 4988 22646 5040 22652
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 5644 21962 5672 22578
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5736 21554 5764 23054
rect 5828 22778 5856 24142
rect 5920 23798 5948 25774
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 6012 23798 6040 24346
rect 5908 23792 5960 23798
rect 5908 23734 5960 23740
rect 6000 23792 6052 23798
rect 6000 23734 6052 23740
rect 5816 22772 5868 22778
rect 5816 22714 5868 22720
rect 6012 22642 6040 23734
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 20754 5488 20878
rect 5460 20726 5580 20754
rect 5552 20534 5580 20726
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 5644 19514 5672 19926
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4436 19236 4488 19242
rect 4436 19178 4488 19184
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 5276 18698 5304 19110
rect 5460 18902 5488 19178
rect 5644 18970 5672 19450
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 6104 18766 6132 26166
rect 6184 24064 6236 24070
rect 6184 24006 6236 24012
rect 6196 21554 6224 24006
rect 6288 23050 6316 27338
rect 6380 26518 6408 33866
rect 7116 33590 7144 34682
rect 7484 34542 7512 35634
rect 7576 34610 7604 35770
rect 9140 35086 9168 36110
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 7564 34604 7616 34610
rect 7564 34546 7616 34552
rect 7472 34536 7524 34542
rect 7472 34478 7524 34484
rect 7932 34536 7984 34542
rect 7932 34478 7984 34484
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 7380 33992 7432 33998
rect 7380 33934 7432 33940
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 7104 33584 7156 33590
rect 7104 33526 7156 33532
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 6564 33318 6592 33458
rect 6828 33448 6880 33454
rect 6828 33390 6880 33396
rect 6552 33312 6604 33318
rect 6552 33254 6604 33260
rect 6564 32910 6592 33254
rect 6552 32904 6604 32910
rect 6552 32846 6604 32852
rect 6564 31754 6592 32846
rect 6840 31958 6868 33390
rect 7012 32292 7064 32298
rect 7012 32234 7064 32240
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6564 31726 6776 31754
rect 6644 31476 6696 31482
rect 6644 31418 6696 31424
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6564 30802 6592 31282
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6552 30796 6604 30802
rect 6552 30738 6604 30744
rect 6472 30258 6500 30738
rect 6656 30682 6684 31418
rect 6748 31210 6776 31726
rect 6840 31346 6868 31894
rect 7024 31822 7052 32234
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6736 31204 6788 31210
rect 6736 31146 6788 31152
rect 6748 30938 6776 31146
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6564 30666 6684 30682
rect 6552 30660 6684 30666
rect 6604 30654 6684 30660
rect 6552 30602 6604 30608
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6840 29238 6868 31282
rect 6932 29238 6960 31758
rect 7012 31680 7064 31686
rect 7012 31622 7064 31628
rect 7024 30938 7052 31622
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 7012 30660 7064 30666
rect 7012 30602 7064 30608
rect 7024 29238 7052 30602
rect 7116 30190 7144 33526
rect 7392 33386 7420 33934
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7392 32910 7420 33322
rect 7852 32910 7880 33934
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7564 32904 7616 32910
rect 7564 32846 7616 32852
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7392 32434 7420 32846
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7380 31408 7432 31414
rect 7380 31350 7432 31356
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7208 31142 7236 31282
rect 7288 31204 7340 31210
rect 7288 31146 7340 31152
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7208 29646 7236 31078
rect 7300 30734 7328 31146
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 6828 29232 6880 29238
rect 6828 29174 6880 29180
rect 6920 29232 6972 29238
rect 6920 29174 6972 29180
rect 7012 29232 7064 29238
rect 7012 29174 7064 29180
rect 6840 28966 6868 29174
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6828 28960 6880 28966
rect 6828 28902 6880 28908
rect 6656 28558 6684 28902
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6552 28484 6604 28490
rect 6552 28426 6604 28432
rect 6564 28150 6592 28426
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 6564 27962 6592 28086
rect 6472 27934 6592 27962
rect 6368 26512 6420 26518
rect 6368 26454 6420 26460
rect 6472 23118 6500 27934
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6564 24206 6592 27814
rect 6656 26994 6684 28494
rect 6840 27878 6868 28902
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6932 26926 6960 29174
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7208 28150 7236 28494
rect 7196 28144 7248 28150
rect 7196 28086 7248 28092
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7116 27849 7144 27950
rect 7102 27840 7158 27849
rect 7102 27775 7158 27784
rect 7208 27606 7236 28086
rect 7196 27600 7248 27606
rect 7196 27542 7248 27548
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6828 25900 6880 25906
rect 6828 25842 6880 25848
rect 6656 25770 6684 25842
rect 6644 25764 6696 25770
rect 6644 25706 6696 25712
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6748 24682 6776 25230
rect 6736 24676 6788 24682
rect 6736 24618 6788 24624
rect 6840 24562 6868 25842
rect 6932 25498 6960 25978
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6932 24818 6960 25434
rect 7116 25158 7144 27406
rect 7300 26994 7328 30670
rect 7392 30326 7420 31350
rect 7380 30320 7432 30326
rect 7380 30262 7432 30268
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7392 28422 7420 29582
rect 7484 29170 7512 30194
rect 7576 29646 7604 32846
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 7760 30734 7788 31622
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7852 30870 7880 31078
rect 7840 30864 7892 30870
rect 7840 30806 7892 30812
rect 7748 30728 7800 30734
rect 7748 30670 7800 30676
rect 7840 30728 7892 30734
rect 7840 30670 7892 30676
rect 7748 30592 7800 30598
rect 7852 30580 7880 30670
rect 7800 30552 7880 30580
rect 7748 30534 7800 30540
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7944 30138 7972 34478
rect 8220 33998 8248 34478
rect 8300 34196 8352 34202
rect 8300 34138 8352 34144
rect 8208 33992 8260 33998
rect 8208 33934 8260 33940
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 8036 32026 8064 32166
rect 8024 32020 8076 32026
rect 8024 31962 8076 31968
rect 8036 31822 8064 31962
rect 8128 31822 8156 32778
rect 8312 31822 8340 34138
rect 8760 33856 8812 33862
rect 8760 33798 8812 33804
rect 8772 33522 8800 33798
rect 8760 33516 8812 33522
rect 8760 33458 8812 33464
rect 8392 33380 8444 33386
rect 8392 33322 8444 33328
rect 8404 32910 8432 33322
rect 8772 33114 8800 33458
rect 8760 33108 8812 33114
rect 8760 33050 8812 33056
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 9140 32502 9168 35022
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 8128 30870 8156 31758
rect 8208 31408 8260 31414
rect 8206 31376 8208 31385
rect 8260 31376 8262 31385
rect 8206 31311 8262 31320
rect 8116 30864 8168 30870
rect 8116 30806 8168 30812
rect 7668 29646 7696 30126
rect 7944 30110 8064 30138
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7484 28558 7512 29106
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7392 27130 7420 28358
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7380 27124 7432 27130
rect 7380 27066 7432 27072
rect 7484 26994 7512 27542
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7300 25906 7328 26930
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6748 24534 6868 24562
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6564 22030 6592 24142
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23254 6684 24006
rect 6748 23730 6776 24534
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 7024 23798 7052 24006
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6656 22098 6684 23054
rect 6748 22098 6776 23666
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6564 19854 6592 21830
rect 6656 21622 6684 22034
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6840 21554 6868 22102
rect 7024 21554 7052 22374
rect 7208 22234 7236 22578
rect 7484 22438 7512 22918
rect 7576 22642 7604 29446
rect 7668 24954 7696 29582
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7760 27946 7788 28970
rect 8036 28626 8064 30110
rect 8208 29572 8260 29578
rect 8208 29514 8260 29520
rect 8220 29102 8248 29514
rect 8208 29096 8260 29102
rect 8208 29038 8260 29044
rect 8024 28620 8076 28626
rect 8024 28562 8076 28568
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7760 27538 7788 27882
rect 7748 27532 7800 27538
rect 7748 27474 7800 27480
rect 7852 27470 7880 28358
rect 8312 27946 8340 31758
rect 8772 31385 8800 32370
rect 9232 31754 9260 36246
rect 9324 35766 9352 37266
rect 11716 37262 11744 39200
rect 15028 39148 15056 39200
rect 15028 39120 15240 39148
rect 15212 37262 15240 39120
rect 18340 37262 18368 39200
rect 21652 39166 21680 39200
rect 21640 39160 21692 39166
rect 21640 39102 21692 39108
rect 22100 39160 22152 39166
rect 22100 39102 22152 39108
rect 22112 37262 22140 39102
rect 24964 37262 24992 39200
rect 28276 37262 28304 39200
rect 31588 39114 31616 39200
rect 31588 39086 31800 39114
rect 31772 37262 31800 39086
rect 34900 37754 34928 39200
rect 34808 37726 34928 37754
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 9680 37188 9732 37194
rect 9680 37130 9732 37136
rect 12072 37188 12124 37194
rect 12072 37130 12124 37136
rect 16212 37188 16264 37194
rect 16212 37130 16264 37136
rect 18788 37188 18840 37194
rect 18788 37130 18840 37136
rect 9588 37120 9640 37126
rect 9588 37062 9640 37068
rect 9600 36922 9628 37062
rect 9588 36916 9640 36922
rect 9588 36858 9640 36864
rect 9600 36106 9628 36858
rect 9692 36242 9720 37130
rect 11060 36916 11112 36922
rect 11060 36858 11112 36864
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 10140 36100 10192 36106
rect 10140 36042 10192 36048
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9864 35692 9916 35698
rect 9864 35634 9916 35640
rect 9876 35562 9904 35634
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 9864 35556 9916 35562
rect 9864 35498 9916 35504
rect 9404 35488 9456 35494
rect 9404 35430 9456 35436
rect 9416 35086 9444 35430
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9876 34746 9904 35498
rect 9968 34950 9996 35566
rect 10152 35086 10180 36042
rect 10600 35216 10652 35222
rect 10600 35158 10652 35164
rect 10140 35080 10192 35086
rect 10140 35022 10192 35028
rect 9956 34944 10008 34950
rect 9956 34886 10008 34892
rect 9968 34746 9996 34886
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 10152 34542 10180 35022
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10612 34066 10640 35158
rect 10600 34060 10652 34066
rect 10600 34002 10652 34008
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9416 33590 9444 33934
rect 9864 33924 9916 33930
rect 9864 33866 9916 33872
rect 9404 33584 9456 33590
rect 9404 33526 9456 33532
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 9324 32298 9352 33390
rect 9312 32292 9364 32298
rect 9312 32234 9364 32240
rect 9324 31822 9352 32234
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9048 31726 9260 31754
rect 8758 31376 8814 31385
rect 8758 31311 8814 31320
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 8300 27940 8352 27946
rect 8300 27882 8352 27888
rect 7840 27464 7892 27470
rect 8300 27464 8352 27470
rect 7840 27406 7892 27412
rect 8128 27412 8300 27418
rect 8128 27406 8352 27412
rect 8128 27390 8340 27406
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7668 24070 7696 24890
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7760 22710 7788 27270
rect 8128 26994 8156 27390
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8220 26994 8248 27066
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8024 26852 8076 26858
rect 8024 26794 8076 26800
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 7852 24886 7880 25162
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 7852 24070 7880 24822
rect 8036 24274 8064 26794
rect 8220 26790 8248 26930
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8128 25906 8156 26522
rect 8404 26450 8432 30262
rect 9048 30258 9076 31726
rect 9324 31362 9352 31758
rect 9140 31334 9352 31362
rect 8760 30252 8812 30258
rect 8760 30194 8812 30200
rect 9036 30252 9088 30258
rect 9036 30194 9088 30200
rect 8772 29170 8800 30194
rect 9036 30048 9088 30054
rect 9036 29990 9088 29996
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 9048 29050 9076 29990
rect 8956 29022 9076 29050
rect 9140 29050 9168 31334
rect 9312 31204 9364 31210
rect 9312 31146 9364 31152
rect 9324 30870 9352 31146
rect 9312 30864 9364 30870
rect 9312 30806 9364 30812
rect 9416 30734 9444 33526
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9692 33046 9720 33458
rect 9680 33040 9732 33046
rect 9680 32982 9732 32988
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9508 31822 9536 32710
rect 9692 32502 9720 32982
rect 9876 32910 9904 33866
rect 10612 33522 10640 34002
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10048 33448 10100 33454
rect 10048 33390 10100 33396
rect 10060 32910 10088 33390
rect 10140 33040 10192 33046
rect 10140 32982 10192 32988
rect 9864 32904 9916 32910
rect 10048 32904 10100 32910
rect 9916 32864 9996 32892
rect 9864 32846 9916 32852
rect 9680 32496 9732 32502
rect 9680 32438 9732 32444
rect 9772 32428 9824 32434
rect 9772 32370 9824 32376
rect 9864 32428 9916 32434
rect 9864 32370 9916 32376
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9692 32026 9720 32302
rect 9784 32026 9812 32370
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9496 31816 9548 31822
rect 9496 31758 9548 31764
rect 9600 31686 9628 31894
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9600 30870 9628 31622
rect 9692 31482 9720 31962
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9588 30864 9640 30870
rect 9784 30818 9812 31758
rect 9588 30806 9640 30812
rect 9692 30802 9812 30818
rect 9680 30796 9812 30802
rect 9732 30790 9812 30796
rect 9680 30738 9732 30744
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9416 30326 9444 30670
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 9140 29022 9260 29050
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 8116 25900 8168 25906
rect 8116 25842 8168 25848
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 8128 24206 8156 25842
rect 8312 25770 8340 26318
rect 8300 25764 8352 25770
rect 8300 25706 8352 25712
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8220 25226 8248 25298
rect 8312 25226 8340 25706
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 8300 25220 8352 25226
rect 8300 25162 8352 25168
rect 8220 25106 8248 25162
rect 8220 25078 8340 25106
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7852 23798 7880 24006
rect 7840 23792 7892 23798
rect 7840 23734 7892 23740
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7196 22228 7248 22234
rect 7196 22170 7248 22176
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6748 19786 6776 21490
rect 6840 21146 6868 21490
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6840 19854 6868 20538
rect 6932 19854 6960 21490
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5644 17678 5672 18702
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 5644 16658 5672 17614
rect 6564 17610 6592 18566
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16250 6592 16458
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6656 16046 6684 19314
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6748 18834 6776 19110
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6840 18630 6868 19654
rect 6932 18834 6960 19790
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 16250 6960 16390
rect 7024 16250 7052 21490
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 20874 7144 21286
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 20058 7144 20402
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7576 19514 7604 22578
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7668 21622 7696 21966
rect 8128 21962 8156 24142
rect 8312 22778 8340 25078
rect 8404 23730 8432 26386
rect 8772 26382 8800 26862
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8496 24886 8524 25094
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7668 21146 7696 21558
rect 8128 21486 8156 21898
rect 8220 21554 8248 22578
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8312 22098 8340 22442
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8312 21622 8340 22034
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7944 19446 7972 19654
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 17882 7420 18770
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7944 16250 7972 19382
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8312 17678 8340 18226
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8312 16658 8340 17614
rect 8404 17270 8432 21286
rect 8496 19378 8524 24822
rect 8588 23526 8616 25842
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 18290 8616 18566
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8680 17202 8708 18702
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 7760 15502 7788 15846
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7852 15094 7880 15438
rect 8404 15434 8432 16458
rect 8680 16114 8708 17138
rect 8772 16794 8800 22646
rect 8956 21350 8984 29022
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9140 28558 9168 28902
rect 9232 28762 9260 29022
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9232 28082 9260 28698
rect 9324 28694 9352 30126
rect 9416 29646 9444 30262
rect 9692 30258 9720 30738
rect 9876 30326 9904 32370
rect 9864 30320 9916 30326
rect 9864 30262 9916 30268
rect 9680 30252 9732 30258
rect 9680 30194 9732 30200
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9968 29170 9996 32864
rect 10048 32846 10100 32852
rect 10060 29170 10088 32846
rect 10152 32434 10180 32982
rect 10612 32978 10640 33458
rect 10600 32972 10652 32978
rect 10600 32914 10652 32920
rect 10600 32768 10652 32774
rect 10600 32710 10652 32716
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 10612 32230 10640 32710
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10336 31890 10364 31962
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10140 31748 10192 31754
rect 10140 31690 10192 31696
rect 10152 29850 10180 31690
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10140 29844 10192 29850
rect 10140 29786 10192 29792
rect 10152 29578 10180 29786
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10244 29458 10272 31282
rect 10336 30326 10364 31826
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10520 31278 10548 31758
rect 10508 31272 10560 31278
rect 10508 31214 10560 31220
rect 10324 30320 10376 30326
rect 10324 30262 10376 30268
rect 10520 30122 10548 31214
rect 10508 30116 10560 30122
rect 10508 30058 10560 30064
rect 10152 29430 10272 29458
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9956 29164 10008 29170
rect 9956 29106 10008 29112
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9508 28694 9536 29106
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9312 28688 9364 28694
rect 9312 28630 9364 28636
rect 9496 28688 9548 28694
rect 9496 28630 9548 28636
rect 9220 28076 9272 28082
rect 9140 28036 9220 28064
rect 9140 27606 9168 28036
rect 9220 28018 9272 28024
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9128 27600 9180 27606
rect 9128 27542 9180 27548
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9048 26994 9076 27270
rect 9232 26994 9260 27814
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9508 26314 9536 28630
rect 9600 28422 9628 29038
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9692 28490 9720 28970
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 10060 28082 10088 29106
rect 10152 28966 10180 29430
rect 10520 29034 10548 30058
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28490 10180 28902
rect 10612 28694 10640 32166
rect 11072 30734 11100 36858
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11716 35834 11744 36042
rect 11888 36032 11940 36038
rect 11888 35974 11940 35980
rect 11900 35894 11928 35974
rect 11808 35866 11928 35894
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11808 35630 11836 35866
rect 12084 35698 12112 37130
rect 14188 36916 14240 36922
rect 14188 36858 14240 36864
rect 13176 36780 13228 36786
rect 13176 36722 13228 36728
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 12716 36576 12768 36582
rect 12716 36518 12768 36524
rect 12728 36174 12756 36518
rect 13188 36378 13216 36722
rect 13176 36372 13228 36378
rect 13176 36314 13228 36320
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12912 35766 12940 36178
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 12900 35760 12952 35766
rect 12900 35702 12952 35708
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11808 35018 11836 35566
rect 12084 35154 12112 35634
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 11796 35012 11848 35018
rect 11796 34954 11848 34960
rect 12084 34542 12112 35090
rect 13280 35086 13308 36110
rect 13268 35080 13320 35086
rect 13268 35022 13320 35028
rect 12624 35012 12676 35018
rect 12624 34954 12676 34960
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 11532 33522 11560 33934
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 11532 32910 11560 33458
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11532 32366 11560 32846
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11532 31906 11560 32302
rect 11900 32298 11928 33934
rect 12256 33516 12308 33522
rect 12176 33476 12256 33504
rect 12176 32434 12204 33476
rect 12256 33458 12308 33464
rect 12544 32910 12572 33934
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 12164 32428 12216 32434
rect 12164 32370 12216 32376
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 11532 31878 11744 31906
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10692 30320 10744 30326
rect 10692 30262 10744 30268
rect 10600 28688 10652 28694
rect 10600 28630 10652 28636
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10140 28484 10192 28490
rect 10140 28426 10192 28432
rect 10152 28082 10180 28426
rect 10520 28082 10548 28494
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9324 25498 9352 26182
rect 9508 25906 9536 26250
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9784 25838 9812 26182
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 9416 24274 9444 25774
rect 9680 25288 9732 25294
rect 9784 25242 9812 25774
rect 9732 25236 9812 25242
rect 9680 25230 9812 25236
rect 9692 25214 9812 25230
rect 9784 24886 9812 25214
rect 9772 24880 9824 24886
rect 9772 24822 9824 24828
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9692 24698 9720 24754
rect 9508 24670 9720 24698
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9508 24614 9536 24670
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24274 9628 24550
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23798 9168 24006
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 19854 8984 21286
rect 9140 20534 9168 21966
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9508 20874 9536 21490
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 9140 19922 9168 20470
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9140 18358 9168 19858
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9232 19514 9260 19722
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9692 19378 9720 24670
rect 9784 23526 9812 24686
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9324 18766 9352 19314
rect 9692 18766 9720 19314
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9324 18426 9352 18702
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9416 18154 9444 18634
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8864 16590 8892 16934
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8956 16250 8984 17070
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 15706 8524 15846
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7852 13938 7880 15030
rect 8404 15026 8432 15370
rect 9140 15094 9168 16594
rect 9508 16046 9536 16730
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 9508 14958 9536 15982
rect 9876 15162 9904 27270
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9968 25226 9996 25638
rect 10152 25362 10180 28018
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10244 26994 10272 27474
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10244 25906 10272 26726
rect 10336 26586 10364 27338
rect 10520 26994 10548 28018
rect 10612 28014 10640 28630
rect 10600 28008 10652 28014
rect 10600 27950 10652 27956
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10416 26784 10468 26790
rect 10416 26726 10468 26732
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10428 26518 10456 26726
rect 10416 26512 10468 26518
rect 10416 26454 10468 26460
rect 10612 26042 10640 27950
rect 10704 27606 10732 30262
rect 11072 28762 11100 30670
rect 11152 29844 11204 29850
rect 11152 29786 11204 29792
rect 11164 29306 11192 29786
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11164 28966 11192 29106
rect 11152 28960 11204 28966
rect 11152 28902 11204 28908
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 11532 28558 11560 31878
rect 11716 31822 11744 31878
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11612 31816 11664 31822
rect 11612 31758 11664 31764
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 11624 31482 11652 31758
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11612 31476 11664 31482
rect 11612 31418 11664 31424
rect 11624 30802 11652 31418
rect 11716 31226 11744 31622
rect 11808 31414 11836 31826
rect 11796 31408 11848 31414
rect 11796 31350 11848 31356
rect 11716 31198 11836 31226
rect 11808 31142 11836 31198
rect 11796 31136 11848 31142
rect 11796 31078 11848 31084
rect 11612 30796 11664 30802
rect 11664 30756 11744 30784
rect 11612 30738 11664 30744
rect 11612 30660 11664 30666
rect 11612 30602 11664 30608
rect 11624 30122 11652 30602
rect 11716 30240 11744 30756
rect 11808 30734 11836 31078
rect 11900 30938 11928 32234
rect 11980 31952 12032 31958
rect 11980 31894 12032 31900
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11992 30734 12020 31894
rect 12084 31890 12112 32370
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11796 30252 11848 30258
rect 11716 30212 11796 30240
rect 11796 30194 11848 30200
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 11888 30116 11940 30122
rect 11888 30058 11940 30064
rect 11900 29578 11928 30058
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11716 29238 11744 29446
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11808 28490 11836 29514
rect 11992 29306 12020 30534
rect 12084 29850 12112 31826
rect 12176 30938 12204 32370
rect 12452 32230 12480 32846
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 12438 31920 12494 31929
rect 12438 31855 12494 31864
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12360 31414 12388 31758
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12256 31340 12308 31346
rect 12256 31282 12308 31288
rect 12164 30932 12216 30938
rect 12164 30874 12216 30880
rect 12268 30734 12296 31282
rect 12256 30728 12308 30734
rect 12256 30670 12308 30676
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 11980 28960 12032 28966
rect 11980 28902 12032 28908
rect 11992 28762 12020 28902
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 11796 28484 11848 28490
rect 11796 28426 11848 28432
rect 10784 28416 10836 28422
rect 10784 28358 10836 28364
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 10796 28150 10824 28358
rect 11716 28218 11744 28358
rect 11808 28218 11836 28426
rect 11704 28212 11756 28218
rect 11704 28154 11756 28160
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 10784 28144 10836 28150
rect 10784 28086 10836 28092
rect 10692 27600 10744 27606
rect 10692 27542 10744 27548
rect 11900 27470 11928 28698
rect 12360 27470 12388 29514
rect 12452 29170 12480 31855
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10416 25900 10468 25906
rect 10692 25900 10744 25906
rect 10416 25842 10468 25848
rect 10612 25860 10692 25888
rect 10232 25696 10284 25702
rect 10232 25638 10284 25644
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 9956 25220 10008 25226
rect 9956 25162 10008 25168
rect 9968 23118 9996 25162
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9968 21690 9996 21898
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10152 21554 10180 22714
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 10244 15502 10272 25638
rect 10336 25430 10364 25638
rect 10324 25424 10376 25430
rect 10324 25366 10376 25372
rect 10336 24206 10364 25366
rect 10428 24886 10456 25842
rect 10612 25294 10640 25860
rect 10692 25842 10744 25848
rect 10796 25786 10824 27406
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25906 11008 26182
rect 11164 26042 11192 26250
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 12268 25974 12296 26522
rect 12256 25968 12308 25974
rect 12256 25910 12308 25916
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10704 25758 10824 25786
rect 11980 25764 12032 25770
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10428 24290 10456 24686
rect 10520 24410 10548 24754
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10428 24262 10548 24290
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10520 23118 10548 24262
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10336 22778 10364 22986
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10520 21554 10548 23054
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 20942 10364 21286
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19446 10548 19654
rect 10508 19440 10560 19446
rect 10508 19382 10560 19388
rect 10612 19378 10640 25230
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18290 10364 18634
rect 10612 18358 10640 19314
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10612 17882 10640 18158
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10520 16454 10548 17206
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10428 15706 10456 16050
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14006 9536 14758
rect 9876 14074 9904 14962
rect 10520 14482 10548 16390
rect 10704 16250 10732 25758
rect 11980 25706 12032 25712
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 24138 10916 24550
rect 10876 24132 10928 24138
rect 10876 24074 10928 24080
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10888 21486 10916 21830
rect 10980 21622 11008 21830
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11072 21554 11100 22714
rect 11992 22710 12020 25706
rect 12360 25294 12388 27406
rect 12452 27334 12480 29106
rect 12544 28558 12572 29990
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12636 28422 12664 34954
rect 13372 34610 13400 36722
rect 14200 36310 14228 36858
rect 15200 36848 15252 36854
rect 15200 36790 15252 36796
rect 15936 36848 15988 36854
rect 15936 36790 15988 36796
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 15108 36712 15160 36718
rect 15108 36654 15160 36660
rect 14188 36304 14240 36310
rect 14188 36246 14240 36252
rect 13452 36032 13504 36038
rect 13452 35974 13504 35980
rect 13464 35154 13492 35974
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 32026 12756 32166
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12820 31822 12848 32778
rect 12992 32292 13044 32298
rect 12992 32234 13044 32240
rect 13004 31958 13032 32234
rect 12992 31952 13044 31958
rect 12992 31894 13044 31900
rect 12808 31816 12860 31822
rect 12860 31776 12940 31804
rect 12808 31758 12860 31764
rect 12912 31754 12940 31776
rect 12912 31726 13032 31754
rect 13004 31346 13032 31726
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 13004 30734 13032 31282
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13004 30190 13032 30670
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 13004 29170 13032 30126
rect 13188 29209 13216 34478
rect 13372 31414 13400 34546
rect 13636 34536 13688 34542
rect 13636 34478 13688 34484
rect 13648 33658 13676 34478
rect 13728 33924 13780 33930
rect 13728 33866 13780 33872
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13544 33448 13596 33454
rect 13544 33390 13596 33396
rect 13556 32910 13584 33390
rect 13740 33114 13768 33866
rect 14188 33856 14240 33862
rect 14188 33798 14240 33804
rect 14096 33516 14148 33522
rect 14096 33458 14148 33464
rect 14108 33114 14136 33458
rect 14200 33318 14228 33798
rect 14568 33522 14596 36654
rect 15120 36174 15148 36654
rect 15212 36378 15240 36790
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15948 36242 15976 36790
rect 16028 36576 16080 36582
rect 16028 36518 16080 36524
rect 16040 36242 16068 36518
rect 15936 36236 15988 36242
rect 15936 36178 15988 36184
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 15108 36168 15160 36174
rect 15108 36110 15160 36116
rect 15120 35698 15148 36110
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 14740 35488 14792 35494
rect 14740 35430 14792 35436
rect 14752 34610 14780 35430
rect 15948 35154 15976 36178
rect 16120 36168 16172 36174
rect 16120 36110 16172 36116
rect 15936 35148 15988 35154
rect 15936 35090 15988 35096
rect 15844 35012 15896 35018
rect 15844 34954 15896 34960
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 15028 34134 15056 34478
rect 15016 34128 15068 34134
rect 15016 34070 15068 34076
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 14752 33658 14780 33934
rect 14740 33652 14792 33658
rect 14740 33594 14792 33600
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14464 33448 14516 33454
rect 14464 33390 14516 33396
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 13728 33108 13780 33114
rect 13728 33050 13780 33056
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14372 32768 14424 32774
rect 14372 32710 14424 32716
rect 13648 32502 13676 32710
rect 13728 32564 13780 32570
rect 13728 32506 13780 32512
rect 13636 32496 13688 32502
rect 13636 32438 13688 32444
rect 13740 32337 13768 32506
rect 14292 32502 14320 32710
rect 14384 32570 14412 32710
rect 14476 32570 14504 33390
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 14556 32836 14608 32842
rect 14608 32796 14688 32824
rect 14556 32778 14608 32784
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14280 32496 14332 32502
rect 14280 32438 14332 32444
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 13726 32328 13782 32337
rect 13726 32263 13782 32272
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13556 31482 13584 31622
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13360 31408 13412 31414
rect 13360 31350 13412 31356
rect 13634 31376 13690 31385
rect 13634 31311 13636 31320
rect 13688 31311 13690 31320
rect 13636 31282 13688 31288
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30802 13768 31214
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13832 30598 13860 32166
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 14200 30734 14228 31078
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 13820 30592 13872 30598
rect 13820 30534 13872 30540
rect 13820 29776 13872 29782
rect 13820 29718 13872 29724
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 13174 29200 13230 29209
rect 12992 29164 13044 29170
rect 13280 29170 13308 29650
rect 13832 29238 13860 29718
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14108 29510 14136 29582
rect 14188 29572 14240 29578
rect 14292 29560 14320 31282
rect 14384 30394 14412 32166
rect 14568 31890 14596 32370
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14660 30938 14688 32796
rect 14752 32026 14780 32846
rect 14844 32042 14872 32914
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14936 32230 14964 32370
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14844 32026 14964 32042
rect 14740 32020 14792 32026
rect 14740 31962 14792 31968
rect 14832 32020 14964 32026
rect 14884 32014 14964 32020
rect 14832 31962 14884 31968
rect 14832 31884 14884 31890
rect 14832 31826 14884 31832
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14648 30932 14700 30938
rect 14648 30874 14700 30880
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14568 30054 14596 30874
rect 14740 30592 14792 30598
rect 14740 30534 14792 30540
rect 14752 30190 14780 30534
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 14464 30048 14516 30054
rect 14464 29990 14516 29996
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14476 29578 14504 29990
rect 14240 29532 14320 29560
rect 14188 29514 14240 29520
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 14108 29170 14136 29446
rect 13174 29135 13230 29144
rect 13268 29164 13320 29170
rect 12992 29106 13044 29112
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 28082 12664 28358
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12820 27130 12848 27338
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 13004 26994 13032 29106
rect 13188 29050 13216 29135
rect 13268 29106 13320 29112
rect 13912 29164 13964 29170
rect 13912 29106 13964 29112
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 13188 29022 13308 29050
rect 13924 29034 13952 29106
rect 13176 28960 13228 28966
rect 13176 28902 13228 28908
rect 13188 27878 13216 28902
rect 13176 27872 13228 27878
rect 13176 27814 13228 27820
rect 13188 27062 13216 27814
rect 13176 27056 13228 27062
rect 13176 26998 13228 27004
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12452 25974 12480 26862
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12084 24070 12112 24346
rect 12360 24206 12388 25230
rect 12452 24818 12480 25910
rect 12544 25838 12572 26182
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12544 25226 12572 25774
rect 12532 25220 12584 25226
rect 12532 25162 12584 25168
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12728 24682 12756 25842
rect 13004 25498 13032 25842
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13188 25294 13216 25638
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 12716 24676 12768 24682
rect 12716 24618 12768 24624
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12360 23798 12388 24142
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12360 23118 12388 23734
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 12360 22642 12388 23054
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 11072 21010 11100 21490
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11072 20806 11100 20946
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11428 20936 11480 20942
rect 11480 20884 11560 20890
rect 11428 20878 11560 20884
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10980 19378 11008 19722
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10980 18426 11008 19314
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11164 17270 11192 20878
rect 11440 20862 11560 20878
rect 11532 20398 11560 20862
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11532 19378 11560 20334
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11256 17678 11284 18022
rect 11532 17678 11560 19314
rect 11716 18358 11744 19790
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 11072 16182 11100 16526
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11532 16114 11560 17614
rect 12084 17202 12112 20742
rect 13280 18970 13308 29022
rect 13912 29028 13964 29034
rect 13912 28970 13964 28976
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13464 28694 13492 28902
rect 13452 28688 13504 28694
rect 13452 28630 13504 28636
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13372 28150 13400 28426
rect 13360 28144 13412 28150
rect 13360 28086 13412 28092
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13372 26994 13400 27950
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13464 25294 13492 27270
rect 14016 27062 14044 27270
rect 14004 27056 14056 27062
rect 14004 26998 14056 27004
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13648 25906 13676 26250
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13648 25362 13676 25842
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13464 24886 13492 25230
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13648 24818 13676 25298
rect 14016 25158 14044 26998
rect 14108 26518 14136 29106
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 14108 26042 14136 26454
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 23798 13952 24686
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 14016 22166 14044 25094
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 20534 13860 20742
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12268 17814 12296 18294
rect 12360 18086 12388 18702
rect 13280 18630 13308 18906
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12728 17746 12756 18566
rect 13372 18290 13400 18770
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13464 18222 13492 18294
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12912 17746 12940 18022
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12268 16522 12296 17478
rect 13096 17270 13124 17478
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12360 16590 12388 17070
rect 13096 16998 13124 17206
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16726 13124 16934
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15570 11192 15846
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 7852 12918 7880 13874
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13394 10272 13670
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 7852 12306 7880 12854
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 7852 11898 7880 12242
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 8772 10674 8800 12242
rect 9416 11898 9444 12786
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 10152 10810 10180 13262
rect 10428 12782 10456 13874
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10520 13462 10548 13806
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10980 12442 11008 13670
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11354 10364 12174
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10796 11694 10824 11766
rect 11072 11762 11100 12582
rect 11716 12306 11744 15574
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11808 15366 11836 15438
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 14414 11836 15302
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 14006 11836 14350
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11900 13870 11928 15438
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11992 15094 12020 15370
rect 12176 15366 12204 16390
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 12360 14958 12388 16526
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15570 13032 16050
rect 13464 15706 13492 18158
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11164 11762 11192 12106
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11762 12020 12038
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 10784 11688 10836 11694
rect 11992 11642 12020 11698
rect 10836 11636 10916 11642
rect 10784 11630 10916 11636
rect 10796 11614 10916 11630
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10796 11150 10824 11494
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 10336 10266 10364 10542
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10428 9654 10456 11086
rect 10888 10266 10916 11614
rect 11900 11614 12020 11642
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11218 11744 11494
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11900 11150 11928 11614
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11150 12020 11494
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10520 9586 10548 9998
rect 10888 9722 10916 10202
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 10796 9178 10824 9522
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 11072 7954 11100 10066
rect 11348 10062 11376 10950
rect 12084 10130 12112 14894
rect 12912 14618 12940 14894
rect 13280 14618 13308 14962
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12268 12986 12296 14282
rect 12912 13870 12940 14282
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 12986 12940 13806
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11354 12204 12174
rect 12268 11898 12296 12922
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12306 12756 12786
rect 13188 12782 13216 14010
rect 13372 13870 13400 14486
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13832 13802 13860 17546
rect 14200 14414 14228 22510
rect 14292 21078 14320 29532
rect 14464 29572 14516 29578
rect 14464 29514 14516 29520
rect 14568 28994 14596 29990
rect 14844 29306 14872 31826
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14568 28966 14688 28994
rect 14660 28218 14688 28966
rect 14752 28558 14780 29038
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14936 28422 14964 32014
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14924 28416 14976 28422
rect 14924 28358 14976 28364
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14844 27946 14872 28358
rect 14832 27940 14884 27946
rect 14832 27882 14884 27888
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14372 26852 14424 26858
rect 14372 26794 14424 26800
rect 14384 26450 14412 26794
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14476 24750 14504 26862
rect 14844 26586 14872 26930
rect 15028 26874 15056 34070
rect 15292 34060 15344 34066
rect 15292 34002 15344 34008
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15212 32994 15240 33458
rect 15304 33114 15332 34002
rect 15476 33856 15528 33862
rect 15476 33798 15528 33804
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 15212 32966 15332 32994
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15120 31906 15148 32302
rect 15212 32026 15240 32846
rect 15304 32722 15332 32966
rect 15396 32960 15424 33458
rect 15488 33318 15516 33798
rect 15660 33448 15712 33454
rect 15660 33390 15712 33396
rect 15568 33380 15620 33386
rect 15568 33322 15620 33328
rect 15476 33312 15528 33318
rect 15476 33254 15528 33260
rect 15476 32972 15528 32978
rect 15396 32932 15476 32960
rect 15476 32914 15528 32920
rect 15580 32910 15608 33322
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15304 32694 15608 32722
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15292 32224 15344 32230
rect 15292 32166 15344 32172
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15120 31878 15240 31906
rect 15212 31686 15240 31878
rect 15200 31680 15252 31686
rect 15200 31622 15252 31628
rect 15304 31142 15332 32166
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15120 30161 15148 30670
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15106 30152 15162 30161
rect 15106 30087 15162 30096
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15120 28558 15148 28970
rect 15212 28558 15240 30534
rect 15396 30258 15424 32370
rect 15580 31958 15608 32694
rect 15568 31952 15620 31958
rect 15568 31894 15620 31900
rect 15476 30796 15528 30802
rect 15476 30738 15528 30744
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15292 30116 15344 30122
rect 15292 30058 15344 30064
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 14936 26846 15056 26874
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14476 21690 14504 22578
rect 14568 22522 14596 23054
rect 14660 22642 14688 23190
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14844 22710 14872 22986
rect 14832 22704 14884 22710
rect 14832 22646 14884 22652
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14568 22494 14780 22522
rect 14556 22160 14608 22166
rect 14556 22102 14608 22108
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14292 15502 14320 21014
rect 14476 20874 14504 21490
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14476 20602 14504 20810
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14568 19854 14596 22102
rect 14752 22098 14780 22494
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 21554 14688 21830
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14646 20904 14702 20913
rect 14646 20839 14648 20848
rect 14700 20839 14702 20848
rect 14648 20810 14700 20816
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20602 14780 20742
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19258 14780 19654
rect 14844 19378 14872 19722
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14752 19242 14872 19258
rect 14752 19236 14884 19242
rect 14752 19230 14832 19236
rect 14832 19178 14884 19184
rect 14844 18834 14872 19178
rect 14936 19174 14964 26846
rect 15120 26382 15148 27066
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15198 26208 15254 26217
rect 15198 26143 15254 26152
rect 15212 25906 15240 26143
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15304 24138 15332 30058
rect 15396 28762 15424 30194
rect 15488 29714 15516 30738
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15580 30394 15608 30670
rect 15568 30388 15620 30394
rect 15568 30330 15620 30336
rect 15672 30122 15700 33390
rect 15856 33114 15884 34954
rect 16132 33658 16160 36110
rect 16224 35562 16252 37130
rect 17040 37120 17092 37126
rect 17040 37062 17092 37068
rect 17052 36786 17080 37062
rect 17040 36780 17092 36786
rect 17040 36722 17092 36728
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 16960 36106 16988 36518
rect 16948 36100 17000 36106
rect 16948 36042 17000 36048
rect 17052 35698 17080 36722
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 16212 35556 16264 35562
rect 16212 35498 16264 35504
rect 16224 35154 16252 35498
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16212 35148 16264 35154
rect 16212 35090 16264 35096
rect 16960 35086 16988 35430
rect 16948 35080 17000 35086
rect 16948 35022 17000 35028
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 17052 33998 17080 34342
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 16120 33652 16172 33658
rect 16120 33594 16172 33600
rect 16224 33590 16252 33934
rect 17776 33924 17828 33930
rect 17776 33866 17828 33872
rect 17868 33924 17920 33930
rect 17868 33866 17920 33872
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 16212 33584 16264 33590
rect 16212 33526 16264 33532
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 16302 32464 16358 32473
rect 16302 32399 16304 32408
rect 16356 32399 16358 32408
rect 16304 32370 16356 32376
rect 16028 32292 16080 32298
rect 16028 32234 16080 32240
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15844 32020 15896 32026
rect 15844 31962 15896 31968
rect 15856 31929 15884 31962
rect 15842 31920 15898 31929
rect 15948 31890 15976 32166
rect 15842 31855 15898 31864
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 16040 31822 16068 32234
rect 16120 32224 16172 32230
rect 16120 32166 16172 32172
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 16132 31686 16160 32166
rect 15752 31680 15804 31686
rect 15752 31622 15804 31628
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 15764 31414 15792 31622
rect 15752 31408 15804 31414
rect 15752 31350 15804 31356
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15764 30326 15792 30806
rect 15856 30734 15884 31282
rect 16672 31204 16724 31210
rect 16672 31146 16724 31152
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 15752 30320 15804 30326
rect 15752 30262 15804 30268
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 16224 29782 16252 31078
rect 16684 30734 16712 31146
rect 16304 30728 16356 30734
rect 16304 30670 16356 30676
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16316 30598 16344 30670
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 15844 29096 15896 29102
rect 15844 29038 15896 29044
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15212 22642 15240 23054
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15304 22094 15332 22918
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15028 22066 15332 22094
rect 15028 22030 15056 22066
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15396 21690 15424 22374
rect 15488 22234 15516 22578
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15580 22166 15608 22578
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15580 21962 15608 22102
rect 15672 22030 15700 22578
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15764 21894 15792 25230
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15212 19514 15240 21082
rect 15672 20942 15700 21286
rect 15856 21026 15884 29038
rect 16132 25294 16160 29514
rect 16224 29306 16252 29718
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16316 28558 16344 30534
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16500 29646 16528 30262
rect 16684 30258 16712 30670
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16776 29646 16804 33594
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 16960 32230 16988 33458
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 17144 31822 17172 32302
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 16868 31414 16896 31758
rect 16856 31408 16908 31414
rect 16856 31350 16908 31356
rect 17040 30660 17092 30666
rect 17040 30602 17092 30608
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 16500 28762 16528 29582
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16592 29238 16620 29446
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16776 28694 16804 29582
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16764 28688 16816 28694
rect 16764 28630 16816 28636
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16120 25288 16172 25294
rect 16172 25248 16252 25276
rect 16120 25230 16172 25236
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 22438 15976 23054
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15948 21418 15976 22374
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16040 21486 16068 21966
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 15856 20998 15976 21026
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15290 20496 15346 20505
rect 15290 20431 15292 20440
rect 15344 20431 15346 20440
rect 15292 20402 15344 20408
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14844 18290 14872 18770
rect 15212 18766 15240 19110
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14832 18284 14884 18290
rect 14752 18244 14832 18272
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17678 14688 18022
rect 14752 17678 14780 18244
rect 14832 18226 14884 18232
rect 14844 18154 14872 18226
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14568 15162 14596 15982
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 13938 14044 14282
rect 14200 14006 14228 14350
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 14016 13190 14044 13874
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12360 11830 12388 12106
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12360 11286 12388 11766
rect 12728 11694 12756 12242
rect 12912 12170 12940 12718
rect 13188 12170 13216 12718
rect 13280 12238 13308 12854
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12912 11626 12940 12106
rect 13280 11830 13308 12174
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 13556 10470 13584 12310
rect 13648 10674 13676 12786
rect 14200 12102 14228 13942
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13326 14596 13874
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11256 9586 11284 9930
rect 11348 9654 11376 9998
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11532 9586 11560 9862
rect 11808 9586 11836 9998
rect 13464 9722 13492 10406
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 11072 4690 11100 7890
rect 11164 7886 11192 9318
rect 11256 8634 11284 9522
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11808 8498 11836 9522
rect 13556 9450 13584 10406
rect 14016 9654 14044 11698
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 8498 12848 9318
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11808 7546 11836 8434
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 12820 7478 12848 8434
rect 13096 7886 13124 8502
rect 14108 8498 14136 11018
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10198 14228 10610
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14200 9654 14228 10134
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8974 14596 9318
rect 14752 8974 14780 10678
rect 14844 10062 14872 17614
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15028 17202 15056 17478
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15304 16522 15332 20402
rect 15580 20398 15608 20538
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15396 20058 15424 20334
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15580 19802 15608 20334
rect 15396 19774 15608 19802
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15396 19174 15424 19774
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19514 15608 19654
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 19440 15528 19446
rect 15672 19394 15700 19790
rect 15476 19382 15528 19388
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15488 18766 15516 19382
rect 15580 19366 15700 19394
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15304 14414 15332 15030
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15120 13938 15148 14282
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 13938 15240 14214
rect 15488 14006 15516 14282
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13530 15056 13806
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15304 13394 15332 13874
rect 15580 13734 15608 19366
rect 15856 19174 15884 20878
rect 15948 20330 15976 20998
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 15948 19786 15976 20266
rect 16040 19922 16068 20742
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18426 15884 19110
rect 15948 18970 15976 19314
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 16040 18154 16068 19246
rect 16224 18358 16252 25248
rect 16316 23594 16344 28494
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16500 26790 16528 28018
rect 16592 28014 16620 28494
rect 16580 28008 16632 28014
rect 16580 27950 16632 27956
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16408 26586 16436 26726
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16486 26208 16542 26217
rect 16486 26143 16542 26152
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16316 21622 16344 23530
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16408 21554 16436 21830
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16316 20398 16344 21422
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16408 19922 16436 21490
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 17338 15792 17478
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15936 17196 15988 17202
rect 15856 17156 15936 17184
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 16794 15700 17002
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15856 16658 15884 17156
rect 15936 17138 15988 17144
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 16114 15884 16594
rect 16040 16182 16068 18090
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16590 16160 17478
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 16224 14958 16252 16730
rect 16408 15026 16436 19654
rect 16500 18698 16528 26143
rect 16592 25294 16620 27270
rect 16776 26926 16804 28630
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16868 28082 16896 28494
rect 16960 28218 16988 29106
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 17052 27606 17080 30602
rect 17236 29850 17264 32914
rect 17604 32910 17632 33798
rect 17788 33522 17816 33866
rect 17880 33658 17908 33866
rect 17972 33658 18000 35022
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17960 33652 18012 33658
rect 17960 33594 18012 33600
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17604 32570 17632 32846
rect 17592 32564 17644 32570
rect 17592 32506 17644 32512
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17328 31278 17356 32370
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 17316 31272 17368 31278
rect 17316 31214 17368 31220
rect 17328 30433 17356 31214
rect 17314 30424 17370 30433
rect 17314 30359 17370 30368
rect 17420 30122 17448 32166
rect 17592 31884 17644 31890
rect 17592 31826 17644 31832
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17408 30116 17460 30122
rect 17408 30058 17460 30064
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 17420 27520 17448 29582
rect 17512 29102 17540 31214
rect 17604 30054 17632 31826
rect 17788 31278 17816 33458
rect 17972 33454 18000 33594
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 18064 33114 18092 36654
rect 18696 36100 18748 36106
rect 18696 36042 18748 36048
rect 18420 35828 18472 35834
rect 18420 35770 18472 35776
rect 18432 35698 18460 35770
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 18604 35692 18656 35698
rect 18604 35634 18656 35640
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18248 33114 18276 35430
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18340 33318 18368 35022
rect 18432 34950 18460 35634
rect 18616 35086 18644 35634
rect 18708 35630 18736 36042
rect 18696 35624 18748 35630
rect 18696 35566 18748 35572
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18708 35018 18736 35566
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 18432 33454 18460 34886
rect 18604 33992 18656 33998
rect 18604 33934 18656 33940
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18328 33312 18380 33318
rect 18328 33254 18380 33260
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 17776 31136 17828 31142
rect 17776 31078 17828 31084
rect 17684 30728 17736 30734
rect 17788 30716 17816 31078
rect 17736 30688 17816 30716
rect 17684 30670 17736 30676
rect 17788 30258 17816 30688
rect 17868 30728 17920 30734
rect 17920 30676 18000 30682
rect 17868 30670 18000 30676
rect 17880 30654 18000 30670
rect 18064 30666 18092 31962
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 17880 30258 17908 30534
rect 17776 30252 17828 30258
rect 17776 30194 17828 30200
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17774 30152 17830 30161
rect 17972 30138 18000 30654
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18156 30598 18184 31282
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 17774 30087 17776 30096
rect 17828 30087 17830 30096
rect 17880 30110 18000 30138
rect 17776 30058 17828 30064
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17604 29170 17632 29718
rect 17880 29646 17908 30110
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17684 29572 17736 29578
rect 17684 29514 17736 29520
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17500 29096 17552 29102
rect 17500 29038 17552 29044
rect 17696 28762 17724 29514
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 17972 28626 18000 29106
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17420 27492 17540 27520
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16960 25974 16988 26998
rect 17052 26858 17080 27270
rect 17144 27130 17172 27406
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 17420 26994 17448 27338
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17040 26852 17092 26858
rect 17040 26794 17092 26800
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17052 26382 17080 26794
rect 17236 26466 17264 26794
rect 17236 26450 17448 26466
rect 17224 26444 17448 26450
rect 17276 26438 17448 26444
rect 17224 26386 17276 26392
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 16948 25968 17000 25974
rect 16948 25910 17000 25916
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16592 23186 16620 24686
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 21010 16620 21354
rect 16684 21146 16712 22510
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16684 20534 16712 21082
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16684 20058 16712 20470
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16776 18714 16804 25162
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16868 24410 16896 24754
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16868 23730 16896 24210
rect 17236 23730 17264 26250
rect 17316 25832 17368 25838
rect 17316 25774 17368 25780
rect 17328 24206 17356 25774
rect 17420 24206 17448 26438
rect 17512 25770 17540 27492
rect 17696 26382 17724 27542
rect 17684 26376 17736 26382
rect 17736 26336 17816 26364
rect 17684 26318 17736 26324
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17500 25764 17552 25770
rect 17500 25706 17552 25712
rect 17696 25498 17724 25842
rect 17788 25838 17816 26336
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17776 25696 17828 25702
rect 17776 25638 17828 25644
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17696 24818 17724 25434
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17788 24206 17816 25638
rect 17880 24721 17908 28494
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 17972 26450 18000 27474
rect 18156 26926 18184 30262
rect 18248 28558 18276 33050
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18340 32570 18368 32846
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18328 32564 18380 32570
rect 18328 32506 18380 32512
rect 18340 30394 18368 32506
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 27606 18276 28494
rect 18340 28082 18368 30194
rect 18432 29306 18460 32710
rect 18524 31346 18552 33798
rect 18616 32978 18644 33934
rect 18708 33522 18736 34954
rect 18800 33969 18828 37130
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19444 36854 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19984 36712 20036 36718
rect 19984 36654 20036 36660
rect 18972 36304 19024 36310
rect 18972 36246 19024 36252
rect 18984 36106 19012 36246
rect 18972 36100 19024 36106
rect 18972 36042 19024 36048
rect 18984 35698 19012 36042
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 18972 35692 19024 35698
rect 18972 35634 19024 35640
rect 18786 33960 18842 33969
rect 18786 33895 18842 33904
rect 18984 33658 19012 35634
rect 19444 35086 19472 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34610 20024 36654
rect 20180 36582 20208 37198
rect 20996 37188 21048 37194
rect 20996 37130 21048 37136
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 22928 37188 22980 37194
rect 22928 37130 22980 37136
rect 21008 36786 21036 37130
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21548 36780 21600 36786
rect 21548 36722 21600 36728
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 20260 36168 20312 36174
rect 20260 36110 20312 36116
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20272 35154 20300 36110
rect 20364 35698 20392 36110
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20456 35170 20484 35974
rect 20548 35698 20576 36518
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20640 35170 20668 36722
rect 21272 36304 21324 36310
rect 21272 36246 21324 36252
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20732 35834 20760 36110
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 21284 35766 21312 36246
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21272 35760 21324 35766
rect 21272 35702 21324 35708
rect 20812 35624 20864 35630
rect 20812 35566 20864 35572
rect 20260 35148 20312 35154
rect 20456 35142 20576 35170
rect 20640 35142 20760 35170
rect 20260 35090 20312 35096
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19984 34128 20036 34134
rect 19984 34070 20036 34076
rect 19248 33924 19300 33930
rect 19248 33866 19300 33872
rect 18972 33652 19024 33658
rect 18972 33594 19024 33600
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 18892 31958 18920 33458
rect 18880 31952 18932 31958
rect 18880 31894 18932 31900
rect 18696 31680 18748 31686
rect 18696 31622 18748 31628
rect 18708 31346 18736 31622
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18604 30660 18656 30666
rect 18604 30602 18656 30608
rect 18616 30190 18644 30602
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18524 29714 18552 29990
rect 18512 29708 18564 29714
rect 18512 29650 18564 29656
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18512 29096 18564 29102
rect 18512 29038 18564 29044
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18236 27600 18288 27606
rect 18236 27542 18288 27548
rect 18248 26994 18276 27542
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 18156 26246 18184 26862
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18064 26042 18092 26182
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 18064 25362 18092 25978
rect 18156 25906 18184 26182
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 18064 24818 18092 25298
rect 18156 25294 18184 25706
rect 18248 25378 18276 26930
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18340 26382 18368 26794
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18248 25362 18368 25378
rect 18248 25356 18380 25362
rect 18248 25350 18328 25356
rect 18328 25298 18380 25304
rect 18524 25294 18552 29038
rect 18604 27532 18656 27538
rect 18708 27520 18736 31282
rect 18892 29034 18920 31894
rect 18984 31793 19012 33594
rect 18970 31784 19026 31793
rect 19260 31754 19288 33866
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19352 33046 19380 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19444 33522 19472 33594
rect 19996 33522 20024 34070
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 19628 33386 19656 33458
rect 19720 33425 19748 33458
rect 19892 33448 19944 33454
rect 19706 33416 19762 33425
rect 19616 33380 19668 33386
rect 19892 33390 19944 33396
rect 19706 33351 19762 33360
rect 19616 33322 19668 33328
rect 19628 33289 19656 33322
rect 19614 33280 19670 33289
rect 19614 33215 19670 33224
rect 19340 33040 19392 33046
rect 19340 32982 19392 32988
rect 19904 32774 19932 33390
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19340 32768 19392 32774
rect 19432 32768 19484 32774
rect 19340 32710 19392 32716
rect 19430 32736 19432 32745
rect 19892 32768 19944 32774
rect 19484 32736 19486 32745
rect 19352 31822 19380 32710
rect 19892 32710 19944 32716
rect 19430 32671 19486 32680
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19798 32056 19854 32065
rect 19798 31991 19854 32000
rect 19812 31958 19840 31991
rect 19800 31952 19852 31958
rect 19800 31894 19852 31900
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 18970 31719 19026 31728
rect 19168 31726 19288 31754
rect 18984 29170 19012 31719
rect 19168 31346 19196 31726
rect 19156 31340 19208 31346
rect 19156 31282 19208 31288
rect 19352 30802 19380 31758
rect 19444 31482 19472 31758
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19522 31376 19578 31385
rect 19522 31311 19578 31320
rect 19536 30938 19564 31311
rect 19524 30932 19576 30938
rect 19524 30874 19576 30880
rect 19340 30796 19392 30802
rect 19340 30738 19392 30744
rect 19628 30734 19656 31418
rect 19996 30938 20024 33254
rect 19984 30932 20036 30938
rect 19984 30874 20036 30880
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 29714 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 29850 20024 30874
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19340 29300 19392 29306
rect 19168 29260 19340 29288
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 19168 29102 19196 29260
rect 19340 29242 19392 29248
rect 19616 29164 19668 29170
rect 19616 29106 19668 29112
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 19248 29096 19300 29102
rect 19248 29038 19300 29044
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 19260 28490 19288 29038
rect 19628 29034 19656 29106
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19616 29028 19668 29034
rect 19616 28970 19668 28976
rect 19812 28762 19840 29038
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28082 20024 28426
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19996 27946 20024 28018
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19352 27674 19380 27882
rect 20088 27878 20116 34682
rect 20272 34474 20300 35090
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 34542 20392 34886
rect 20456 34678 20484 35022
rect 20548 35018 20576 35142
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20536 35012 20588 35018
rect 20536 34954 20588 34960
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20548 34626 20576 34954
rect 20640 34746 20668 35022
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 20168 34468 20220 34474
rect 20168 34410 20220 34416
rect 20260 34468 20312 34474
rect 20260 34410 20312 34416
rect 20180 33522 20208 34410
rect 20260 34128 20312 34134
rect 20260 34070 20312 34076
rect 20272 33998 20300 34070
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20272 33538 20300 33934
rect 20364 33658 20392 34478
rect 20456 34202 20484 34614
rect 20548 34610 20668 34626
rect 20548 34604 20680 34610
rect 20548 34598 20628 34604
rect 20628 34546 20680 34552
rect 20536 34536 20588 34542
rect 20536 34478 20588 34484
rect 20444 34196 20496 34202
rect 20444 34138 20496 34144
rect 20548 34134 20576 34478
rect 20536 34128 20588 34134
rect 20536 34070 20588 34076
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 20352 33652 20404 33658
rect 20352 33594 20404 33600
rect 20168 33516 20220 33522
rect 20272 33510 20392 33538
rect 20168 33458 20220 33464
rect 20364 33046 20392 33510
rect 20352 33040 20404 33046
rect 20258 33008 20314 33017
rect 20352 32982 20404 32988
rect 20180 32952 20258 32960
rect 20180 32932 20260 32952
rect 20180 31346 20208 32932
rect 20312 32943 20314 32952
rect 20260 32914 20312 32920
rect 20352 32904 20404 32910
rect 20352 32846 20404 32852
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20272 32502 20300 32710
rect 20260 32496 20312 32502
rect 20260 32438 20312 32444
rect 20364 31958 20392 32846
rect 20456 32434 20484 33934
rect 20536 33584 20588 33590
rect 20536 33526 20588 33532
rect 20548 33017 20576 33526
rect 20534 33008 20590 33017
rect 20534 32943 20590 32952
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20444 32224 20496 32230
rect 20548 32212 20576 32846
rect 20496 32184 20576 32212
rect 20444 32166 20496 32172
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20272 31414 20300 31622
rect 20260 31408 20312 31414
rect 20260 31350 20312 31356
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 20272 30258 20300 31214
rect 20352 31204 20404 31210
rect 20352 31146 20404 31152
rect 20364 30394 20392 31146
rect 20456 30938 20484 32166
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20352 30388 20404 30394
rect 20352 30330 20404 30336
rect 20364 30258 20392 30330
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20168 29232 20220 29238
rect 20168 29174 20220 29180
rect 20180 28218 20208 29174
rect 20272 29102 20300 29582
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 28212 20220 28218
rect 20168 28154 20220 28160
rect 20180 28082 20208 28154
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20260 28008 20312 28014
rect 20260 27950 20312 27956
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 18656 27492 18736 27520
rect 18604 27474 18656 27480
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 19352 27418 19380 27610
rect 20088 27470 20116 27814
rect 20076 27464 20128 27470
rect 19076 27062 19104 27406
rect 19352 27390 19472 27418
rect 20076 27406 20128 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19064 27056 19116 27062
rect 19064 26998 19116 27004
rect 19352 25974 19380 27270
rect 19444 26738 19472 27390
rect 19892 27328 19944 27334
rect 19944 27288 20024 27316
rect 19892 27270 19944 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19614 27024 19670 27033
rect 19614 26959 19670 26968
rect 19800 26988 19852 26994
rect 19444 26710 19564 26738
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19444 26353 19472 26522
rect 19430 26344 19486 26353
rect 19430 26279 19486 26288
rect 19536 26228 19564 26710
rect 19628 26382 19656 26959
rect 19800 26930 19852 26936
rect 19812 26382 19840 26930
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19720 26246 19748 26318
rect 19444 26200 19564 26228
rect 19708 26240 19760 26246
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 17866 24712 17922 24721
rect 17866 24647 17922 24656
rect 18420 24608 18472 24614
rect 18418 24576 18420 24585
rect 18472 24576 18474 24585
rect 18418 24511 18474 24520
rect 18708 24342 18736 25230
rect 19076 24818 19104 25298
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18696 24336 18748 24342
rect 18748 24296 18828 24324
rect 18696 24278 18748 24284
rect 18800 24206 18828 24296
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 17972 23866 18000 24142
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18248 23798 18276 24142
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16868 22506 16896 23666
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16592 18686 16804 18714
rect 16592 15178 16620 18686
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18290 16804 18566
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16776 15314 16804 18226
rect 16868 16114 16896 22034
rect 16960 21486 16988 23462
rect 17144 22098 17172 23598
rect 17236 22642 17264 23666
rect 17224 22636 17276 22642
rect 17276 22596 17356 22624
rect 17224 22578 17276 22584
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16960 19174 16988 20198
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 17678 16988 19110
rect 17052 17678 17080 20810
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17144 18970 17172 19722
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17144 17882 17172 18158
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17236 17814 17264 19858
rect 17328 19718 17356 22596
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17604 20913 17632 21558
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17590 20904 17646 20913
rect 17590 20839 17646 20848
rect 17604 20806 17632 20839
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17604 20058 17632 20402
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17420 19718 17448 19926
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17328 19378 17356 19654
rect 17420 19378 17448 19654
rect 17512 19514 17540 19790
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17512 17678 17540 19450
rect 17696 19378 17724 19858
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17144 16726 17172 17546
rect 17236 16998 17264 17614
rect 17604 17066 17632 18158
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 17134 17908 17614
rect 18064 17610 18092 21490
rect 18248 19446 18276 23734
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18524 22642 18552 22918
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18892 21690 18920 22578
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18340 20097 18368 20334
rect 18326 20088 18382 20097
rect 18326 20023 18382 20032
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18236 19440 18288 19446
rect 18234 19408 18236 19417
rect 18288 19408 18290 19417
rect 18234 19343 18290 19352
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17202 18276 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 16868 15434 16896 16050
rect 17512 15434 17540 16050
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 16776 15286 16896 15314
rect 16592 15150 16804 15178
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 11898 15240 12786
rect 15304 12714 15332 13330
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 15212 9926 15240 11834
rect 15488 11762 15516 12854
rect 15580 12306 15608 12854
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15672 12102 15700 13126
rect 15764 12238 15792 13330
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15304 10062 15332 10610
rect 15672 10606 15700 11698
rect 15764 11626 15792 12174
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9654 15240 9862
rect 15304 9722 15332 9998
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14384 8498 14412 8842
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14096 8492 14148 8498
rect 14372 8492 14424 8498
rect 14148 8452 14228 8480
rect 14096 8434 14148 8440
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12912 7002 12940 7822
rect 13096 7342 13124 7822
rect 13740 7410 13768 8298
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14108 7410 14136 7958
rect 14200 7886 14228 8452
rect 14372 8434 14424 8440
rect 14384 7886 14412 8434
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13740 6934 13768 7346
rect 13728 6928 13780 6934
rect 14108 6914 14136 7346
rect 14660 7342 14688 8570
rect 15488 8090 15516 9522
rect 15672 9110 15700 10542
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15488 7886 15516 8026
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15672 7410 15700 8230
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 13728 6870 13780 6876
rect 14016 6886 14136 6914
rect 14016 6798 14044 6886
rect 14660 6866 14688 7278
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14752 6798 14780 7346
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 14752 6186 14780 6734
rect 15488 6322 15516 6734
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15580 6254 15608 7142
rect 15672 6866 15700 7346
rect 15856 6914 15884 13738
rect 16120 13320 16172 13326
rect 16118 13288 16120 13297
rect 16172 13288 16174 13297
rect 16118 13223 16174 13232
rect 16132 12918 16160 13223
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11694 15976 12174
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 11830 16160 12106
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 11150 16068 11630
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9586 16068 9998
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16224 9178 16252 14758
rect 16500 11898 16528 15030
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 12850 16620 13330
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 11286 16528 11834
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16592 11150 16620 12786
rect 16776 12374 16804 15150
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16684 12102 16712 12242
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 16040 8498 16068 8842
rect 16316 8498 16344 11018
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 8974 16528 9318
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16040 8090 16068 8434
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16500 7410 16528 8298
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 15856 6886 15976 6914
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15948 6798 15976 6886
rect 16500 6798 16528 7346
rect 16868 6914 16896 15286
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 8498 16988 14758
rect 17236 14618 17264 14962
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 9042 17080 13874
rect 17236 13870 17264 14214
rect 17328 14074 17356 14962
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17512 13938 17540 14826
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17236 12782 17264 13806
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11830 17172 12242
rect 17236 12238 17264 12582
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17236 11150 17264 12174
rect 17328 11762 17356 12786
rect 17420 12170 17448 13806
rect 17604 13326 17632 14350
rect 17500 13320 17552 13326
rect 17498 13288 17500 13297
rect 17592 13320 17644 13326
rect 17552 13288 17554 13297
rect 17592 13262 17644 13268
rect 17498 13223 17554 13232
rect 17696 12850 17724 15846
rect 17880 15502 17908 15982
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17788 14278 17816 14962
rect 18064 14890 18092 15098
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14482 17908 14758
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13938 17816 14214
rect 18156 14006 18184 14826
rect 18248 14618 18276 14894
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18248 14006 18276 14554
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12306 17540 12718
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17696 12102 17724 12650
rect 17880 12646 17908 13262
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17868 12436 17920 12442
rect 18340 12434 18368 18702
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17746 18644 18022
rect 18708 17746 18736 19654
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19076 19174 19104 19246
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18902 19104 19110
rect 19168 18902 19196 21490
rect 19260 20534 19288 24890
rect 19352 24886 19380 25910
rect 19444 25242 19472 26200
rect 19708 26182 19760 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 19904 25430 19932 25978
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19996 25294 20024 27288
rect 20272 27130 20300 27950
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20166 26344 20222 26353
rect 20166 26279 20222 26288
rect 20076 26240 20128 26246
rect 20076 26182 20128 26188
rect 20088 25838 20116 26182
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 19984 25288 20036 25294
rect 19444 25214 19656 25242
rect 19984 25230 20036 25236
rect 19432 25152 19484 25158
rect 19628 25140 19656 25214
rect 19628 25112 20024 25140
rect 19432 25094 19484 25100
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 19246 20360 19302 20369
rect 19246 20295 19248 20304
rect 19300 20295 19302 20304
rect 19248 20266 19300 20272
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19260 19009 19288 19450
rect 19352 19310 19380 24074
rect 19444 23730 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19996 23186 20024 25112
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 20088 23066 20116 25366
rect 19996 23038 20116 23066
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 23038
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 20088 22778 20116 22918
rect 20180 22778 20208 26279
rect 20272 25974 20300 26930
rect 20364 26450 20392 29446
rect 20456 29238 20484 30738
rect 20548 30734 20576 31894
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20456 28490 20484 29174
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20548 28150 20576 30670
rect 20536 28144 20588 28150
rect 20456 28092 20536 28098
rect 20456 28086 20588 28092
rect 20456 28070 20576 28086
rect 20456 27538 20484 28070
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20548 27062 20576 27814
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20444 26512 20496 26518
rect 20444 26454 20496 26460
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20272 25362 20300 25910
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20364 25242 20392 26386
rect 20272 25214 20392 25242
rect 20272 24698 20300 25214
rect 20456 24818 20484 26454
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20548 25294 20576 26318
rect 20640 25906 20668 34546
rect 20732 33998 20760 35142
rect 20824 34542 20852 35566
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 21100 34610 21128 35090
rect 21180 35012 21232 35018
rect 21180 34954 21232 34960
rect 21088 34604 21140 34610
rect 21088 34546 21140 34552
rect 20812 34536 20864 34542
rect 20812 34478 20864 34484
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20720 33040 20772 33046
rect 20720 32982 20772 32988
rect 20732 32366 20760 32982
rect 20812 32836 20864 32842
rect 20812 32778 20864 32784
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20824 32230 20852 32778
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20916 32570 20944 32710
rect 20904 32564 20956 32570
rect 20904 32506 20956 32512
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20824 31278 20852 32166
rect 20994 31784 21050 31793
rect 20994 31719 21050 31728
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20732 29034 20760 29990
rect 20824 29073 20852 30874
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20810 29064 20866 29073
rect 20720 29028 20772 29034
rect 20810 28999 20866 29008
rect 20720 28970 20772 28976
rect 20718 28656 20774 28665
rect 20718 28591 20774 28600
rect 20732 27402 20760 28591
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20732 25974 20760 26726
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20824 25838 20852 28999
rect 20916 26926 20944 30534
rect 21008 29170 21036 31719
rect 21100 30734 21128 34546
rect 21192 31754 21220 34954
rect 21284 34610 21312 35702
rect 21376 34610 21404 35770
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 21364 34604 21416 34610
rect 21364 34546 21416 34552
rect 21272 34196 21324 34202
rect 21272 34138 21324 34144
rect 21284 31890 21312 34138
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 21376 31929 21404 34002
rect 21560 33930 21588 36722
rect 22296 36378 22324 37130
rect 22376 36780 22428 36786
rect 22376 36722 22428 36728
rect 22284 36372 22336 36378
rect 22284 36314 22336 36320
rect 22296 36242 22324 36314
rect 22284 36236 22336 36242
rect 22284 36178 22336 36184
rect 22388 35834 22416 36722
rect 22468 36236 22520 36242
rect 22468 36178 22520 36184
rect 22376 35828 22428 35834
rect 22376 35770 22428 35776
rect 22480 35222 22508 36178
rect 22940 36038 22968 37130
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 26608 37120 26660 37126
rect 26608 37062 26660 37068
rect 23020 36576 23072 36582
rect 23020 36518 23072 36524
rect 23032 36174 23060 36518
rect 23020 36168 23072 36174
rect 23020 36110 23072 36116
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 22928 36032 22980 36038
rect 22928 35974 22980 35980
rect 22940 35698 22968 35974
rect 23032 35834 23060 36110
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23400 35766 23428 36110
rect 23676 36106 23704 37062
rect 23756 36848 23808 36854
rect 23756 36790 23808 36796
rect 25596 36848 25648 36854
rect 25596 36790 25648 36796
rect 23664 36100 23716 36106
rect 23664 36042 23716 36048
rect 23388 35760 23440 35766
rect 23388 35702 23440 35708
rect 23572 35760 23624 35766
rect 23572 35702 23624 35708
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 22468 35216 22520 35222
rect 22468 35158 22520 35164
rect 23400 35170 23428 35430
rect 23480 35216 23532 35222
rect 23400 35164 23480 35170
rect 23400 35158 23532 35164
rect 23400 35142 23520 35158
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22112 34746 22140 35022
rect 23020 35012 23072 35018
rect 23020 34954 23072 34960
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22376 34536 22428 34542
rect 22376 34478 22428 34484
rect 22192 34400 22244 34406
rect 22192 34342 22244 34348
rect 21548 33924 21600 33930
rect 21548 33866 21600 33872
rect 21640 33924 21692 33930
rect 21640 33866 21692 33872
rect 21560 32502 21588 33866
rect 21652 33658 21680 33866
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21652 32978 21680 33594
rect 21730 33416 21786 33425
rect 21730 33351 21786 33360
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21468 31958 21496 32166
rect 21456 31952 21508 31958
rect 21362 31920 21418 31929
rect 21272 31884 21324 31890
rect 21456 31894 21508 31900
rect 21362 31855 21418 31864
rect 21272 31826 21324 31832
rect 21376 31822 21404 31855
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 21192 31726 21312 31754
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21192 31482 21220 31622
rect 21284 31498 21312 31726
rect 21180 31476 21232 31482
rect 21284 31470 21404 31498
rect 21180 31418 21232 31424
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21284 30734 21312 31282
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 21100 28966 21128 30670
rect 21376 28994 21404 31470
rect 21456 30184 21508 30190
rect 21456 30126 21508 30132
rect 21468 30025 21496 30126
rect 21454 30016 21510 30025
rect 21454 29951 21510 29960
rect 21744 29850 21772 33351
rect 22204 33318 22232 34342
rect 22388 33998 22416 34478
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22744 34400 22796 34406
rect 22744 34342 22796 34348
rect 22572 33998 22600 34342
rect 22756 34202 22784 34342
rect 22744 34196 22796 34202
rect 22744 34138 22796 34144
rect 22652 34128 22704 34134
rect 22652 34070 22704 34076
rect 22376 33992 22428 33998
rect 22376 33934 22428 33940
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21732 29844 21784 29850
rect 21732 29786 21784 29792
rect 21638 29744 21694 29753
rect 21638 29679 21640 29688
rect 21692 29679 21694 29688
rect 21640 29650 21692 29656
rect 21928 29646 21956 32302
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 22112 30938 22140 31962
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21284 28966 21404 28994
rect 21456 29028 21508 29034
rect 21456 28970 21508 28976
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 21008 27674 21036 28154
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20548 24886 20576 25230
rect 20916 25226 20944 25638
rect 20904 25220 20956 25226
rect 20904 25162 20956 25168
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20536 24880 20588 24886
rect 20536 24822 20588 24828
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20272 24670 20484 24698
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20272 23186 20300 24006
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20364 23032 20392 23530
rect 20456 23186 20484 24670
rect 20640 23594 20668 25094
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20824 23730 20852 24210
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20272 23004 20392 23032
rect 20536 23044 20588 23050
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19444 20466 19472 21966
rect 20180 21894 20208 22578
rect 20272 22094 20300 23004
rect 20536 22986 20588 22992
rect 20548 22778 20576 22986
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20456 22658 20484 22714
rect 20456 22630 20576 22658
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20272 22066 20392 22094
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 21558
rect 20364 20618 20392 22066
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20180 20590 20392 20618
rect 19720 20482 19748 20538
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19524 20460 19576 20466
rect 19720 20454 19840 20482
rect 19524 20402 19576 20408
rect 19444 20233 19472 20402
rect 19430 20224 19486 20233
rect 19430 20159 19486 20168
rect 19536 20058 19564 20402
rect 19812 20262 19840 20454
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19720 19922 19748 20198
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19996 19786 20024 20538
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 20088 20369 20116 20470
rect 20074 20360 20130 20369
rect 20074 20295 20130 20304
rect 20180 20312 20208 20590
rect 20456 20448 20484 22170
rect 20364 20420 20484 20448
rect 20180 20284 20300 20312
rect 20074 20224 20130 20233
rect 20074 20159 20130 20168
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 19360 20116 20159
rect 20166 20088 20222 20097
rect 20166 20023 20222 20032
rect 20180 19514 20208 20023
rect 20272 19718 20300 20284
rect 20364 20262 20392 20420
rect 20548 20346 20576 22630
rect 20640 22234 20668 23122
rect 20732 22574 20760 23462
rect 20916 23118 20944 25162
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 21008 20398 21036 26930
rect 21100 26790 21128 27338
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21192 26382 21220 27610
rect 21284 26518 21312 28966
rect 21468 28626 21496 28970
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21272 26512 21324 26518
rect 21272 26454 21324 26460
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21192 25294 21220 26318
rect 21376 26042 21404 28494
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21468 26518 21496 28358
rect 21744 26926 21772 29582
rect 22204 29578 22232 33254
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22296 31346 22324 32166
rect 22388 31346 22416 33526
rect 22572 32910 22600 33934
rect 22664 33318 22692 34070
rect 23032 33998 23060 34954
rect 23400 34950 23428 35142
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23400 34474 23428 34886
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23204 34468 23256 34474
rect 23204 34410 23256 34416
rect 23388 34468 23440 34474
rect 23388 34410 23440 34416
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22572 31890 22600 31962
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22376 31340 22428 31346
rect 22376 31282 22428 31288
rect 22480 31226 22508 31622
rect 22388 31198 22508 31226
rect 22192 29572 22244 29578
rect 22192 29514 22244 29520
rect 22204 29170 22232 29514
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22112 28506 22140 28970
rect 21916 28484 21968 28490
rect 21916 28426 21968 28432
rect 22020 28478 22140 28506
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 27470 21864 28358
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21732 26920 21784 26926
rect 21732 26862 21784 26868
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21468 26217 21496 26318
rect 21454 26208 21510 26217
rect 21454 26143 21510 26152
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20456 20318 20576 20346
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20720 20324 20772 20330
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20272 19378 20300 19654
rect 20350 19408 20406 19417
rect 19536 19334 20116 19360
rect 19444 19332 20116 19334
rect 20260 19372 20312 19378
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19444 19306 19564 19332
rect 20350 19343 20406 19352
rect 20260 19314 20312 19320
rect 19246 19000 19302 19009
rect 19246 18935 19302 18944
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18984 18426 19012 18634
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 19168 16726 19196 18838
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 17066 19288 17546
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16726 19288 17002
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18432 15094 18460 15574
rect 18420 15088 18472 15094
rect 18420 15030 18472 15036
rect 18524 14346 18552 15574
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18800 14414 18828 15030
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 14074 18920 14214
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 17868 12378 17920 12384
rect 18248 12406 18368 12434
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17500 11756 17552 11762
rect 17696 11744 17724 12038
rect 17788 11830 17816 12038
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17552 11716 17724 11744
rect 17500 11698 17552 11704
rect 17328 11558 17356 11698
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17328 10810 17356 11086
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17420 10266 17448 11086
rect 17512 10690 17540 11698
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10810 17724 10950
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17788 10742 17816 11766
rect 17880 11014 17908 12378
rect 18248 12374 18276 12406
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18892 12306 18920 13874
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 17972 11354 18000 12242
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18524 11558 18552 11698
rect 18708 11626 18736 12174
rect 18984 12102 19012 14350
rect 19352 12434 19380 19246
rect 19444 17270 19472 19306
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19616 18896 19668 18902
rect 19614 18864 19616 18873
rect 19668 18864 19670 18873
rect 19614 18799 19670 18808
rect 19904 18766 19932 18906
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18222 20024 19110
rect 20074 19000 20130 19009
rect 20074 18935 20076 18944
rect 20128 18935 20130 18944
rect 20076 18906 20128 18912
rect 20272 18222 20300 19314
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19444 13954 19472 16594
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16114 20024 16934
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 14906 20116 17750
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 19996 14890 20116 14906
rect 19984 14884 20116 14890
rect 20036 14878 20116 14884
rect 19984 14826 20036 14832
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14006 20024 14214
rect 19984 14000 20036 14006
rect 19444 13926 19564 13954
rect 19984 13942 20036 13948
rect 20088 13938 20116 14878
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20180 14482 20208 14758
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19260 12406 19380 12434
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18524 11286 18552 11494
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18984 11218 19012 12038
rect 19260 11642 19288 12406
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19352 11762 19380 12310
rect 19444 11812 19472 13806
rect 19536 13258 19564 13926
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19444 11784 19564 11812
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19260 11614 19380 11642
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17776 10736 17828 10742
rect 17512 10662 17724 10690
rect 17776 10678 17828 10684
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 17696 10266 17724 10662
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17696 10130 17724 10202
rect 17788 10130 17816 10474
rect 18156 10130 18184 10678
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17604 9110 17632 9522
rect 17788 9518 17816 10066
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 8498 17172 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16684 6886 16896 6914
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 16224 5778 16252 6190
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 4690 16528 5714
rect 16684 5302 16712 6886
rect 17788 5710 17816 9114
rect 19168 8974 19196 11494
rect 19352 9178 19380 11614
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19444 11354 19472 11562
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19536 11234 19564 11784
rect 19996 11778 20024 13806
rect 20272 12238 20300 15574
rect 20364 15502 20392 19343
rect 20456 18850 20484 20318
rect 20720 20266 20772 20272
rect 20732 19854 20760 20266
rect 21008 19990 21036 20334
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 18970 20576 19314
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20456 18822 20576 18850
rect 20548 18340 20576 18822
rect 20640 18630 20668 19654
rect 21008 19310 21036 19926
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20628 18352 20680 18358
rect 20548 18312 20628 18340
rect 20628 18294 20680 18300
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20456 18086 20484 18226
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20456 15065 20484 18022
rect 20536 15496 20588 15502
rect 20534 15464 20536 15473
rect 20588 15464 20590 15473
rect 20534 15399 20590 15408
rect 20442 15056 20498 15065
rect 20442 14991 20498 15000
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20364 14822 20392 14894
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 13870 20392 14758
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20456 13716 20484 14991
rect 20640 14958 20668 18294
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20732 15366 20760 15914
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 21008 14346 21036 18702
rect 21100 18222 21128 24006
rect 21284 23798 21312 24822
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 23866 21496 24142
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21178 19408 21234 19417
rect 21178 19343 21180 19352
rect 21232 19343 21234 19352
rect 21180 19314 21232 19320
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 18426 21312 18702
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21100 14278 21128 18158
rect 21284 18086 21312 18226
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 16114 21312 18022
rect 21376 16153 21404 22918
rect 21468 22030 21496 22918
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21560 21078 21588 26726
rect 21638 26616 21694 26625
rect 21638 26551 21694 26560
rect 21652 26450 21680 26551
rect 21744 26518 21772 26862
rect 21732 26512 21784 26518
rect 21732 26454 21784 26460
rect 21822 26480 21878 26489
rect 21640 26444 21692 26450
rect 21822 26415 21878 26424
rect 21640 26386 21692 26392
rect 21638 26072 21694 26081
rect 21638 26007 21694 26016
rect 21652 23662 21680 26007
rect 21732 25968 21784 25974
rect 21732 25910 21784 25916
rect 21744 24206 21772 25910
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21640 23656 21692 23662
rect 21692 23616 21772 23644
rect 21640 23598 21692 23604
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 21362 16144 21418 16153
rect 21272 16108 21324 16114
rect 21362 16079 21418 16088
rect 21272 16050 21324 16056
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20364 13688 20484 13716
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 19444 11206 19564 11234
rect 19628 11750 20024 11778
rect 20180 11762 20208 12106
rect 20168 11756 20220 11762
rect 19444 10198 19472 11206
rect 19524 11144 19576 11150
rect 19628 11132 19656 11750
rect 20168 11698 20220 11704
rect 19984 11688 20036 11694
rect 19812 11648 19984 11676
rect 19812 11558 19840 11648
rect 19984 11630 20036 11636
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19812 11150 19840 11494
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19904 11150 19932 11290
rect 19576 11104 19656 11132
rect 19800 11144 19852 11150
rect 19524 11086 19576 11092
rect 19800 11086 19852 11092
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19812 8974 19840 9318
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18432 8498 18460 8842
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8498 19012 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8566 20024 9862
rect 20088 9042 20116 10066
rect 20364 9674 20392 13688
rect 20824 13326 20852 14214
rect 21376 13394 21404 14486
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12986 21312 13262
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20456 11354 20484 11494
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20548 11150 20576 12174
rect 20640 11558 20668 12242
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20272 9646 20392 9674
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8566 20116 8978
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17972 6866 18000 7754
rect 18248 7410 18276 8366
rect 18432 7478 18460 8434
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 7002 18276 7346
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18340 6798 18368 7278
rect 18432 6866 18460 7414
rect 18524 7410 18552 7822
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18984 7478 19012 7754
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18340 6322 18368 6734
rect 18524 6322 18552 6938
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18064 5778 18092 5850
rect 19168 5778 19196 6190
rect 19260 5914 19288 7210
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19352 5846 19380 6326
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 19352 4978 19380 5782
rect 19444 5778 19472 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20272 6914 20300 9646
rect 20548 9450 20576 11086
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9722 20760 10066
rect 20916 10062 20944 10406
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20824 8498 20852 9046
rect 20916 8634 20944 9862
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20732 7886 20760 8298
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20824 7410 20852 8434
rect 21008 7954 21036 12582
rect 21192 12442 21220 12786
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21284 12238 21312 12922
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21100 11082 21128 12174
rect 21284 11626 21312 12174
rect 21376 11898 21404 12786
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21376 10606 21404 11834
rect 21468 11150 21496 19926
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21652 17678 21680 19790
rect 21744 19446 21772 23616
rect 21836 22438 21864 26415
rect 21928 24818 21956 28426
rect 22020 27962 22048 28478
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22296 28082 22324 28358
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22020 27934 22232 27962
rect 22100 26784 22152 26790
rect 22006 26752 22062 26761
rect 22100 26726 22152 26732
rect 22006 26687 22062 26696
rect 22020 26489 22048 26687
rect 22006 26480 22062 26489
rect 22006 26415 22062 26424
rect 22020 26382 22048 26415
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 22020 25906 22048 26182
rect 22112 26081 22140 26726
rect 22098 26072 22154 26081
rect 22098 26007 22154 26016
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25158 22140 25842
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 22112 22642 22140 25094
rect 22204 23798 22232 27934
rect 22388 26246 22416 31198
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22480 29102 22508 29786
rect 22572 29646 22600 31078
rect 22664 30734 22692 33254
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22756 32774 22784 33050
rect 22848 32978 22876 33458
rect 23216 33454 23244 34410
rect 23492 33998 23520 34478
rect 23584 34202 23612 35702
rect 23676 35698 23704 36042
rect 23768 35698 23796 36790
rect 24860 36712 24912 36718
rect 24860 36654 24912 36660
rect 24872 36281 24900 36654
rect 25608 36378 25636 36790
rect 26620 36786 26648 37062
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26608 36780 26660 36786
rect 26608 36722 26660 36728
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 24952 36372 25004 36378
rect 24952 36314 25004 36320
rect 25596 36372 25648 36378
rect 25596 36314 25648 36320
rect 24858 36272 24914 36281
rect 24858 36207 24914 36216
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23664 35080 23716 35086
rect 23664 35022 23716 35028
rect 23676 34474 23704 35022
rect 23664 34468 23716 34474
rect 23664 34410 23716 34416
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23388 33924 23440 33930
rect 23388 33866 23440 33872
rect 23400 33522 23428 33866
rect 23388 33516 23440 33522
rect 23388 33458 23440 33464
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23400 32978 23428 33458
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 22744 32768 22796 32774
rect 22742 32736 22744 32745
rect 22796 32736 22798 32745
rect 22742 32671 22798 32680
rect 22848 32042 22876 32914
rect 22928 32904 22980 32910
rect 22980 32864 23060 32892
rect 22928 32846 22980 32852
rect 22848 32026 22968 32042
rect 22836 32020 22968 32026
rect 22888 32014 22968 32020
rect 22836 31962 22888 31968
rect 22940 31822 22968 32014
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 23032 31482 23060 32864
rect 23112 31952 23164 31958
rect 23112 31894 23164 31900
rect 23124 31754 23152 31894
rect 23400 31754 23428 32914
rect 23492 32570 23520 33934
rect 23572 33448 23624 33454
rect 23572 33390 23624 33396
rect 23584 32774 23612 33390
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23492 32434 23520 32506
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23584 31754 23612 32710
rect 23768 31793 23796 35634
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23860 34542 23888 35022
rect 24492 34740 24544 34746
rect 24492 34682 24544 34688
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23860 32434 23888 34138
rect 24308 34060 24360 34066
rect 24308 34002 24360 34008
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 23848 32428 23900 32434
rect 23848 32370 23900 32376
rect 23848 32224 23900 32230
rect 23848 32166 23900 32172
rect 23860 31822 23888 32166
rect 23848 31816 23900 31822
rect 23754 31784 23810 31793
rect 23124 31726 23244 31754
rect 23020 31476 23072 31482
rect 23020 31418 23072 31424
rect 22744 31136 22796 31142
rect 22744 31078 22796 31084
rect 22756 30802 22784 31078
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22744 30660 22796 30666
rect 22744 30602 22796 30608
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22664 29594 22692 29990
rect 22756 29782 22784 30602
rect 22836 30592 22888 30598
rect 22834 30560 22836 30569
rect 22888 30560 22890 30569
rect 22834 30495 22890 30504
rect 22848 30104 22876 30495
rect 23216 30258 23244 31726
rect 23388 31748 23440 31754
rect 23584 31726 23704 31754
rect 23388 31690 23440 31696
rect 23400 31346 23428 31690
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23480 31272 23532 31278
rect 23480 31214 23532 31220
rect 23388 31204 23440 31210
rect 23388 31146 23440 31152
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23308 30705 23336 30874
rect 23400 30734 23428 31146
rect 23388 30728 23440 30734
rect 23294 30696 23350 30705
rect 23388 30670 23440 30676
rect 23294 30631 23350 30640
rect 23308 30580 23336 30631
rect 23308 30552 23428 30580
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 22928 30116 22980 30122
rect 22848 30076 22928 30104
rect 22928 30058 22980 30064
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23020 29844 23072 29850
rect 23020 29786 23072 29792
rect 22744 29776 22796 29782
rect 22744 29718 22796 29724
rect 22664 29566 22784 29594
rect 22652 29504 22704 29510
rect 22756 29481 22784 29566
rect 22652 29446 22704 29452
rect 22742 29472 22798 29481
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22192 23792 22244 23798
rect 22192 23734 22244 23740
rect 22204 23050 22232 23734
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22296 22778 22324 23258
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22480 22642 22508 27270
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22020 21010 22048 22374
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22112 20890 22140 22578
rect 22374 21992 22430 22001
rect 22374 21927 22430 21936
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22020 20874 22140 20890
rect 22020 20868 22152 20874
rect 22020 20862 22100 20868
rect 22020 20058 22048 20862
rect 22100 20810 22152 20816
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22008 19848 22060 19854
rect 22006 19816 22008 19825
rect 22060 19816 22062 19825
rect 21916 19780 21968 19786
rect 22006 19751 22062 19760
rect 21916 19722 21968 19728
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21652 16658 21680 17614
rect 21928 17610 21956 19722
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 18426 22048 18702
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22112 18193 22140 18226
rect 22098 18184 22154 18193
rect 22098 18119 22154 18128
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 16250 21588 16526
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21652 15502 21680 16594
rect 21928 16590 21956 17546
rect 22204 17218 22232 20946
rect 22296 19786 22324 20946
rect 22388 20942 22416 21927
rect 22480 21010 22508 22578
rect 22572 22094 22600 28426
rect 22664 27470 22692 29446
rect 22742 29407 22798 29416
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22664 26994 22692 27406
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22756 26874 22784 29407
rect 22926 29336 22982 29345
rect 22926 29271 22982 29280
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22848 28150 22876 28358
rect 22836 28144 22888 28150
rect 22836 28086 22888 28092
rect 22836 27940 22888 27946
rect 22836 27882 22888 27888
rect 22664 26846 22784 26874
rect 22664 24274 22692 26846
rect 22848 26382 22876 27882
rect 22940 27606 22968 29271
rect 23032 29034 23060 29786
rect 23124 29646 23152 29990
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23020 29028 23072 29034
rect 23020 28970 23072 28976
rect 22928 27600 22980 27606
rect 22928 27542 22980 27548
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 22940 26246 22968 26930
rect 23032 26790 23060 28970
rect 23110 28656 23166 28665
rect 23110 28591 23166 28600
rect 23124 28558 23152 28591
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23216 28082 23244 30194
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23308 29850 23336 30126
rect 23400 29850 23428 30552
rect 23296 29844 23348 29850
rect 23296 29786 23348 29792
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23308 28490 23336 29582
rect 23400 29306 23428 29582
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23388 29096 23440 29102
rect 23492 29073 23520 31214
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23584 30258 23612 30670
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23570 30016 23626 30025
rect 23570 29951 23626 29960
rect 23388 29038 23440 29044
rect 23478 29064 23534 29073
rect 23296 28484 23348 28490
rect 23296 28426 23348 28432
rect 23296 28144 23348 28150
rect 23296 28086 23348 28092
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23124 27334 23152 28018
rect 23204 27600 23256 27606
rect 23204 27542 23256 27548
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23020 26580 23072 26586
rect 23020 26522 23072 26528
rect 22928 26240 22980 26246
rect 23032 26217 23060 26522
rect 22928 26182 22980 26188
rect 23018 26208 23074 26217
rect 23018 26143 23074 26152
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22756 24886 22784 25910
rect 23124 25294 23152 27270
rect 23216 26994 23244 27542
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23308 26874 23336 28086
rect 23216 26846 23336 26874
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 22744 24880 22796 24886
rect 22744 24822 22796 24828
rect 23110 24848 23166 24857
rect 23110 24783 23112 24792
rect 23164 24783 23166 24792
rect 23112 24754 23164 24760
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22664 22982 22692 24210
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 23322 22876 24006
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22572 22066 22692 22094
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22572 20534 22600 21966
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22480 20058 22508 20334
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22112 17190 22232 17218
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 15026 21680 15438
rect 21824 15428 21876 15434
rect 21928 15416 21956 16526
rect 22006 16144 22062 16153
rect 22006 16079 22062 16088
rect 22020 15502 22048 16079
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21876 15388 21956 15416
rect 21824 15370 21876 15376
rect 21928 15094 21956 15388
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21652 14414 21680 14962
rect 21928 14414 21956 15030
rect 22006 14512 22062 14521
rect 22006 14447 22062 14456
rect 22020 14414 22048 14447
rect 21640 14408 21692 14414
rect 21732 14408 21784 14414
rect 21640 14350 21692 14356
rect 21730 14376 21732 14385
rect 21916 14408 21968 14414
rect 21784 14376 21786 14385
rect 21916 14350 21968 14356
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21730 14311 21786 14320
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21560 12238 21588 13262
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21652 11694 21680 12582
rect 21744 11762 21772 13330
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21744 11218 21772 11698
rect 21928 11354 21956 12650
rect 22020 12238 22048 13262
rect 22112 12374 22140 17190
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12850 22232 13126
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21468 10062 21496 11086
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21100 9042 21128 9522
rect 21468 9518 21496 9998
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 22020 9042 22048 12174
rect 22296 11370 22324 19314
rect 22480 18290 22508 19994
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22388 17814 22416 18226
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 22480 13530 22508 18226
rect 22572 17270 22600 20470
rect 22664 19854 22692 22066
rect 22756 21690 22784 22578
rect 23032 22098 23060 24142
rect 23124 23730 23152 24754
rect 23216 24410 23244 26846
rect 23400 26466 23428 29038
rect 23478 28999 23534 29008
rect 23492 28558 23520 28999
rect 23480 28552 23532 28558
rect 23480 28494 23532 28500
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23492 27538 23520 27814
rect 23584 27606 23612 29951
rect 23676 29306 23704 31726
rect 23848 31758 23900 31764
rect 24030 31784 24086 31793
rect 23754 31719 23810 31728
rect 24030 31719 24086 31728
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23860 31260 23888 31418
rect 23940 31272 23992 31278
rect 23860 31232 23940 31260
rect 23768 29578 23796 31214
rect 23860 30734 23888 31232
rect 23940 31214 23992 31220
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 24044 29782 24072 31719
rect 24032 29776 24084 29782
rect 24032 29718 24084 29724
rect 23756 29572 23808 29578
rect 23756 29514 23808 29520
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23676 27674 23704 29242
rect 23768 29170 23796 29514
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23860 28694 23888 29106
rect 23848 28688 23900 28694
rect 23848 28630 23900 28636
rect 23860 27690 23888 28630
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23768 27662 23888 27690
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23308 26438 23428 26466
rect 23308 25906 23336 26438
rect 23584 26382 23612 26794
rect 23662 26616 23718 26625
rect 23662 26551 23664 26560
rect 23716 26551 23718 26560
rect 23664 26522 23716 26528
rect 23676 26382 23704 26522
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23308 24818 23336 25706
rect 23400 24818 23428 26318
rect 23584 25294 23612 26318
rect 23768 25906 23796 27662
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 23952 26994 23980 27338
rect 23940 26988 23992 26994
rect 23940 26930 23992 26936
rect 23848 26444 23900 26450
rect 23848 26386 23900 26392
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23216 23882 23244 24210
rect 23308 24070 23336 24754
rect 23400 24274 23428 24754
rect 23478 24712 23534 24721
rect 23478 24647 23534 24656
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23388 24132 23440 24138
rect 23388 24074 23440 24080
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23216 23854 23336 23882
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23202 22128 23258 22137
rect 23020 22092 23072 22098
rect 23202 22063 23258 22072
rect 23020 22034 23072 22040
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22756 20466 22784 21626
rect 23216 20942 23244 22063
rect 23308 21962 23336 23854
rect 23400 23730 23428 24074
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23492 23594 23520 24647
rect 23860 24206 23888 26386
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23492 23497 23520 23530
rect 23478 23488 23534 23497
rect 23478 23423 23534 23432
rect 23952 22166 23980 26930
rect 24044 26518 24072 29718
rect 24136 28558 24164 32506
rect 24320 31890 24348 34002
rect 24504 32434 24532 34682
rect 24596 33844 24624 36110
rect 24860 36100 24912 36106
rect 24860 36042 24912 36048
rect 24872 35222 24900 36042
rect 24860 35216 24912 35222
rect 24860 35158 24912 35164
rect 24872 34950 24900 35158
rect 24964 35057 24992 36314
rect 26160 36242 26188 36654
rect 26344 36242 26372 36722
rect 26424 36576 26476 36582
rect 26424 36518 26476 36524
rect 26436 36242 26464 36518
rect 27172 36378 27200 37198
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 26148 36236 26200 36242
rect 26148 36178 26200 36184
rect 26332 36236 26384 36242
rect 26332 36178 26384 36184
rect 26424 36236 26476 36242
rect 26424 36178 26476 36184
rect 27724 36106 27752 37198
rect 31024 37188 31076 37194
rect 31024 37130 31076 37136
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 28540 37120 28592 37126
rect 28540 37062 28592 37068
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28276 36378 28304 36722
rect 28264 36372 28316 36378
rect 28264 36314 28316 36320
rect 27712 36100 27764 36106
rect 27712 36042 27764 36048
rect 25228 35692 25280 35698
rect 25228 35634 25280 35640
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25044 35488 25096 35494
rect 25044 35430 25096 35436
rect 24950 35048 25006 35057
rect 24950 34983 25006 34992
rect 25056 34950 25084 35430
rect 25148 35086 25176 35566
rect 25240 35290 25268 35634
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 25228 35284 25280 35290
rect 25228 35226 25280 35232
rect 25240 35154 25268 35226
rect 25516 35222 25544 35566
rect 26056 35556 26108 35562
rect 26056 35498 26108 35504
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 25504 35216 25556 35222
rect 25504 35158 25556 35164
rect 25228 35148 25280 35154
rect 25228 35090 25280 35096
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24676 34400 24728 34406
rect 24676 34342 24728 34348
rect 24688 33998 24716 34342
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24596 33816 24716 33844
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24308 31884 24360 31890
rect 24308 31826 24360 31832
rect 24216 30728 24268 30734
rect 24216 30670 24268 30676
rect 24228 30394 24256 30670
rect 24216 30388 24268 30394
rect 24216 30330 24268 30336
rect 24320 30258 24348 31826
rect 24412 31804 24440 32370
rect 24492 31816 24544 31822
rect 24412 31776 24492 31804
rect 24492 31758 24544 31764
rect 24504 31346 24532 31758
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 24308 30252 24360 30258
rect 24308 30194 24360 30200
rect 24320 29753 24348 30194
rect 24306 29744 24362 29753
rect 24306 29679 24362 29688
rect 24320 29238 24348 29679
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 24412 28994 24440 31214
rect 24504 30326 24532 31282
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24412 28966 24532 28994
rect 24124 28552 24176 28558
rect 24124 28494 24176 28500
rect 24124 28144 24176 28150
rect 24124 28086 24176 28092
rect 24136 27606 24164 28086
rect 24124 27600 24176 27606
rect 24124 27542 24176 27548
rect 24136 26994 24164 27542
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 24136 25158 24164 26930
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24136 24410 24164 25094
rect 24320 24970 24348 25434
rect 24504 25362 24532 28966
rect 24596 27130 24624 32846
rect 24688 32434 24716 33816
rect 24872 33318 24900 34886
rect 25148 34610 25176 35022
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 24952 34536 25004 34542
rect 24952 34478 25004 34484
rect 24964 34134 24992 34478
rect 24952 34128 25004 34134
rect 24952 34070 25004 34076
rect 25056 33998 25084 34546
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24768 31476 24820 31482
rect 24768 31418 24820 31424
rect 24780 30190 24808 31418
rect 24872 31346 24900 33254
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24768 30184 24820 30190
rect 24768 30126 24820 30132
rect 24964 29306 24992 32914
rect 25056 31754 25084 33934
rect 25148 33454 25176 34546
rect 25240 34406 25268 35090
rect 25976 35057 26004 35226
rect 25962 35048 26018 35057
rect 25504 35012 25556 35018
rect 26068 35018 26096 35498
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 25962 34983 26018 34992
rect 26056 35012 26108 35018
rect 25504 34954 25556 34960
rect 26056 34954 26108 34960
rect 25228 34400 25280 34406
rect 25228 34342 25280 34348
rect 25240 33930 25268 34342
rect 25228 33924 25280 33930
rect 25228 33866 25280 33872
rect 25136 33448 25188 33454
rect 25136 33390 25188 33396
rect 25240 33318 25268 33866
rect 25228 33312 25280 33318
rect 25228 33254 25280 33260
rect 25410 33280 25466 33289
rect 25410 33215 25466 33224
rect 25424 33046 25452 33215
rect 25412 33040 25464 33046
rect 25412 32982 25464 32988
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25240 32570 25268 32846
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25136 32224 25188 32230
rect 25240 32178 25268 32302
rect 25188 32172 25268 32178
rect 25136 32166 25268 32172
rect 25148 32150 25268 32166
rect 25148 31754 25176 32150
rect 25044 31748 25096 31754
rect 25148 31726 25268 31754
rect 25044 31690 25096 31696
rect 25056 31498 25084 31690
rect 25056 31470 25176 31498
rect 25148 30802 25176 31470
rect 25240 31142 25268 31726
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 25412 30932 25464 30938
rect 25412 30874 25464 30880
rect 25136 30796 25188 30802
rect 25136 30738 25188 30744
rect 25424 30258 25452 30874
rect 25516 30734 25544 34954
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25608 33998 25636 34886
rect 25596 33992 25648 33998
rect 25596 33934 25648 33940
rect 25608 33590 25636 33934
rect 25700 33930 25728 34886
rect 26160 34678 26188 35090
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26148 34672 26200 34678
rect 26148 34614 26200 34620
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 25688 33924 25740 33930
rect 25688 33866 25740 33872
rect 25700 33658 25728 33866
rect 25688 33652 25740 33658
rect 25688 33594 25740 33600
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25608 30410 25636 33526
rect 26068 33402 26096 34546
rect 26160 33522 26188 34614
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26528 33590 26556 33866
rect 26620 33658 26648 35022
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26896 34678 26924 34954
rect 27264 34746 27292 35634
rect 27724 35630 27752 36042
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27344 35216 27396 35222
rect 27344 35158 27396 35164
rect 27252 34740 27304 34746
rect 27252 34682 27304 34688
rect 26884 34672 26936 34678
rect 26884 34614 26936 34620
rect 26700 34060 26752 34066
rect 26700 34002 26752 34008
rect 26608 33652 26660 33658
rect 26608 33594 26660 33600
rect 26516 33584 26568 33590
rect 26516 33526 26568 33532
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26332 33448 26384 33454
rect 26068 33396 26332 33402
rect 26068 33390 26384 33396
rect 25780 33380 25832 33386
rect 25780 33322 25832 33328
rect 26068 33374 26372 33390
rect 25688 33108 25740 33114
rect 25688 33050 25740 33056
rect 25700 32337 25728 33050
rect 25686 32328 25742 32337
rect 25686 32263 25742 32272
rect 25688 31952 25740 31958
rect 25688 31894 25740 31900
rect 25700 31822 25728 31894
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25700 31482 25728 31758
rect 25792 31634 25820 33322
rect 25872 33312 25924 33318
rect 25872 33254 25924 33260
rect 25884 31822 25912 33254
rect 26068 32842 26096 33374
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26056 32836 26108 32842
rect 26056 32778 26108 32784
rect 26068 32434 26096 32778
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26160 31958 26188 32710
rect 26252 32434 26280 32846
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 26148 31952 26200 31958
rect 26148 31894 26200 31900
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25792 31606 26096 31634
rect 25688 31476 25740 31482
rect 25688 31418 25740 31424
rect 25872 31476 25924 31482
rect 25872 31418 25924 31424
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 25516 30382 25636 30410
rect 25516 30326 25544 30382
rect 25504 30320 25556 30326
rect 25700 30274 25728 31282
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25792 30870 25820 31078
rect 25884 30938 25912 31418
rect 25872 30932 25924 30938
rect 25872 30874 25924 30880
rect 25780 30864 25832 30870
rect 25780 30806 25832 30812
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25504 30262 25556 30268
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24780 28218 24808 28426
rect 24872 28218 24900 28970
rect 24964 28694 24992 29106
rect 25044 29096 25096 29102
rect 25042 29064 25044 29073
rect 25096 29064 25098 29073
rect 25042 28999 25098 29008
rect 25044 28960 25096 28966
rect 25044 28902 25096 28908
rect 25056 28694 25084 28902
rect 24952 28688 25004 28694
rect 24952 28630 25004 28636
rect 25044 28688 25096 28694
rect 25044 28630 25096 28636
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24860 28212 24912 28218
rect 24860 28154 24912 28160
rect 25056 28082 25084 28358
rect 25148 28150 25176 29446
rect 25332 29238 25360 30126
rect 25412 30116 25464 30122
rect 25412 30058 25464 30064
rect 25320 29232 25372 29238
rect 25320 29174 25372 29180
rect 25332 29102 25360 29174
rect 25228 29096 25280 29102
rect 25226 29064 25228 29073
rect 25320 29096 25372 29102
rect 25280 29064 25282 29073
rect 25320 29038 25372 29044
rect 25226 28999 25282 29008
rect 25136 28144 25188 28150
rect 25136 28086 25188 28092
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24780 26994 24808 27270
rect 24872 26994 24900 27474
rect 24964 27130 24992 27950
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24872 26858 24900 26930
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24952 26852 25004 26858
rect 24952 26794 25004 26800
rect 24964 26761 24992 26794
rect 25056 26790 25084 28018
rect 25240 28014 25268 28999
rect 25424 28082 25452 30058
rect 25516 29170 25544 30262
rect 25608 30258 25728 30274
rect 25596 30252 25728 30258
rect 25648 30246 25728 30252
rect 25596 30194 25648 30200
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25608 28966 25636 30194
rect 25792 29850 25820 30670
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25688 29300 25740 29306
rect 25688 29242 25740 29248
rect 25700 29102 25728 29242
rect 25688 29096 25740 29102
rect 25688 29038 25740 29044
rect 25596 28960 25648 28966
rect 25596 28902 25648 28908
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25792 27538 25820 29786
rect 25780 27532 25832 27538
rect 25780 27474 25832 27480
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 25148 26994 25176 27270
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25044 26784 25096 26790
rect 24950 26752 25006 26761
rect 25044 26726 25096 26732
rect 24950 26687 25006 26696
rect 25056 26602 25084 26726
rect 24964 26574 25084 26602
rect 24964 26382 24992 26574
rect 25148 26382 25176 26930
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 24676 26308 24728 26314
rect 24676 26250 24728 26256
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 24320 24954 24440 24970
rect 24308 24948 24440 24954
rect 24360 24942 24440 24948
rect 24308 24890 24360 24896
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24320 24410 24348 24754
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24320 23118 24348 24346
rect 24412 24274 24440 24942
rect 24400 24268 24452 24274
rect 24400 24210 24452 24216
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24504 22642 24532 25298
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 24596 23662 24624 24754
rect 24688 24206 24716 26250
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24872 25430 24900 25774
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24964 25226 24992 26318
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24964 24818 24992 25162
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24780 24070 24808 24686
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22848 18154 22876 18294
rect 22836 18148 22888 18154
rect 22836 18090 22888 18096
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22756 16794 22784 16934
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22756 16590 22784 16730
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22756 16182 22784 16526
rect 22940 16266 22968 20810
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23124 20534 23152 20742
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23124 19378 23152 19654
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 22848 16238 22968 16266
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22388 12850 22416 13194
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12986 22508 13126
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22480 12850 22508 12922
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22572 11762 22600 16118
rect 22848 12434 22876 16238
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22940 15502 22968 16118
rect 23032 16046 23060 19314
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23124 17678 23152 18226
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17066 23152 17614
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22664 12406 22876 12434
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22296 11342 22508 11370
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 22112 10606 22140 10950
rect 22204 10674 22232 11086
rect 22296 10742 22324 11222
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10742 22416 10950
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22204 10266 22232 10610
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22480 9654 22508 11342
rect 22572 9722 22600 11698
rect 22664 10538 22692 12406
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22480 8906 22508 9590
rect 22572 9586 22600 9658
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20996 7948 21048 7954
rect 20916 7908 20996 7936
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20916 7342 20944 7908
rect 20996 7890 21048 7896
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7546 21128 7822
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20364 7002 20392 7142
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20088 6886 20300 6914
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19444 5166 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19536 4978 19564 5102
rect 19352 4950 19564 4978
rect 20088 4826 20116 6886
rect 20364 6322 20392 6938
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6458 20668 6734
rect 21284 6730 21312 8366
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 7886 21588 8230
rect 22940 8090 22968 15438
rect 23124 14822 23152 16186
rect 23216 15348 23244 19858
rect 23308 19378 23336 21898
rect 23584 21350 23612 21966
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23386 20632 23442 20641
rect 23386 20567 23442 20576
rect 23400 19854 23428 20567
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23584 19378 23612 21286
rect 24504 20942 24532 21422
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24596 20466 24624 22714
rect 24688 22642 24716 23190
rect 24780 22778 24808 23666
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24688 21350 24716 22578
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24780 21350 24808 22510
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24872 21486 24900 21626
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24766 21176 24822 21185
rect 24766 21111 24822 21120
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24780 20058 24808 21111
rect 24964 20942 24992 23054
rect 25056 22438 25084 26318
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25148 25294 25176 25842
rect 25332 25498 25360 27406
rect 25412 27396 25464 27402
rect 25412 27338 25464 27344
rect 25504 27396 25556 27402
rect 25504 27338 25556 27344
rect 25424 27033 25452 27338
rect 25516 27062 25544 27338
rect 25504 27056 25556 27062
rect 25410 27024 25466 27033
rect 25504 26998 25556 27004
rect 25410 26959 25466 26968
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25148 24750 25176 25230
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25228 24336 25280 24342
rect 25228 24278 25280 24284
rect 25136 23588 25188 23594
rect 25136 23530 25188 23536
rect 25044 22432 25096 22438
rect 25044 22374 25096 22380
rect 25148 22234 25176 23530
rect 25240 23050 25268 24278
rect 25332 23202 25360 25434
rect 25504 25424 25556 25430
rect 25504 25366 25556 25372
rect 25516 23610 25544 25366
rect 25688 24880 25740 24886
rect 25688 24822 25740 24828
rect 25516 23582 25636 23610
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 25332 23174 25452 23202
rect 25424 23118 25452 23174
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 25056 21418 25084 21830
rect 25044 21412 25096 21418
rect 25044 21354 25096 21360
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 20398 24900 20742
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24400 19236 24452 19242
rect 24400 19178 24452 19184
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 23308 18290 23336 18838
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23584 18290 23612 18702
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23308 17678 23336 18226
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23296 17264 23348 17270
rect 23348 17212 23428 17218
rect 23296 17206 23428 17212
rect 23308 17190 23428 17206
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23308 16522 23336 17070
rect 23400 16658 23428 17190
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 15502 23336 16458
rect 23400 15978 23428 16594
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23216 15320 23428 15348
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23216 8022 23244 14962
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23308 13530 23336 13738
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23400 8566 23428 15320
rect 23584 15026 23612 18226
rect 23676 17270 23704 18294
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24228 17882 24256 18158
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24320 17678 24348 17818
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 23756 17604 23808 17610
rect 23808 17564 23888 17592
rect 23756 17546 23808 17552
rect 23860 17270 23888 17564
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 15162 23888 16390
rect 24044 15978 24072 17138
rect 24412 16402 24440 19178
rect 24504 18766 24532 19178
rect 24596 18970 24624 19314
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24688 18698 24716 19858
rect 24780 19854 24808 19994
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24688 18358 24716 18634
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24780 18290 24808 19110
rect 24872 18426 24900 20334
rect 24964 20330 24992 20878
rect 25056 20466 25084 20878
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17678 24624 18022
rect 24780 17678 24808 18226
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24872 17746 24900 18158
rect 24964 18086 24992 20266
rect 25056 20058 25084 20402
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24768 17672 24820 17678
rect 25148 17626 25176 22170
rect 25332 22098 25360 22918
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25228 22024 25280 22030
rect 25226 21992 25228 22001
rect 25280 21992 25282 22001
rect 25226 21927 25282 21936
rect 24768 17614 24820 17620
rect 24596 17202 24624 17614
rect 25056 17598 25176 17626
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24412 16374 24624 16402
rect 24398 16280 24454 16289
rect 24398 16215 24454 16224
rect 24412 16182 24440 16215
rect 24400 16176 24452 16182
rect 24306 16144 24362 16153
rect 24400 16118 24452 16124
rect 24306 16079 24362 16088
rect 24032 15972 24084 15978
rect 24032 15914 24084 15920
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23480 14272 23532 14278
rect 23532 14232 23612 14260
rect 23480 14214 23532 14220
rect 23584 13977 23612 14232
rect 23570 13968 23626 13977
rect 23480 13932 23532 13938
rect 23570 13903 23626 13912
rect 23756 13932 23808 13938
rect 23480 13874 23532 13880
rect 23492 13326 23520 13874
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23480 12844 23532 12850
rect 23584 12832 23612 13903
rect 23756 13874 23808 13880
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13394 23704 13670
rect 23768 13530 23796 13874
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23676 12986 23704 13330
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23952 12850 23980 14350
rect 24044 13938 24072 15914
rect 24122 15056 24178 15065
rect 24122 14991 24124 15000
rect 24176 14991 24178 15000
rect 24124 14962 24176 14968
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24044 13326 24072 13874
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23532 12804 23612 12832
rect 23940 12844 23992 12850
rect 23480 12786 23532 12792
rect 23940 12786 23992 12792
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21560 6798 21588 7822
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 22020 7546 22048 7754
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21272 6724 21324 6730
rect 21272 6666 21324 6672
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 21100 6322 21128 6666
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21468 6390 21496 6598
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21652 6322 21680 6598
rect 22112 6390 22140 7346
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 22098 6216 22154 6225
rect 22098 6151 22154 6160
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20732 5234 20760 5714
rect 21008 5710 21036 6054
rect 22112 5914 22140 6151
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22204 5778 22232 6734
rect 23204 6724 23256 6730
rect 23204 6666 23256 6672
rect 23216 6458 23244 6666
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 22204 5166 22232 5714
rect 23492 5302 23520 12786
rect 24136 10282 24164 14010
rect 24228 13938 24256 14214
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24228 13394 24256 13874
rect 24320 13870 24348 16079
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15026 24440 15846
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24412 14618 24440 14962
rect 24504 14822 24532 15370
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24412 14414 24440 14554
rect 24504 14414 24532 14758
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24492 13796 24544 13802
rect 24492 13738 24544 13744
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24504 13326 24532 13738
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24596 12306 24624 16374
rect 25056 16114 25084 17598
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25148 17202 25176 17478
rect 25240 17270 25268 21927
rect 25516 20233 25544 23462
rect 25608 22982 25636 23582
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25700 22642 25728 24822
rect 25792 24274 25820 27474
rect 25884 26586 25912 30874
rect 25976 30394 26004 31418
rect 26068 30734 26096 31606
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 25964 30388 26016 30394
rect 25964 30330 26016 30336
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 25976 28218 26004 30194
rect 26068 29102 26096 30670
rect 26160 30190 26188 31894
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26252 30870 26280 31282
rect 26344 30938 26372 31282
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26240 30864 26292 30870
rect 26240 30806 26292 30812
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 26424 29776 26476 29782
rect 26424 29718 26476 29724
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 26068 28626 26096 29038
rect 26252 29034 26280 29582
rect 26240 29028 26292 29034
rect 26240 28970 26292 28976
rect 26436 28994 26464 29718
rect 26528 29345 26556 33526
rect 26712 32910 26740 34002
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26700 32904 26752 32910
rect 26700 32846 26752 32852
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26620 29594 26648 32710
rect 26700 32020 26752 32026
rect 26700 31962 26752 31968
rect 26712 30666 26740 31962
rect 26700 30660 26752 30666
rect 26700 30602 26752 30608
rect 26620 29566 26740 29594
rect 26514 29336 26570 29345
rect 26514 29271 26570 29280
rect 26436 28966 26648 28994
rect 26056 28620 26108 28626
rect 26056 28562 26108 28568
rect 25964 28212 26016 28218
rect 25964 28154 26016 28160
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27062 26188 27406
rect 26252 27334 26280 28018
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 26344 26518 26372 26726
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26252 25294 26280 25978
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 25964 25152 26016 25158
rect 25964 25094 26016 25100
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25872 22432 25924 22438
rect 25872 22374 25924 22380
rect 25884 22030 25912 22374
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25608 20466 25636 21490
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25502 20224 25558 20233
rect 25502 20159 25558 20168
rect 25516 19310 25544 20159
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25228 17264 25280 17270
rect 25228 17206 25280 17212
rect 25332 17202 25360 18022
rect 25608 17814 25636 18226
rect 25596 17808 25648 17814
rect 25596 17750 25648 17756
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25700 16250 25728 21830
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25688 16244 25740 16250
rect 25688 16186 25740 16192
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 25056 15502 25084 15914
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 24872 15162 24900 15438
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24872 13870 24900 15098
rect 25056 14958 25084 15438
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24964 14482 24992 14894
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24964 14278 24992 14418
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24860 13864 24912 13870
rect 24780 13812 24860 13818
rect 24780 13806 24912 13812
rect 24780 13790 24900 13806
rect 24780 13258 24808 13790
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 25240 11898 25268 15846
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25424 15026 25452 15302
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25608 14618 25636 14962
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25332 14385 25360 14418
rect 25318 14376 25374 14385
rect 25318 14311 25374 14320
rect 25596 14000 25648 14006
rect 25594 13968 25596 13977
rect 25648 13968 25650 13977
rect 25700 13938 25728 16050
rect 25594 13903 25650 13912
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25608 12850 25636 13670
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 24950 11384 25006 11393
rect 24950 11319 25006 11328
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24136 10254 24256 10282
rect 24688 10266 24716 10610
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23768 6662 23796 7482
rect 23940 7472 23992 7478
rect 23940 7414 23992 7420
rect 23952 7002 23980 7414
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23952 6458 23980 6938
rect 24136 6866 24164 7142
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24136 6390 24164 6802
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24228 6322 24256 10254
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24872 8974 24900 11018
rect 24964 8974 24992 11319
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25148 10062 25176 10406
rect 25240 10130 25268 11834
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25240 9654 25268 10066
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25332 9602 25360 12242
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 10470 25544 11018
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25608 9654 25636 12038
rect 25686 11384 25742 11393
rect 25686 11319 25688 11328
rect 25740 11319 25742 11328
rect 25688 11290 25740 11296
rect 25792 11286 25820 21286
rect 25976 16182 26004 25094
rect 26252 24993 26280 25230
rect 26238 24984 26294 24993
rect 26238 24919 26294 24928
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26160 24342 26188 24686
rect 26436 24682 26464 27814
rect 26620 27470 26648 28966
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26516 26580 26568 26586
rect 26516 26522 26568 26528
rect 26528 25294 26556 26522
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26148 24336 26200 24342
rect 26148 24278 26200 24284
rect 26252 23798 26280 24618
rect 26240 23792 26292 23798
rect 26240 23734 26292 23740
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 26160 22642 26188 23598
rect 26252 23322 26280 23734
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26252 22710 26280 23258
rect 26240 22704 26292 22710
rect 26240 22646 26292 22652
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26160 21010 26188 21966
rect 26148 21004 26200 21010
rect 26148 20946 26200 20952
rect 26252 19990 26280 22510
rect 26424 22500 26476 22506
rect 26424 22442 26476 22448
rect 26436 21690 26464 22442
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26424 20936 26476 20942
rect 26422 20904 26424 20913
rect 26476 20904 26478 20913
rect 26422 20839 26478 20848
rect 26528 20058 26556 22578
rect 26712 22094 26740 29566
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26804 26314 26832 27338
rect 26792 26308 26844 26314
rect 26792 26250 26844 26256
rect 26896 25294 26924 33934
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 27172 31822 27200 33390
rect 27250 31920 27306 31929
rect 27250 31855 27306 31864
rect 27264 31822 27292 31855
rect 27160 31816 27212 31822
rect 27160 31758 27212 31764
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 27068 31748 27120 31754
rect 27068 31690 27120 31696
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 26988 29102 27016 31282
rect 27080 30734 27108 31690
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27068 29504 27120 29510
rect 27066 29472 27068 29481
rect 27120 29472 27122 29481
rect 27066 29407 27122 29416
rect 27172 29306 27200 31758
rect 27264 31346 27292 31758
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 27252 30660 27304 30666
rect 27252 30602 27304 30608
rect 27264 30394 27292 30602
rect 27252 30388 27304 30394
rect 27252 30330 27304 30336
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27068 29232 27120 29238
rect 27068 29174 27120 29180
rect 26976 29096 27028 29102
rect 26976 29038 27028 29044
rect 26988 27946 27016 29038
rect 27080 28558 27108 29174
rect 27264 29170 27292 29514
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27252 29164 27304 29170
rect 27252 29106 27304 29112
rect 27172 28762 27200 29106
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 27252 28484 27304 28490
rect 27252 28426 27304 28432
rect 26976 27940 27028 27946
rect 26976 27882 27028 27888
rect 27068 27940 27120 27946
rect 27068 27882 27120 27888
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26896 24206 26924 25230
rect 27080 24256 27108 27882
rect 27160 27872 27212 27878
rect 27160 27814 27212 27820
rect 27172 27130 27200 27814
rect 27264 27334 27292 28426
rect 27356 28082 27384 35158
rect 27620 34536 27672 34542
rect 27620 34478 27672 34484
rect 27632 33930 27660 34478
rect 27620 33924 27672 33930
rect 27620 33866 27672 33872
rect 27436 33652 27488 33658
rect 27436 33594 27488 33600
rect 27448 30326 27476 33594
rect 27632 33046 27660 33866
rect 27620 33040 27672 33046
rect 27620 32982 27672 32988
rect 27528 30864 27580 30870
rect 27528 30806 27580 30812
rect 27540 30734 27568 30806
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27528 30592 27580 30598
rect 27528 30534 27580 30540
rect 27436 30320 27488 30326
rect 27436 30262 27488 30268
rect 27436 30184 27488 30190
rect 27436 30126 27488 30132
rect 27448 29646 27476 30126
rect 27436 29640 27488 29646
rect 27436 29582 27488 29588
rect 27448 28490 27476 29582
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 27344 28076 27396 28082
rect 27344 28018 27396 28024
rect 27436 28008 27488 28014
rect 27436 27950 27488 27956
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 27264 25294 27292 27270
rect 27356 26994 27384 27406
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27448 26926 27476 27950
rect 27540 27878 27568 30534
rect 27632 30258 27660 32982
rect 27724 32473 27752 35566
rect 28080 34128 28132 34134
rect 28080 34070 28132 34076
rect 27710 32464 27766 32473
rect 27710 32399 27766 32408
rect 27896 32428 27948 32434
rect 27896 32370 27948 32376
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 27712 32360 27764 32366
rect 27712 32302 27764 32308
rect 27724 31754 27752 32302
rect 27908 31890 27936 32370
rect 28000 32298 28028 32370
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 28000 31822 28028 32234
rect 27988 31816 28040 31822
rect 27988 31758 28040 31764
rect 27724 31726 27936 31754
rect 27804 31136 27856 31142
rect 27804 31078 27856 31084
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27528 27872 27580 27878
rect 27528 27814 27580 27820
rect 27632 27713 27660 28358
rect 27618 27704 27674 27713
rect 27618 27639 27674 27648
rect 27724 27470 27752 30330
rect 27816 28150 27844 31078
rect 27908 28626 27936 31726
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28000 29238 28028 31282
rect 27988 29232 28040 29238
rect 27988 29174 28040 29180
rect 27896 28620 27948 28626
rect 27896 28562 27948 28568
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 27896 28212 27948 28218
rect 27896 28154 27948 28160
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27816 27606 27844 28086
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27632 26994 27660 27066
rect 27724 27033 27752 27406
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27710 27024 27766 27033
rect 27620 26988 27672 26994
rect 27710 26959 27766 26968
rect 27620 26930 27672 26936
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27632 25974 27660 26930
rect 27712 26512 27764 26518
rect 27712 26454 27764 26460
rect 27620 25968 27672 25974
rect 27620 25910 27672 25916
rect 27724 25906 27752 26454
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27252 25288 27304 25294
rect 27252 25230 27304 25236
rect 27540 24993 27568 25638
rect 27724 25430 27752 25842
rect 27712 25424 27764 25430
rect 27712 25366 27764 25372
rect 27526 24984 27582 24993
rect 27526 24919 27582 24928
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27632 24410 27660 24550
rect 27620 24404 27672 24410
rect 27620 24346 27672 24352
rect 27080 24228 27292 24256
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26896 23254 26924 24142
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 26884 23248 26936 23254
rect 26884 23190 26936 23196
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 26792 22094 26844 22098
rect 26712 22092 26844 22094
rect 26712 22066 26792 22092
rect 26792 22034 26844 22040
rect 26792 21888 26844 21894
rect 26792 21830 26844 21836
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26146 18864 26202 18873
rect 26146 18799 26202 18808
rect 26160 18766 26188 18799
rect 26528 18766 26556 19858
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26436 17610 26464 18702
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25884 13326 25912 15438
rect 25976 13394 26004 15846
rect 26054 15192 26110 15201
rect 26054 15127 26110 15136
rect 26068 14006 26096 15127
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12442 25912 13262
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25884 11354 25912 11698
rect 25976 11626 26004 12106
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25780 11280 25832 11286
rect 25780 11222 25832 11228
rect 26160 10674 26188 16934
rect 26252 16658 26280 17478
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26252 16522 26280 16594
rect 26344 16590 26372 17070
rect 26528 16590 26556 18702
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26436 15638 26464 16458
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26252 14550 26280 14962
rect 26240 14544 26292 14550
rect 26240 14486 26292 14492
rect 26620 14414 26648 21490
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26344 12782 26372 13466
rect 26620 13394 26648 14350
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 26528 12918 26556 13194
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 26620 12850 26648 13330
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26252 11558 26280 11698
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 25596 9648 25648 9654
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24308 8900 24360 8906
rect 24308 8842 24360 8848
rect 24320 8430 24348 8842
rect 24872 8650 24900 8910
rect 24780 8622 24900 8650
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24780 7546 24808 8622
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24872 8090 24900 8434
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24320 6390 24348 7142
rect 24964 6866 24992 8910
rect 25056 8498 25084 9454
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8634 25176 8910
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24964 6390 24992 6802
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 22204 4622 22232 5102
rect 23032 4826 23060 5170
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 23584 4554 23612 5306
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23676 4486 23704 6190
rect 24596 5370 24624 6258
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 25056 5166 25084 8434
rect 25148 7886 25176 8570
rect 25240 8022 25268 9590
rect 25332 9574 25452 9602
rect 25596 9590 25648 9596
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25332 9178 25360 9454
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25424 8838 25452 9574
rect 26252 9382 26280 11494
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25228 8016 25280 8022
rect 25228 7958 25280 7964
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25424 6866 25452 8774
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25516 7342 25544 7890
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 25332 6322 25360 6666
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25332 5914 25360 6258
rect 25424 5914 25452 6598
rect 25504 6112 25556 6118
rect 25504 6054 25556 6060
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25516 5778 25544 6054
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25240 5234 25268 5646
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4622 24716 4966
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24964 4486 24992 5102
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 24964 4146 24992 4422
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 25884 4078 25912 7278
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 6338 26096 6734
rect 26252 6730 26280 7482
rect 26344 7002 26372 12718
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26528 10742 26556 11086
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26528 9722 26556 10678
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26712 8974 26740 21082
rect 26804 13326 26832 21830
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26896 10810 26924 20742
rect 26988 19836 27016 23054
rect 27172 22166 27200 24074
rect 27160 22160 27212 22166
rect 27160 22102 27212 22108
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27080 21894 27108 21966
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 27080 21486 27108 21830
rect 27172 21554 27200 22102
rect 27264 22094 27292 24228
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27356 22778 27384 23598
rect 27526 23488 27582 23497
rect 27526 23423 27582 23432
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27264 22066 27384 22094
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 27264 20482 27292 21626
rect 27356 20602 27384 22066
rect 27448 21146 27476 22714
rect 27540 21622 27568 23423
rect 27632 23118 27660 24346
rect 27724 24138 27752 24754
rect 27712 24132 27764 24138
rect 27712 24074 27764 24080
rect 27724 23730 27752 24074
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27632 21962 27660 22578
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27724 22234 27752 22510
rect 27712 22228 27764 22234
rect 27712 22170 27764 22176
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27436 21140 27488 21146
rect 27436 21082 27488 21088
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27264 20466 27384 20482
rect 27264 20460 27396 20466
rect 27264 20454 27344 20460
rect 27068 19848 27120 19854
rect 26988 19808 27068 19836
rect 27068 19790 27120 19796
rect 27080 19446 27108 19790
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 27068 19440 27120 19446
rect 27068 19382 27120 19388
rect 27172 19378 27200 19654
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27264 18698 27292 20454
rect 27344 20402 27396 20408
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27252 18692 27304 18698
rect 27252 18634 27304 18640
rect 27264 17134 27292 18634
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27356 16114 27384 16390
rect 27448 16114 27476 20198
rect 27540 19961 27568 21422
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 20942 27660 21286
rect 27724 21078 27752 22170
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27724 20602 27752 20878
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27632 19990 27660 20402
rect 27620 19984 27672 19990
rect 27526 19952 27582 19961
rect 27620 19926 27672 19932
rect 27526 19887 27582 19896
rect 27724 19242 27752 20538
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 27816 18222 27844 27270
rect 27908 26382 27936 28154
rect 28000 26518 28028 28494
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 27896 26376 27948 26382
rect 27988 26376 28040 26382
rect 27896 26318 27948 26324
rect 27986 26344 27988 26353
rect 28040 26344 28042 26353
rect 27908 25974 27936 26318
rect 27986 26279 28042 26288
rect 27896 25968 27948 25974
rect 27896 25910 27948 25916
rect 28092 25498 28120 34070
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28184 32230 28212 32846
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28172 32224 28224 32230
rect 28172 32166 28224 32172
rect 28184 30734 28212 32166
rect 28276 31890 28304 32302
rect 28356 32224 28408 32230
rect 28356 32166 28408 32172
rect 28264 31884 28316 31890
rect 28264 31826 28316 31832
rect 28276 31482 28304 31826
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28172 30728 28224 30734
rect 28264 30728 28316 30734
rect 28172 30670 28224 30676
rect 28262 30696 28264 30705
rect 28316 30696 28318 30705
rect 28262 30631 28318 30640
rect 28264 29232 28316 29238
rect 28262 29200 28264 29209
rect 28316 29200 28318 29209
rect 28262 29135 28318 29144
rect 28264 29096 28316 29102
rect 28264 29038 28316 29044
rect 28172 29028 28224 29034
rect 28172 28970 28224 28976
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27908 24585 27936 24754
rect 27894 24576 27950 24585
rect 27894 24511 27950 24520
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27908 23594 27936 24142
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 28000 23798 28028 24006
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 28092 23594 28120 25230
rect 28184 24857 28212 28970
rect 28276 28558 28304 29038
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28264 26512 28316 26518
rect 28264 26454 28316 26460
rect 28276 26353 28304 26454
rect 28262 26344 28318 26353
rect 28262 26279 28318 26288
rect 28170 24848 28226 24857
rect 28170 24783 28226 24792
rect 28368 24154 28396 32166
rect 28448 29504 28500 29510
rect 28448 29446 28500 29452
rect 28460 24392 28488 29446
rect 28552 26382 28580 37062
rect 28816 36848 28868 36854
rect 28816 36790 28868 36796
rect 28724 36576 28776 36582
rect 28724 36518 28776 36524
rect 28736 36038 28764 36518
rect 28724 36032 28776 36038
rect 28724 35974 28776 35980
rect 28632 34944 28684 34950
rect 28632 34886 28684 34892
rect 28644 33522 28672 34886
rect 28736 34134 28764 35974
rect 28828 35698 28856 36790
rect 30104 36576 30156 36582
rect 30104 36518 30156 36524
rect 30116 36378 30144 36518
rect 30104 36372 30156 36378
rect 30104 36314 30156 36320
rect 30196 36168 30248 36174
rect 30196 36110 30248 36116
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 28816 35692 28868 35698
rect 28816 35634 28868 35640
rect 29092 35692 29144 35698
rect 29092 35634 29144 35640
rect 29104 35290 29132 35634
rect 29092 35284 29144 35290
rect 29092 35226 29144 35232
rect 29196 35154 29224 35974
rect 30208 35494 30236 36110
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 29184 35148 29236 35154
rect 29184 35090 29236 35096
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 28920 34746 28948 35022
rect 28908 34740 28960 34746
rect 28908 34682 28960 34688
rect 28920 34134 28948 34682
rect 29184 34400 29236 34406
rect 29184 34342 29236 34348
rect 28724 34128 28776 34134
rect 28724 34070 28776 34076
rect 28908 34128 28960 34134
rect 28908 34070 28960 34076
rect 29196 33998 29224 34342
rect 29184 33992 29236 33998
rect 29184 33934 29236 33940
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 28632 33380 28684 33386
rect 28632 33322 28684 33328
rect 28644 32450 28672 33322
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 28736 32570 28764 32846
rect 28816 32836 28868 32842
rect 28816 32778 28868 32784
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28644 32422 28764 32450
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28644 31346 28672 31758
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28632 29232 28684 29238
rect 28632 29174 28684 29180
rect 28644 28422 28672 29174
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28644 28218 28672 28358
rect 28632 28212 28684 28218
rect 28632 28154 28684 28160
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28552 25430 28580 26318
rect 28540 25424 28592 25430
rect 28540 25366 28592 25372
rect 28632 25220 28684 25226
rect 28632 25162 28684 25168
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28552 24562 28580 24686
rect 28644 24682 28672 25162
rect 28632 24676 28684 24682
rect 28632 24618 28684 24624
rect 28552 24534 28672 24562
rect 28460 24364 28580 24392
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28276 24126 28396 24154
rect 27896 23588 27948 23594
rect 27896 23530 27948 23536
rect 28080 23588 28132 23594
rect 28080 23530 28132 23536
rect 27908 22982 27936 23530
rect 27986 23352 28042 23361
rect 27986 23287 28042 23296
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 28000 22710 28028 23287
rect 27988 22704 28040 22710
rect 27988 22646 28040 22652
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27908 20398 27936 21422
rect 28000 21418 28028 21966
rect 28080 21956 28132 21962
rect 28080 21898 28132 21904
rect 27988 21412 28040 21418
rect 27988 21354 28040 21360
rect 27986 21312 28042 21321
rect 27986 21247 28042 21256
rect 28000 20942 28028 21247
rect 28092 20942 28120 21898
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 28184 20534 28212 24074
rect 28276 21321 28304 24126
rect 28552 23526 28580 24364
rect 28644 24206 28672 24534
rect 28736 24274 28764 32422
rect 28828 32230 28856 32778
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 28828 29714 28856 32166
rect 29012 31278 29040 33390
rect 29184 31952 29236 31958
rect 29184 31894 29236 31900
rect 29196 31346 29224 31894
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 29000 31272 29052 31278
rect 29052 31232 29132 31260
rect 29000 31214 29052 31220
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28920 29782 28948 30534
rect 29104 30326 29132 31232
rect 29184 30728 29236 30734
rect 29184 30670 29236 30676
rect 29092 30320 29144 30326
rect 29092 30262 29144 30268
rect 29092 30184 29144 30190
rect 29092 30126 29144 30132
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 29012 29850 29040 29990
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 28816 29708 28868 29714
rect 28816 29650 28868 29656
rect 29104 29170 29132 30126
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29000 29096 29052 29102
rect 29196 29050 29224 30670
rect 29288 29646 29316 35022
rect 30208 34610 30236 35430
rect 30840 35080 30892 35086
rect 30932 35080 30984 35086
rect 30840 35022 30892 35028
rect 30930 35048 30932 35057
rect 30984 35048 30986 35057
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 29472 33590 29500 34546
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29460 33584 29512 33590
rect 29460 33526 29512 33532
rect 29748 32434 29776 33934
rect 29840 33561 29868 33934
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 29826 33552 29882 33561
rect 29826 33487 29882 33496
rect 29918 33144 29974 33153
rect 29918 33079 29974 33088
rect 29932 32910 29960 33079
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 30024 32842 30052 33866
rect 30116 33833 30144 33866
rect 30102 33824 30158 33833
rect 30102 33759 30158 33768
rect 30116 33658 30144 33759
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 30012 32836 30064 32842
rect 30012 32778 30064 32784
rect 30024 32502 30052 32778
rect 30012 32496 30064 32502
rect 30012 32438 30064 32444
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29460 32360 29512 32366
rect 29460 32302 29512 32308
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29380 30394 29408 31690
rect 29368 30388 29420 30394
rect 29368 30330 29420 30336
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 29000 29038 29052 29044
rect 28908 28960 28960 28966
rect 29012 28914 29040 29038
rect 29104 29034 29224 29050
rect 29092 29028 29224 29034
rect 29144 29022 29224 29028
rect 29092 28970 29144 28976
rect 28960 28908 29040 28914
rect 28908 28902 29040 28908
rect 28920 28886 29040 28902
rect 28816 24744 28868 24750
rect 28816 24686 28868 24692
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 28828 24138 28856 24686
rect 28816 24132 28868 24138
rect 28816 24074 28868 24080
rect 28630 24032 28686 24041
rect 28630 23967 28686 23976
rect 28644 23730 28672 23967
rect 28828 23882 28856 24074
rect 28920 24041 28948 28886
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 29012 25974 29040 26930
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 29012 24993 29040 25094
rect 28998 24984 29054 24993
rect 28998 24919 29054 24928
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28906 24032 28962 24041
rect 28906 23967 28962 23976
rect 28828 23854 28948 23882
rect 28632 23724 28684 23730
rect 28632 23666 28684 23672
rect 28920 23662 28948 23854
rect 28908 23656 28960 23662
rect 28908 23598 28960 23604
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28540 23520 28592 23526
rect 28540 23462 28592 23468
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28368 22234 28396 22578
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28460 21622 28488 23462
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28632 23044 28684 23050
rect 28632 22986 28684 22992
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28552 21690 28580 21966
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28448 21344 28500 21350
rect 28262 21312 28318 21321
rect 28448 21286 28500 21292
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28262 21247 28318 21256
rect 28460 21026 28488 21286
rect 28368 20998 28488 21026
rect 28368 20942 28396 20998
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 28078 19952 28134 19961
rect 27908 19689 27936 19926
rect 28078 19887 28134 19896
rect 27988 19780 28040 19786
rect 27988 19722 28040 19728
rect 27894 19680 27950 19689
rect 27894 19615 27950 19624
rect 28000 19378 28028 19722
rect 28092 19446 28120 19887
rect 28184 19854 28212 20470
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28368 19700 28396 20878
rect 28552 20777 28580 21286
rect 28538 20768 28594 20777
rect 28538 20703 28594 20712
rect 28644 20074 28672 22986
rect 28724 22160 28776 22166
rect 28722 22128 28724 22137
rect 28776 22128 28778 22137
rect 28722 22063 28778 22072
rect 28724 22024 28776 22030
rect 28828 22012 28856 23054
rect 28776 21984 28856 22012
rect 28724 21966 28776 21972
rect 28736 20466 28764 21966
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28184 19672 28396 19700
rect 28460 20058 28672 20074
rect 28460 20052 28684 20058
rect 28460 20046 28632 20052
rect 28080 19440 28132 19446
rect 28080 19382 28132 19388
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27988 18624 28040 18630
rect 27988 18566 28040 18572
rect 27908 18358 27936 18566
rect 27896 18352 27948 18358
rect 27896 18294 27948 18300
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 17678 27660 18022
rect 27816 17678 27844 18158
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 27540 16658 27568 16730
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27632 16182 27660 16526
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27172 15706 27200 16050
rect 27160 15700 27212 15706
rect 27160 15642 27212 15648
rect 27540 15502 27568 16050
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14618 27384 14962
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27172 13938 27200 14350
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27448 13870 27476 15098
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27540 14618 27568 14894
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27264 12986 27292 13262
rect 27448 13258 27476 13806
rect 27436 13252 27488 13258
rect 27436 13194 27488 13200
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27448 12238 27476 13194
rect 27618 12336 27674 12345
rect 27618 12271 27674 12280
rect 27632 12238 27660 12271
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27528 12096 27580 12102
rect 27526 12064 27528 12073
rect 27580 12064 27582 12073
rect 27526 11999 27582 12008
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27632 11218 27660 11290
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27172 10810 27200 11018
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27632 10742 27660 11154
rect 27724 11150 27752 17614
rect 28000 17202 28028 18566
rect 28080 17264 28132 17270
rect 28080 17206 28132 17212
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 28092 16522 28120 17206
rect 28184 16590 28212 19672
rect 28460 19553 28488 20046
rect 28632 19994 28684 20000
rect 28630 19952 28686 19961
rect 28630 19887 28686 19896
rect 28644 19836 28672 19887
rect 28724 19848 28776 19854
rect 28644 19808 28724 19836
rect 28724 19790 28776 19796
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28722 19680 28778 19689
rect 28446 19544 28502 19553
rect 28446 19479 28502 19488
rect 28552 19310 28580 19654
rect 28644 19417 28672 19654
rect 28722 19615 28778 19624
rect 28630 19408 28686 19417
rect 28630 19343 28686 19352
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28276 18426 28304 18634
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 28368 18222 28396 19246
rect 28538 19136 28594 19145
rect 28538 19071 28594 19080
rect 28552 18766 28580 19071
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28448 18148 28500 18154
rect 28448 18090 28500 18096
rect 28460 17202 28488 18090
rect 28644 17270 28672 19343
rect 28736 18698 28764 19615
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28828 17490 28856 21626
rect 28920 19854 28948 23462
rect 29012 23186 29040 24754
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 29104 22982 29132 28970
rect 29472 25906 29500 32302
rect 29748 30938 29776 32370
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 29748 30258 29776 30874
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29748 29646 29776 30194
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29644 29572 29696 29578
rect 29644 29514 29696 29520
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29564 26586 29592 27950
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29564 26314 29592 26522
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29460 25900 29512 25906
rect 29460 25842 29512 25848
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29368 24336 29420 24342
rect 29368 24278 29420 24284
rect 29276 24064 29328 24070
rect 29276 24006 29328 24012
rect 29288 23730 29316 24006
rect 29380 23730 29408 24278
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29368 23520 29420 23526
rect 29368 23462 29420 23468
rect 29184 23180 29236 23186
rect 29184 23122 29236 23128
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 29104 22030 29132 22918
rect 29196 22030 29224 23122
rect 29276 22160 29328 22166
rect 29276 22102 29328 22108
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 29184 22024 29236 22030
rect 29184 21966 29236 21972
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 29012 20466 29040 20538
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29104 20369 29132 21966
rect 29090 20360 29146 20369
rect 29090 20295 29146 20304
rect 29288 20097 29316 22102
rect 29380 21894 29408 23462
rect 29368 21888 29420 21894
rect 29368 21830 29420 21836
rect 29368 21412 29420 21418
rect 29368 21354 29420 21360
rect 29380 21010 29408 21354
rect 29368 21004 29420 21010
rect 29368 20946 29420 20952
rect 29472 20942 29500 24754
rect 29552 24676 29604 24682
rect 29552 24618 29604 24624
rect 29564 24206 29592 24618
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29552 23656 29604 23662
rect 29552 23598 29604 23604
rect 29564 23186 29592 23598
rect 29552 23180 29604 23186
rect 29552 23122 29604 23128
rect 29656 21978 29684 29514
rect 29748 28082 29776 29582
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29748 27674 29776 28018
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29734 27568 29790 27577
rect 29734 27503 29790 27512
rect 29748 26994 29776 27503
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29736 24132 29788 24138
rect 29736 24074 29788 24080
rect 29748 23730 29776 24074
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 29748 23118 29776 23666
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29564 21950 29684 21978
rect 29564 21570 29592 21950
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29656 21690 29684 21830
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29564 21542 29684 21570
rect 29656 21146 29684 21542
rect 29644 21140 29696 21146
rect 29644 21082 29696 21088
rect 29642 21040 29698 21049
rect 29552 21004 29604 21010
rect 29642 20975 29698 20984
rect 29552 20946 29604 20952
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29274 20088 29330 20097
rect 29274 20023 29330 20032
rect 29090 19952 29146 19961
rect 29090 19887 29092 19896
rect 29144 19887 29146 19896
rect 29092 19858 29144 19864
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 29012 19689 29040 19790
rect 29184 19712 29236 19718
rect 28998 19680 29054 19689
rect 28998 19615 29054 19624
rect 29182 19680 29184 19689
rect 29236 19680 29238 19689
rect 29182 19615 29238 19624
rect 28906 19544 28962 19553
rect 29090 19544 29146 19553
rect 28906 19479 28962 19488
rect 29012 19502 29090 19530
rect 28920 18408 28948 19479
rect 29012 18630 29040 19502
rect 29090 19479 29146 19488
rect 29092 19440 29144 19446
rect 29090 19408 29092 19417
rect 29144 19408 29146 19417
rect 29274 19408 29330 19417
rect 29090 19343 29146 19352
rect 29196 19366 29274 19394
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 28920 18380 29040 18408
rect 28908 18284 28960 18290
rect 28908 18226 28960 18232
rect 28920 17610 28948 18226
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 28828 17462 28948 17490
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28448 17196 28500 17202
rect 28500 17156 28580 17184
rect 28448 17138 28500 17144
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28276 16590 28304 17070
rect 28448 17060 28500 17066
rect 28448 17002 28500 17008
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28460 16522 28488 17002
rect 28080 16516 28132 16522
rect 28080 16458 28132 16464
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 27986 15192 28042 15201
rect 27986 15127 28042 15136
rect 28000 14006 28028 15127
rect 27988 14000 28040 14006
rect 27988 13942 28040 13948
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27908 12850 27936 13874
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 28000 13394 28028 13670
rect 27988 13388 28040 13394
rect 27988 13330 28040 13336
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27816 12442 27844 12718
rect 27804 12436 27856 12442
rect 27804 12378 27856 12384
rect 27896 11280 27948 11286
rect 27896 11222 27948 11228
rect 27712 11144 27764 11150
rect 27712 11086 27764 11092
rect 27724 10742 27752 11086
rect 27908 10810 27936 11222
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27712 10736 27764 10742
rect 27712 10678 27764 10684
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26436 7886 26464 8842
rect 26896 8838 26924 9318
rect 27264 9042 27292 9522
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 27448 8634 27476 9522
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27632 8498 27660 10678
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27816 10130 27844 10542
rect 27804 10124 27856 10130
rect 27804 10066 27856 10072
rect 27816 9722 27844 10066
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27632 8378 27660 8434
rect 27448 8350 27660 8378
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26332 6996 26384 7002
rect 26332 6938 26384 6944
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 26240 6724 26292 6730
rect 26240 6666 26292 6672
rect 26160 6458 26188 6666
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26068 6322 26188 6338
rect 26252 6322 26280 6666
rect 26436 6322 26464 7822
rect 27160 7812 27212 7818
rect 27160 7754 27212 7760
rect 27172 7546 27200 7754
rect 27160 7540 27212 7546
rect 27160 7482 27212 7488
rect 27448 7478 27476 8350
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27540 7546 27568 7686
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27816 7342 27844 8230
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 26068 6316 26200 6322
rect 26068 6310 26148 6316
rect 26148 6258 26200 6264
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25976 4758 26004 5170
rect 26068 4758 26096 6190
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 26068 4282 26096 4694
rect 27264 4622 27292 6258
rect 27908 5914 27936 6258
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26528 4282 26556 4490
rect 26056 4276 26108 4282
rect 26056 4218 26108 4224
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 27264 4146 27292 4558
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 28092 2446 28120 15846
rect 28460 15434 28488 16458
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 28446 15192 28502 15201
rect 28446 15127 28502 15136
rect 28354 15056 28410 15065
rect 28354 14991 28356 15000
rect 28408 14991 28410 15000
rect 28356 14962 28408 14968
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28184 5778 28212 14758
rect 28460 14006 28488 15127
rect 28552 14006 28580 17156
rect 28920 16114 28948 17462
rect 29012 17202 29040 18380
rect 29104 18222 29132 19246
rect 29196 19174 29224 19366
rect 29274 19343 29330 19352
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29276 19168 29328 19174
rect 29276 19110 29328 19116
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 29012 16114 29040 16390
rect 29104 16114 29132 18158
rect 29196 16590 29224 19110
rect 29288 18154 29316 19110
rect 29276 18148 29328 18154
rect 29276 18090 29328 18096
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 28828 15706 28856 16050
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 29104 15502 29132 16050
rect 29182 15600 29238 15609
rect 29182 15535 29238 15544
rect 29196 15502 29224 15535
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29184 15496 29236 15502
rect 29184 15438 29236 15444
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 29012 14278 29040 14894
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 29104 14006 29132 14214
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28540 14000 28592 14006
rect 29092 14000 29144 14006
rect 28540 13942 28592 13948
rect 28998 13968 29054 13977
rect 28552 13870 28580 13942
rect 29092 13942 29144 13948
rect 28998 13903 29000 13912
rect 29052 13903 29054 13912
rect 29000 13874 29052 13880
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 28908 13796 28960 13802
rect 28908 13738 28960 13744
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28460 10742 28488 10950
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28264 8424 28316 8430
rect 28264 8366 28316 8372
rect 28276 7886 28304 8366
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28276 6866 28304 7822
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 28184 5234 28212 5714
rect 28276 5710 28304 6394
rect 28460 6118 28488 9658
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28552 8634 28580 9318
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28828 6866 28856 8774
rect 28920 7546 28948 13738
rect 29104 13326 29132 13942
rect 29196 13530 29224 15438
rect 29288 14618 29316 16594
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29104 11694 29132 12378
rect 29092 11688 29144 11694
rect 29092 11630 29144 11636
rect 29104 11218 29132 11630
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29012 8090 29040 9522
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 29104 7954 29132 11154
rect 29288 11098 29316 14554
rect 29380 12850 29408 20742
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29472 19378 29500 19654
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29472 17746 29500 19314
rect 29564 18426 29592 20946
rect 29656 19378 29684 20975
rect 29748 20398 29776 23054
rect 29840 21690 29868 30670
rect 30024 30326 30052 32438
rect 30012 30320 30064 30326
rect 30012 30262 30064 30268
rect 30024 29646 30052 30262
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 30116 30161 30144 30194
rect 30102 30152 30158 30161
rect 30102 30087 30104 30096
rect 30156 30087 30158 30096
rect 30104 30058 30156 30064
rect 29920 29640 29972 29646
rect 29920 29582 29972 29588
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 29932 28558 29960 29582
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29932 28422 29960 28494
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 30024 28150 30052 29582
rect 30104 29572 30156 29578
rect 30104 29514 30156 29520
rect 30116 29306 30144 29514
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 30116 29073 30144 29242
rect 30102 29064 30158 29073
rect 30102 28999 30158 29008
rect 30012 28144 30064 28150
rect 30012 28086 30064 28092
rect 29920 27464 29972 27470
rect 30024 27452 30052 28086
rect 30104 27464 30156 27470
rect 30024 27424 30104 27452
rect 29920 27406 29972 27412
rect 30104 27406 30156 27412
rect 29932 26518 29960 27406
rect 30116 26994 30144 27406
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 29920 26512 29972 26518
rect 29920 26454 29972 26460
rect 30208 26450 30236 34546
rect 30288 33992 30340 33998
rect 30288 33934 30340 33940
rect 30300 33538 30328 33934
rect 30300 33510 30420 33538
rect 30288 33448 30340 33454
rect 30288 33390 30340 33396
rect 30300 33046 30328 33390
rect 30288 33040 30340 33046
rect 30288 32982 30340 32988
rect 30288 32904 30340 32910
rect 30392 32858 30420 33510
rect 30668 33114 30696 34546
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30340 32852 30420 32858
rect 30288 32846 30420 32852
rect 30300 32830 30420 32846
rect 30300 32450 30328 32830
rect 30300 32422 30420 32450
rect 30392 32366 30420 32422
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30288 32360 30340 32366
rect 30288 32302 30340 32308
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30300 32026 30328 32302
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30392 31906 30420 32302
rect 30300 31890 30420 31906
rect 30288 31884 30420 31890
rect 30340 31878 30420 31884
rect 30288 31826 30340 31832
rect 30300 30258 30328 31826
rect 30484 31657 30512 32370
rect 30760 31754 30788 34546
rect 30852 34202 30880 35022
rect 30930 34983 30986 34992
rect 30932 34944 30984 34950
rect 30932 34886 30984 34892
rect 30944 34610 30972 34886
rect 31036 34610 31064 37130
rect 31864 36718 31892 37130
rect 32772 36848 32824 36854
rect 32772 36790 32824 36796
rect 32404 36780 32456 36786
rect 32404 36722 32456 36728
rect 31852 36712 31904 36718
rect 31852 36654 31904 36660
rect 31484 36236 31536 36242
rect 31484 36178 31536 36184
rect 31208 35216 31260 35222
rect 31208 35158 31260 35164
rect 31220 35018 31248 35158
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 31496 34746 31524 36178
rect 31864 36106 31892 36654
rect 32416 36378 32444 36722
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32680 36168 32732 36174
rect 32680 36110 32732 36116
rect 31852 36100 31904 36106
rect 31852 36042 31904 36048
rect 32496 36100 32548 36106
rect 32496 36042 32548 36048
rect 32508 35698 32536 36042
rect 32692 35698 32720 36110
rect 32496 35692 32548 35698
rect 32496 35634 32548 35640
rect 32680 35692 32732 35698
rect 32680 35634 32732 35640
rect 32508 35290 32536 35634
rect 32496 35284 32548 35290
rect 32496 35226 32548 35232
rect 31576 35080 31628 35086
rect 31576 35022 31628 35028
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 31588 34610 31616 35022
rect 32496 35012 32548 35018
rect 32496 34954 32548 34960
rect 32508 34678 32536 34954
rect 32692 34746 32720 35634
rect 32680 34740 32732 34746
rect 32680 34682 32732 34688
rect 32496 34672 32548 34678
rect 32496 34614 32548 34620
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 31024 34604 31076 34610
rect 31024 34546 31076 34552
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 30840 34196 30892 34202
rect 30840 34138 30892 34144
rect 30944 33930 30972 34546
rect 31392 34468 31444 34474
rect 31392 34410 31444 34416
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 30932 33924 30984 33930
rect 30932 33866 30984 33872
rect 30944 33590 30972 33866
rect 30932 33584 30984 33590
rect 30932 33526 30984 33532
rect 30760 31726 30880 31754
rect 30470 31648 30526 31657
rect 30470 31583 30526 31592
rect 30484 30841 30512 31583
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30470 30832 30526 30841
rect 30470 30767 30526 30776
rect 30472 30660 30524 30666
rect 30472 30602 30524 30608
rect 30484 30326 30512 30602
rect 30668 30394 30696 31282
rect 30760 31249 30788 31282
rect 30746 31240 30802 31249
rect 30746 31175 30802 31184
rect 30748 30728 30800 30734
rect 30748 30670 30800 30676
rect 30656 30388 30708 30394
rect 30656 30330 30708 30336
rect 30472 30320 30524 30326
rect 30472 30262 30524 30268
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30300 29646 30328 30194
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30300 28082 30328 29582
rect 30392 28218 30420 29582
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 30288 28076 30340 28082
rect 30288 28018 30340 28024
rect 30300 27606 30328 28018
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30288 27600 30340 27606
rect 30288 27542 30340 27548
rect 30288 27328 30340 27334
rect 30288 27270 30340 27276
rect 30196 26444 30248 26450
rect 30116 26404 30196 26432
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 29932 24818 29960 26318
rect 30116 25226 30144 26404
rect 30196 26386 30248 26392
rect 30196 26240 30248 26246
rect 30196 26182 30248 26188
rect 30208 25906 30236 26182
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 30300 25838 30328 27270
rect 30392 26353 30420 27950
rect 30378 26344 30434 26353
rect 30378 26279 30434 26288
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30104 25220 30156 25226
rect 30104 25162 30156 25168
rect 30288 25220 30340 25226
rect 30392 25208 30420 26279
rect 30340 25180 30420 25208
rect 30288 25162 30340 25168
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 29920 24676 29972 24682
rect 29920 24618 29972 24624
rect 29932 24206 29960 24618
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 29932 23866 29960 24142
rect 30024 24138 30052 24550
rect 30012 24132 30064 24138
rect 30012 24074 30064 24080
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 30104 23248 30156 23254
rect 30104 23190 30156 23196
rect 30010 22808 30066 22817
rect 30010 22743 30066 22752
rect 30024 22710 30052 22743
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 29920 22160 29972 22166
rect 29920 22102 29972 22108
rect 29932 21690 29960 22102
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 30024 21570 30052 22646
rect 30116 21944 30144 23190
rect 30300 23050 30328 25162
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30392 24410 30420 24754
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 30484 22098 30512 30262
rect 30760 29850 30788 30670
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30748 29708 30800 29714
rect 30748 29650 30800 29656
rect 30656 29164 30708 29170
rect 30656 29106 30708 29112
rect 30668 27538 30696 29106
rect 30656 27532 30708 27538
rect 30576 27492 30656 27520
rect 30576 25362 30604 27492
rect 30656 27474 30708 27480
rect 30760 25906 30788 29650
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30748 25900 30800 25906
rect 30748 25842 30800 25848
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30668 23798 30696 25842
rect 30746 25800 30802 25809
rect 30746 25735 30802 25744
rect 30760 25702 30788 25735
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30656 23792 30708 23798
rect 30656 23734 30708 23740
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30576 23118 30604 23666
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 22092 30524 22098
rect 30472 22034 30524 22040
rect 30380 22024 30432 22030
rect 30378 21992 30380 22001
rect 30432 21992 30434 22001
rect 30196 21956 30248 21962
rect 30116 21916 30196 21944
rect 30378 21927 30434 21936
rect 30196 21898 30248 21904
rect 29828 21548 29880 21554
rect 29828 21490 29880 21496
rect 29932 21542 30052 21570
rect 30104 21616 30156 21622
rect 30104 21558 30156 21564
rect 29840 20806 29868 21490
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29734 20088 29790 20097
rect 29840 20058 29868 20198
rect 29734 20023 29790 20032
rect 29828 20052 29880 20058
rect 29748 19854 29776 20023
rect 29828 19994 29880 20000
rect 29932 19854 29960 21542
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 30024 21185 30052 21422
rect 30010 21176 30066 21185
rect 30010 21111 30066 21120
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29748 18698 29776 19314
rect 29840 19242 29868 19790
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 30010 19680 30066 19689
rect 29828 19236 29880 19242
rect 29828 19178 29880 19184
rect 29736 18692 29788 18698
rect 29736 18634 29788 18640
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29828 17264 29880 17270
rect 29828 17206 29880 17212
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 13938 29500 16934
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29380 11218 29408 12786
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29288 11070 29408 11098
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 29104 6914 29132 7890
rect 29104 6886 29224 6914
rect 28816 6860 28868 6866
rect 28816 6802 28868 6808
rect 28828 6662 28856 6802
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28632 6316 28684 6322
rect 28632 6258 28684 6264
rect 28448 6112 28500 6118
rect 28448 6054 28500 6060
rect 28460 5778 28488 6054
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28184 4690 28212 5170
rect 28172 4684 28224 4690
rect 28172 4626 28224 4632
rect 28644 4622 28672 6258
rect 29196 4690 29224 6886
rect 29288 6798 29316 9522
rect 29380 9330 29408 11070
rect 29564 9500 29592 15846
rect 29656 14958 29684 17138
rect 29840 16658 29868 17206
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29644 14000 29696 14006
rect 29748 13977 29776 16526
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29644 13942 29696 13948
rect 29734 13968 29790 13977
rect 29656 13462 29684 13942
rect 29734 13903 29790 13912
rect 29736 13864 29788 13870
rect 29734 13832 29736 13841
rect 29788 13832 29790 13841
rect 29734 13767 29790 13776
rect 29644 13456 29696 13462
rect 29644 13398 29696 13404
rect 29840 13394 29868 14282
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29932 12434 29960 19654
rect 30010 19615 30066 19624
rect 30024 16590 30052 19615
rect 30116 19417 30144 21558
rect 30208 21486 30236 21898
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 30208 19446 30236 21422
rect 30196 19440 30248 19446
rect 30102 19408 30158 19417
rect 30196 19382 30248 19388
rect 30102 19343 30158 19352
rect 30104 19236 30156 19242
rect 30104 19178 30156 19184
rect 30116 18834 30144 19178
rect 30104 18828 30156 18834
rect 30104 18770 30156 18776
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 30102 13968 30158 13977
rect 30102 13903 30104 13912
rect 30156 13903 30158 13912
rect 30104 13874 30156 13880
rect 30012 13728 30064 13734
rect 30012 13670 30064 13676
rect 29840 12406 29960 12434
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29656 9654 29684 11086
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29564 9472 29684 9500
rect 29380 9302 29592 9330
rect 29368 8900 29420 8906
rect 29368 8842 29420 8848
rect 29380 8498 29408 8842
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29472 6866 29500 8298
rect 29564 6866 29592 9302
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29288 6254 29316 6734
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29472 6186 29500 6802
rect 29460 6180 29512 6186
rect 29460 6122 29512 6128
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28276 4214 28304 4422
rect 28644 4282 28672 4558
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28264 4208 28316 4214
rect 28264 4150 28316 4156
rect 29656 3942 29684 9472
rect 29840 8634 29868 12406
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29932 10810 29960 11018
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 29920 6724 29972 6730
rect 29920 6666 29972 6672
rect 29932 6458 29960 6666
rect 29920 6452 29972 6458
rect 29920 6394 29972 6400
rect 30024 6118 30052 13670
rect 30208 12434 30236 18022
rect 30392 17270 30420 21927
rect 30576 21622 30604 22918
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 30668 21010 30696 23734
rect 30760 22094 30788 25638
rect 30852 24070 30880 31726
rect 30944 31414 30972 33526
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 31036 32570 31064 33458
rect 31220 33114 31248 33934
rect 31404 33522 31432 34410
rect 31588 33946 31616 34546
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 31668 33992 31720 33998
rect 31588 33940 31668 33946
rect 31588 33934 31720 33940
rect 31588 33918 31708 33934
rect 31760 33924 31812 33930
rect 31588 33522 31616 33918
rect 31760 33866 31812 33872
rect 31666 33824 31722 33833
rect 31772 33810 31800 33866
rect 31722 33782 31800 33810
rect 32128 33856 32180 33862
rect 32128 33798 32180 33804
rect 31666 33759 31722 33768
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31576 33516 31628 33522
rect 31576 33458 31628 33464
rect 31208 33108 31260 33114
rect 31208 33050 31260 33056
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 31312 32910 31340 33050
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31116 32836 31168 32842
rect 31116 32778 31168 32784
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 31128 32502 31156 32778
rect 31116 32496 31168 32502
rect 31116 32438 31168 32444
rect 31312 32298 31340 32846
rect 31300 32292 31352 32298
rect 31300 32234 31352 32240
rect 31404 31754 31432 33458
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 31496 32434 31524 32846
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31312 31726 31432 31754
rect 31116 31680 31168 31686
rect 31116 31622 31168 31628
rect 30932 31408 30984 31414
rect 30932 31350 30984 31356
rect 30944 30734 30972 31350
rect 31128 31346 31156 31622
rect 31208 31408 31260 31414
rect 31208 31350 31260 31356
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31128 30802 31156 31282
rect 31116 30796 31168 30802
rect 31116 30738 31168 30744
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31024 30048 31076 30054
rect 31024 29990 31076 29996
rect 31036 29850 31064 29990
rect 31024 29844 31076 29850
rect 31024 29786 31076 29792
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30944 29073 30972 29106
rect 30930 29064 30986 29073
rect 30930 28999 30986 29008
rect 30932 27668 30984 27674
rect 30932 27610 30984 27616
rect 30944 27402 30972 27610
rect 30932 27396 30984 27402
rect 30932 27338 30984 27344
rect 31036 25906 31064 29786
rect 31128 28966 31156 30602
rect 31220 29209 31248 31350
rect 31312 31210 31340 31726
rect 31588 31686 31616 33458
rect 31944 33040 31996 33046
rect 31944 32982 31996 32988
rect 31668 32836 31720 32842
rect 31668 32778 31720 32784
rect 31680 32570 31708 32778
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31668 32564 31720 32570
rect 31668 32506 31720 32512
rect 31576 31680 31628 31686
rect 31576 31622 31628 31628
rect 31300 31204 31352 31210
rect 31300 31146 31352 31152
rect 31312 31113 31340 31146
rect 31298 31104 31354 31113
rect 31298 31039 31354 31048
rect 31484 30728 31536 30734
rect 31484 30670 31536 30676
rect 31300 30592 31352 30598
rect 31300 30534 31352 30540
rect 31312 29578 31340 30534
rect 31496 29646 31524 30670
rect 31680 29850 31708 32506
rect 31668 29844 31720 29850
rect 31668 29786 31720 29792
rect 31484 29640 31536 29646
rect 31404 29600 31484 29628
rect 31300 29572 31352 29578
rect 31300 29514 31352 29520
rect 31206 29200 31262 29209
rect 31206 29135 31262 29144
rect 31116 28960 31168 28966
rect 31116 28902 31168 28908
rect 31128 28626 31156 28902
rect 31312 28762 31340 29514
rect 31404 29170 31432 29600
rect 31484 29582 31536 29588
rect 31484 29504 31536 29510
rect 31482 29472 31484 29481
rect 31536 29472 31538 29481
rect 31482 29407 31538 29416
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31484 29164 31536 29170
rect 31484 29106 31536 29112
rect 31404 28762 31432 29106
rect 31300 28756 31352 28762
rect 31300 28698 31352 28704
rect 31392 28756 31444 28762
rect 31392 28698 31444 28704
rect 31116 28620 31168 28626
rect 31116 28562 31168 28568
rect 31208 28552 31260 28558
rect 31208 28494 31260 28500
rect 31220 27674 31248 28494
rect 31392 28484 31444 28490
rect 31392 28426 31444 28432
rect 31116 27668 31168 27674
rect 31116 27610 31168 27616
rect 31208 27668 31260 27674
rect 31208 27610 31260 27616
rect 31128 27130 31156 27610
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 31024 25900 31076 25906
rect 30944 25860 31024 25888
rect 30944 24886 30972 25860
rect 31024 25842 31076 25848
rect 31024 25356 31076 25362
rect 31024 25298 31076 25304
rect 30932 24880 30984 24886
rect 30932 24822 30984 24828
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 31036 23730 31064 25298
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31036 22642 31064 23666
rect 31128 23662 31156 27066
rect 31404 26926 31432 28426
rect 31496 26994 31524 29106
rect 31772 28994 31800 32710
rect 31852 32360 31904 32366
rect 31852 32302 31904 32308
rect 31588 28966 31800 28994
rect 31484 26988 31536 26994
rect 31484 26930 31536 26936
rect 31392 26920 31444 26926
rect 31392 26862 31444 26868
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 31208 24200 31260 24206
rect 31206 24168 31208 24177
rect 31260 24168 31262 24177
rect 31206 24103 31262 24112
rect 31312 24070 31340 24686
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31128 22710 31156 23598
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 31116 22568 31168 22574
rect 31116 22510 31168 22516
rect 30760 22066 31064 22094
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30944 21418 30972 21966
rect 30932 21412 30984 21418
rect 30932 21354 30984 21360
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30760 20913 30788 21286
rect 30840 21004 30892 21010
rect 30840 20946 30892 20952
rect 30746 20904 30802 20913
rect 30746 20839 30802 20848
rect 30760 20466 30788 20839
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30668 20233 30696 20402
rect 30748 20256 30800 20262
rect 30654 20224 30710 20233
rect 30748 20198 30800 20204
rect 30654 20159 30710 20168
rect 30668 19922 30696 20159
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30380 17264 30432 17270
rect 30380 17206 30432 17212
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30286 16688 30342 16697
rect 30392 16658 30420 17070
rect 30484 16794 30512 17614
rect 30760 17610 30788 20198
rect 30852 18766 30880 20946
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30944 19514 30972 20402
rect 31036 19825 31064 22066
rect 31022 19816 31078 19825
rect 31022 19751 31024 19760
rect 31076 19751 31078 19760
rect 31024 19722 31076 19728
rect 30932 19508 30984 19514
rect 30932 19450 30984 19456
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30748 17604 30800 17610
rect 30748 17546 30800 17552
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30472 16788 30524 16794
rect 30472 16730 30524 16736
rect 30286 16623 30288 16632
rect 30340 16623 30342 16632
rect 30380 16652 30432 16658
rect 30288 16594 30340 16600
rect 30380 16594 30432 16600
rect 30378 16416 30434 16425
rect 30378 16351 30434 16360
rect 30392 16114 30420 16351
rect 30484 16182 30512 16730
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30392 15570 30420 16050
rect 30380 15564 30432 15570
rect 30380 15506 30432 15512
rect 30668 15473 30696 17206
rect 30760 16522 30788 17546
rect 30852 17202 30880 18702
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30944 17338 30972 17478
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30840 17196 30892 17202
rect 30840 17138 30892 17144
rect 31036 16590 31064 18770
rect 31128 17746 31156 22510
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31220 21622 31248 21966
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 31128 17270 31156 17682
rect 31116 17264 31168 17270
rect 31116 17206 31168 17212
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 30748 16516 30800 16522
rect 30748 16458 30800 16464
rect 30944 16289 30972 16526
rect 30930 16280 30986 16289
rect 31128 16250 31156 17206
rect 30930 16215 30986 16224
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31220 16130 31248 21558
rect 31312 21146 31340 24006
rect 31404 23338 31432 26862
rect 31484 24268 31536 24274
rect 31588 24256 31616 28966
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31680 27606 31708 28494
rect 31772 28218 31800 28494
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31864 28150 31892 32302
rect 31852 28144 31904 28150
rect 31852 28086 31904 28092
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31956 26738 31984 32982
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 32048 31142 32076 31758
rect 32036 31136 32088 31142
rect 32036 31078 32088 31084
rect 32048 30870 32076 31078
rect 32036 30864 32088 30870
rect 32036 30806 32088 30812
rect 32036 28484 32088 28490
rect 32036 28426 32088 28432
rect 32048 27334 32076 28426
rect 32036 27328 32088 27334
rect 32036 27270 32088 27276
rect 31864 26710 31984 26738
rect 31668 25832 31720 25838
rect 31668 25774 31720 25780
rect 31536 24228 31616 24256
rect 31484 24210 31536 24216
rect 31496 23526 31524 24210
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31484 23520 31536 23526
rect 31484 23462 31536 23468
rect 31588 23338 31616 23666
rect 31404 23310 31616 23338
rect 31588 22642 31616 23310
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31484 22024 31536 22030
rect 31484 21966 31536 21972
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31404 21078 31432 21830
rect 31496 21554 31524 21966
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31392 21072 31444 21078
rect 31444 21020 31616 21026
rect 31392 21014 31616 21020
rect 31404 21010 31616 21014
rect 31404 21004 31628 21010
rect 31404 20998 31576 21004
rect 31404 20482 31432 20998
rect 31576 20946 31628 20952
rect 31484 20868 31536 20874
rect 31484 20810 31536 20816
rect 31312 20454 31432 20482
rect 31312 18766 31340 20454
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 31312 16590 31340 18702
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 30944 16114 31248 16130
rect 30932 16108 31248 16114
rect 30984 16102 31248 16108
rect 30932 16050 30984 16056
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 30852 15638 30880 15982
rect 30840 15632 30892 15638
rect 30840 15574 30892 15580
rect 30654 15464 30710 15473
rect 30654 15399 30710 15408
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30208 12406 30328 12434
rect 30196 9580 30248 9586
rect 30196 9522 30248 9528
rect 30208 8974 30236 9522
rect 30300 9518 30328 12406
rect 30392 11762 30420 14894
rect 30668 14414 30696 15399
rect 30944 15026 30972 16050
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31036 15094 31064 15302
rect 31312 15094 31340 16526
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 31300 15088 31352 15094
rect 31300 15030 31352 15036
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 31300 14544 31352 14550
rect 31114 14512 31170 14521
rect 31300 14486 31352 14492
rect 31114 14447 31170 14456
rect 30656 14408 30708 14414
rect 30656 14350 30708 14356
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30944 13326 30972 14010
rect 31128 13938 31156 14447
rect 31312 13938 31340 14486
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31300 13932 31352 13938
rect 31300 13874 31352 13880
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 31036 13530 31064 13806
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31404 12374 31432 20266
rect 31496 19281 31524 20810
rect 31680 20618 31708 25774
rect 31864 25294 31892 26710
rect 32048 25770 32076 27270
rect 32036 25764 32088 25770
rect 32036 25706 32088 25712
rect 31852 25288 31904 25294
rect 31852 25230 31904 25236
rect 32036 25288 32088 25294
rect 32036 25230 32088 25236
rect 31864 24426 31892 25230
rect 31944 25152 31996 25158
rect 31944 25094 31996 25100
rect 31772 24398 31892 24426
rect 31772 23730 31800 24398
rect 31852 24336 31904 24342
rect 31852 24278 31904 24284
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31772 22506 31800 23666
rect 31760 22500 31812 22506
rect 31760 22442 31812 22448
rect 31864 22234 31892 24278
rect 31852 22228 31904 22234
rect 31852 22170 31904 22176
rect 31852 21072 31904 21078
rect 31852 21014 31904 21020
rect 31588 20590 31708 20618
rect 31588 20262 31616 20590
rect 31668 20528 31720 20534
rect 31668 20470 31720 20476
rect 31576 20256 31628 20262
rect 31576 20198 31628 20204
rect 31576 19984 31628 19990
rect 31576 19926 31628 19932
rect 31482 19272 31538 19281
rect 31482 19207 31538 19216
rect 31496 18834 31524 19207
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31484 15904 31536 15910
rect 31484 15846 31536 15852
rect 31496 15570 31524 15846
rect 31484 15564 31536 15570
rect 31484 15506 31536 15512
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31484 12300 31536 12306
rect 31484 12242 31536 12248
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30576 11762 30604 12038
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 31208 9376 31260 9382
rect 31208 9318 31260 9324
rect 30576 9110 30604 9318
rect 30656 9172 30708 9178
rect 30656 9114 30708 9120
rect 30564 9104 30616 9110
rect 30564 9046 30616 9052
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30208 8566 30236 8910
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 30208 7886 30236 8502
rect 30484 8498 30512 8910
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30576 6866 30604 9046
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30392 6458 30420 6734
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 30576 5914 30604 6802
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29748 4690 29776 5646
rect 30472 5636 30524 5642
rect 30472 5578 30524 5584
rect 30484 5370 30512 5578
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 29736 4684 29788 4690
rect 29736 4626 29788 4632
rect 30104 4548 30156 4554
rect 30104 4490 30156 4496
rect 30116 4282 30144 4490
rect 30104 4276 30156 4282
rect 30104 4218 30156 4224
rect 30576 4214 30604 5170
rect 30668 5166 30696 9114
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30760 8498 30788 8842
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30944 7886 30972 8910
rect 31220 8906 31248 9318
rect 31208 8900 31260 8906
rect 31208 8842 31260 8848
rect 31312 8566 31340 11018
rect 31496 11014 31524 12242
rect 31588 12238 31616 19926
rect 31680 19446 31708 20470
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 31864 19310 31892 21014
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 31864 18766 31892 19246
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 31668 18080 31720 18086
rect 31668 18022 31720 18028
rect 31680 14618 31708 18022
rect 31864 17762 31892 18702
rect 31772 17734 31892 17762
rect 31772 16046 31800 17734
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 31864 17202 31892 17614
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31956 16590 31984 25094
rect 32048 24886 32076 25230
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 32048 24274 32076 24822
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 32048 21486 32076 24006
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 32048 16980 32076 19722
rect 32140 17134 32168 33798
rect 32232 32910 32260 34478
rect 32404 34400 32456 34406
rect 32404 34342 32456 34348
rect 32416 33658 32444 34342
rect 32508 34202 32536 34614
rect 32496 34196 32548 34202
rect 32496 34138 32548 34144
rect 32680 33856 32732 33862
rect 32680 33798 32732 33804
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32692 33454 32720 33798
rect 32680 33448 32732 33454
rect 32680 33390 32732 33396
rect 32588 32972 32640 32978
rect 32588 32914 32640 32920
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32324 32230 32352 32846
rect 32312 32224 32364 32230
rect 32312 32166 32364 32172
rect 32220 31748 32272 31754
rect 32220 31690 32272 31696
rect 32232 31482 32260 31690
rect 32404 31680 32456 31686
rect 32324 31628 32404 31634
rect 32324 31622 32456 31628
rect 32324 31606 32444 31622
rect 32220 31476 32272 31482
rect 32220 31418 32272 31424
rect 32324 31414 32352 31606
rect 32312 31408 32364 31414
rect 32312 31350 32364 31356
rect 32324 30734 32352 31350
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32508 29850 32536 30194
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 32312 29504 32364 29510
rect 32312 29446 32364 29452
rect 32324 29238 32352 29446
rect 32312 29232 32364 29238
rect 32312 29174 32364 29180
rect 32416 28966 32444 29582
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 32508 29306 32536 29514
rect 32496 29300 32548 29306
rect 32496 29242 32548 29248
rect 32404 28960 32456 28966
rect 32404 28902 32456 28908
rect 32416 28762 32444 28902
rect 32404 28756 32456 28762
rect 32404 28698 32456 28704
rect 32600 28098 32628 32914
rect 32784 32366 32812 36790
rect 33968 36780 34020 36786
rect 33968 36722 34020 36728
rect 33416 36576 33468 36582
rect 33416 36518 33468 36524
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 33060 35834 33088 36178
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 32956 35080 33008 35086
rect 32956 35022 33008 35028
rect 32968 34542 32996 35022
rect 33048 34944 33100 34950
rect 33048 34886 33100 34892
rect 33060 34610 33088 34886
rect 33428 34678 33456 36518
rect 33980 36378 34008 36722
rect 34244 36712 34296 36718
rect 34244 36654 34296 36660
rect 33968 36372 34020 36378
rect 33968 36314 34020 36320
rect 34256 36242 34284 36654
rect 34244 36236 34296 36242
rect 34244 36178 34296 36184
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 33520 35290 33548 35634
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 33416 34672 33468 34678
rect 33416 34614 33468 34620
rect 33048 34604 33100 34610
rect 33048 34546 33100 34552
rect 32956 34536 33008 34542
rect 32956 34478 33008 34484
rect 33060 34354 33088 34546
rect 32968 34326 33088 34354
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32876 32026 32904 32370
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32968 31822 32996 34326
rect 33140 34196 33192 34202
rect 33140 34138 33192 34144
rect 33152 33522 33180 34138
rect 33232 34060 33284 34066
rect 33232 34002 33284 34008
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33140 33516 33192 33522
rect 33140 33458 33192 33464
rect 33060 33114 33088 33458
rect 33152 33153 33180 33458
rect 33138 33144 33194 33153
rect 33048 33108 33100 33114
rect 33138 33079 33194 33088
rect 33048 33050 33100 33056
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 32968 31482 32996 31758
rect 32956 31476 33008 31482
rect 32956 31418 33008 31424
rect 32680 30660 32732 30666
rect 32680 30602 32732 30608
rect 32692 30258 32720 30602
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 32692 29306 32720 30194
rect 33140 30048 33192 30054
rect 33140 29990 33192 29996
rect 33152 29578 33180 29990
rect 33140 29572 33192 29578
rect 33140 29514 33192 29520
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 33048 29232 33100 29238
rect 33048 29174 33100 29180
rect 33060 28558 33088 29174
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32508 28070 32628 28098
rect 32324 27674 32352 28018
rect 32312 27668 32364 27674
rect 32312 27610 32364 27616
rect 32220 27056 32272 27062
rect 32220 26998 32272 27004
rect 32232 25226 32260 26998
rect 32416 26042 32444 28018
rect 32404 26036 32456 26042
rect 32404 25978 32456 25984
rect 32312 25356 32364 25362
rect 32312 25298 32364 25304
rect 32220 25220 32272 25226
rect 32220 25162 32272 25168
rect 32232 23798 32260 25162
rect 32324 24206 32352 25298
rect 32508 25226 32536 28070
rect 32588 27940 32640 27946
rect 32588 27882 32640 27888
rect 32600 26994 32628 27882
rect 32956 27464 33008 27470
rect 32956 27406 33008 27412
rect 32968 27130 32996 27406
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 32496 25220 32548 25226
rect 32496 25162 32548 25168
rect 32404 24268 32456 24274
rect 32404 24210 32456 24216
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32220 23792 32272 23798
rect 32220 23734 32272 23740
rect 32324 23662 32352 24142
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32416 22658 32444 24210
rect 32508 24070 32536 25162
rect 32496 24064 32548 24070
rect 32496 24006 32548 24012
rect 32600 22778 32628 26930
rect 32680 26920 32732 26926
rect 32680 26862 32732 26868
rect 32692 26518 32720 26862
rect 32968 26858 32996 27066
rect 33060 26994 33088 28494
rect 33048 26988 33100 26994
rect 33048 26930 33100 26936
rect 32956 26852 33008 26858
rect 32956 26794 33008 26800
rect 32680 26512 32732 26518
rect 32680 26454 32732 26460
rect 33138 26480 33194 26489
rect 32692 24682 32720 26454
rect 33138 26415 33194 26424
rect 33152 25974 33180 26415
rect 33140 25968 33192 25974
rect 33140 25910 33192 25916
rect 32680 24676 32732 24682
rect 32680 24618 32732 24624
rect 32692 23497 32720 24618
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 32772 23520 32824 23526
rect 32678 23488 32734 23497
rect 32772 23462 32824 23468
rect 32678 23423 32734 23432
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32416 22630 32628 22658
rect 32496 22568 32548 22574
rect 32496 22510 32548 22516
rect 32312 22500 32364 22506
rect 32312 22442 32364 22448
rect 32324 22012 32352 22442
rect 32508 22030 32536 22510
rect 32600 22234 32628 22630
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32232 21984 32352 22012
rect 32496 22024 32548 22030
rect 32232 19854 32260 21984
rect 32496 21966 32548 21972
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32416 21622 32444 21830
rect 32404 21616 32456 21622
rect 32404 21558 32456 21564
rect 32508 19922 32536 21966
rect 32600 21146 32628 22170
rect 32680 21956 32732 21962
rect 32680 21898 32732 21904
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32692 20398 32720 21898
rect 32784 21554 32812 23462
rect 32876 22030 32904 23802
rect 33046 23760 33102 23769
rect 33046 23695 33048 23704
rect 33100 23695 33102 23704
rect 33048 23666 33100 23672
rect 33060 23118 33088 23666
rect 33048 23112 33100 23118
rect 33048 23054 33100 23060
rect 33048 22500 33100 22506
rect 33048 22442 33100 22448
rect 33060 22030 33088 22442
rect 33244 22098 33272 34002
rect 33428 33590 33456 34614
rect 34256 34610 34284 36178
rect 34520 36100 34572 36106
rect 34520 36042 34572 36048
rect 34532 35834 34560 36042
rect 34520 35828 34572 35834
rect 34520 35770 34572 35776
rect 34808 35193 34836 37726
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36636 37324 36688 37330
rect 36636 37266 36688 37272
rect 36648 36718 36676 37266
rect 38212 37262 38240 39200
rect 39026 38312 39082 38321
rect 39026 38247 39082 38256
rect 39040 37330 39068 38247
rect 39028 37324 39080 37330
rect 39028 37266 39080 37272
rect 36912 37256 36964 37262
rect 36912 37198 36964 37204
rect 38200 37256 38252 37262
rect 38200 37198 38252 37204
rect 36820 37188 36872 37194
rect 36820 37130 36872 37136
rect 36728 36780 36780 36786
rect 36728 36722 36780 36728
rect 36636 36712 36688 36718
rect 36636 36654 36688 36660
rect 35716 36576 35768 36582
rect 35716 36518 35768 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34794 35184 34850 35193
rect 35728 35154 35756 36518
rect 36360 36168 36412 36174
rect 36360 36110 36412 36116
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 34794 35119 34850 35128
rect 35716 35148 35768 35154
rect 35716 35090 35768 35096
rect 35900 35148 35952 35154
rect 35900 35090 35952 35096
rect 34796 35012 34848 35018
rect 34796 34954 34848 34960
rect 34244 34604 34296 34610
rect 34244 34546 34296 34552
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 33416 33584 33468 33590
rect 33416 33526 33468 33532
rect 34440 33522 34468 33594
rect 34808 33522 34836 34954
rect 35348 34400 35400 34406
rect 35348 34342 35400 34348
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 33862 35388 34342
rect 35716 34128 35768 34134
rect 35716 34070 35768 34076
rect 35348 33856 35400 33862
rect 35348 33798 35400 33804
rect 35530 33824 35586 33833
rect 34428 33516 34480 33522
rect 34704 33516 34756 33522
rect 34428 33458 34480 33464
rect 34532 33476 34704 33504
rect 34532 32570 34560 33476
rect 34704 33458 34756 33464
rect 34796 33516 34848 33522
rect 34796 33458 34848 33464
rect 34704 33380 34756 33386
rect 34704 33322 34756 33328
rect 34520 32564 34572 32570
rect 34520 32506 34572 32512
rect 34152 32224 34204 32230
rect 34152 32166 34204 32172
rect 34164 31278 34192 32166
rect 34334 31648 34390 31657
rect 34334 31583 34390 31592
rect 34348 31346 34376 31583
rect 34532 31346 34560 32506
rect 34716 32298 34744 33322
rect 34704 32292 34756 32298
rect 34704 32234 34756 32240
rect 34716 31346 34744 32234
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34164 31142 34192 31214
rect 34152 31136 34204 31142
rect 34152 31078 34204 31084
rect 33876 30796 33928 30802
rect 33876 30738 33928 30744
rect 33888 30326 33916 30738
rect 33876 30320 33928 30326
rect 33876 30262 33928 30268
rect 33324 30184 33376 30190
rect 33324 30126 33376 30132
rect 33336 29578 33364 30126
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33428 29646 33456 30058
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 34532 29578 34560 31282
rect 34612 29844 34664 29850
rect 34612 29786 34664 29792
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 34520 29572 34572 29578
rect 34520 29514 34572 29520
rect 33336 28014 33364 29514
rect 33506 29064 33562 29073
rect 33506 28999 33562 29008
rect 33416 28620 33468 28626
rect 33416 28562 33468 28568
rect 33428 28150 33456 28562
rect 33416 28144 33468 28150
rect 33416 28086 33468 28092
rect 33324 28008 33376 28014
rect 33324 27950 33376 27956
rect 33336 26926 33364 27950
rect 33416 27532 33468 27538
rect 33416 27474 33468 27480
rect 33428 26926 33456 27474
rect 33324 26920 33376 26926
rect 33324 26862 33376 26868
rect 33416 26920 33468 26926
rect 33416 26862 33468 26868
rect 33428 26450 33456 26862
rect 33416 26444 33468 26450
rect 33416 26386 33468 26392
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 33428 25294 33456 25638
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 33520 23730 33548 28999
rect 34624 28994 34652 29786
rect 34532 28966 34652 28994
rect 33876 28620 33928 28626
rect 33876 28562 33928 28568
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33612 27538 33640 28018
rect 33692 27600 33744 27606
rect 33692 27542 33744 27548
rect 33600 27532 33652 27538
rect 33600 27474 33652 27480
rect 33612 26518 33640 27474
rect 33704 27470 33732 27542
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 33600 26512 33652 26518
rect 33600 26454 33652 26460
rect 33704 26042 33732 27406
rect 33888 27402 33916 28562
rect 34244 28212 34296 28218
rect 34244 28154 34296 28160
rect 33968 27464 34020 27470
rect 33968 27406 34020 27412
rect 33876 27396 33928 27402
rect 33876 27338 33928 27344
rect 33888 27282 33916 27338
rect 33796 27254 33916 27282
rect 33692 26036 33744 26042
rect 33692 25978 33744 25984
rect 33796 25838 33824 27254
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 33888 25906 33916 26522
rect 33980 26382 34008 27406
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 34164 26518 34192 26930
rect 34256 26518 34284 28154
rect 34532 27470 34560 28966
rect 34808 27690 34836 33458
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35256 32428 35308 32434
rect 35256 32370 35308 32376
rect 35268 32298 35296 32370
rect 35256 32292 35308 32298
rect 35256 32234 35308 32240
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35256 31816 35308 31822
rect 35360 31804 35388 33798
rect 35530 33759 35586 33768
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 35452 32570 35480 32846
rect 35440 32564 35492 32570
rect 35440 32506 35492 32512
rect 35544 32502 35572 33759
rect 35728 33454 35756 34070
rect 35912 33522 35940 35090
rect 36096 34066 36124 35974
rect 36372 35154 36400 36110
rect 36740 35698 36768 36722
rect 36832 36378 36860 37130
rect 36820 36372 36872 36378
rect 36820 36314 36872 36320
rect 36924 35834 36952 37198
rect 39028 37120 39080 37126
rect 39028 37062 39080 37068
rect 39040 36961 39068 37062
rect 39026 36952 39082 36961
rect 39026 36887 39082 36896
rect 37924 36780 37976 36786
rect 37924 36722 37976 36728
rect 37464 36100 37516 36106
rect 37464 36042 37516 36048
rect 37476 35834 37504 36042
rect 37832 36032 37884 36038
rect 37832 35974 37884 35980
rect 36912 35828 36964 35834
rect 36912 35770 36964 35776
rect 37464 35828 37516 35834
rect 37464 35770 37516 35776
rect 37844 35698 37872 35974
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 37648 35692 37700 35698
rect 37648 35634 37700 35640
rect 37832 35692 37884 35698
rect 37832 35634 37884 35640
rect 36360 35148 36412 35154
rect 36360 35090 36412 35096
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 35992 33652 36044 33658
rect 35992 33594 36044 33600
rect 36004 33522 36032 33594
rect 35808 33516 35860 33522
rect 35808 33458 35860 33464
rect 35900 33516 35952 33522
rect 35900 33458 35952 33464
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 35716 33448 35768 33454
rect 35716 33390 35768 33396
rect 35820 33318 35848 33458
rect 35808 33312 35860 33318
rect 35808 33254 35860 33260
rect 35820 32774 35848 33254
rect 36096 32910 36124 34002
rect 36268 33516 36320 33522
rect 36268 33458 36320 33464
rect 36280 32910 36308 33458
rect 36372 32978 36400 35090
rect 36360 32972 36412 32978
rect 36360 32914 36412 32920
rect 36084 32904 36136 32910
rect 36084 32846 36136 32852
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 35808 32768 35860 32774
rect 35808 32710 35860 32716
rect 35900 32768 35952 32774
rect 35952 32728 36032 32756
rect 35900 32710 35952 32716
rect 35532 32496 35584 32502
rect 35532 32438 35584 32444
rect 35716 32496 35768 32502
rect 35716 32438 35768 32444
rect 35624 32360 35676 32366
rect 35624 32302 35676 32308
rect 35440 31816 35492 31822
rect 35360 31776 35440 31804
rect 35256 31758 35308 31764
rect 35440 31758 35492 31764
rect 35268 31482 35296 31758
rect 35256 31476 35308 31482
rect 35256 31418 35308 31424
rect 35348 31340 35400 31346
rect 35348 31282 35400 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29730 35388 31282
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 35452 29850 35480 30194
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 35360 29702 35480 29730
rect 35452 29646 35480 29702
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 35072 29572 35124 29578
rect 35072 29514 35124 29520
rect 35164 29572 35216 29578
rect 35164 29514 35216 29520
rect 35084 29238 35112 29514
rect 35072 29232 35124 29238
rect 35176 29209 35204 29514
rect 35348 29232 35400 29238
rect 35072 29174 35124 29180
rect 35162 29200 35218 29209
rect 35348 29174 35400 29180
rect 35162 29135 35218 29144
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34624 27662 34836 27690
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 34152 26512 34204 26518
rect 34152 26454 34204 26460
rect 34244 26512 34296 26518
rect 34244 26454 34296 26460
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 33876 25900 33928 25906
rect 33876 25842 33928 25848
rect 33784 25832 33836 25838
rect 33784 25774 33836 25780
rect 33600 25288 33652 25294
rect 33600 25230 33652 25236
rect 33612 23730 33640 25230
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33704 24274 33732 24754
rect 33796 24410 33824 25774
rect 34072 25158 34100 26318
rect 34060 25152 34112 25158
rect 34060 25094 34112 25100
rect 33876 24744 33928 24750
rect 33876 24686 33928 24692
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33692 24268 33744 24274
rect 33692 24210 33744 24216
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33612 23526 33640 23666
rect 33600 23520 33652 23526
rect 33600 23462 33652 23468
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33508 22636 33560 22642
rect 33508 22578 33560 22584
rect 33232 22092 33284 22098
rect 33232 22034 33284 22040
rect 33520 22030 33548 22578
rect 33612 22098 33640 22646
rect 33704 22574 33732 24210
rect 33888 24206 33916 24686
rect 34072 24206 34100 25094
rect 34256 24410 34284 26318
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 34060 24200 34112 24206
rect 34532 24177 34560 26386
rect 34624 24290 34652 27662
rect 34980 27464 35032 27470
rect 34980 27406 35032 27412
rect 34796 27056 34848 27062
rect 34796 26998 34848 27004
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34716 24410 34744 26930
rect 34808 25294 34836 26998
rect 34992 26858 35020 27406
rect 34980 26852 35032 26858
rect 34980 26794 35032 26800
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26382 35388 29174
rect 35452 29170 35480 29582
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35452 27606 35480 29106
rect 35532 28960 35584 28966
rect 35532 28902 35584 28908
rect 35544 28558 35572 28902
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 35440 27600 35492 27606
rect 35440 27542 35492 27548
rect 35532 27464 35584 27470
rect 35532 27406 35584 27412
rect 35544 26586 35572 27406
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 34980 26376 35032 26382
rect 35256 26376 35308 26382
rect 34980 26318 35032 26324
rect 35254 26344 35256 26353
rect 35348 26376 35400 26382
rect 35308 26344 35310 26353
rect 34992 26042 35020 26318
rect 35348 26318 35400 26324
rect 35254 26279 35310 26288
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34624 24262 34744 24290
rect 34060 24142 34112 24148
rect 34518 24168 34574 24177
rect 33888 23866 33916 24142
rect 34518 24103 34574 24112
rect 33876 23860 33928 23866
rect 33876 23802 33928 23808
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 33692 22568 33744 22574
rect 33692 22510 33744 22516
rect 33600 22092 33652 22098
rect 33600 22034 33652 22040
rect 34060 22092 34112 22098
rect 34060 22034 34112 22040
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 32496 19916 32548 19922
rect 32496 19858 32548 19864
rect 32220 19848 32272 19854
rect 32404 19848 32456 19854
rect 32220 19790 32272 19796
rect 32402 19816 32404 19825
rect 32456 19816 32458 19825
rect 32232 18766 32260 19790
rect 32402 19751 32458 19760
rect 32508 18834 32536 19858
rect 32784 19802 32812 21490
rect 32692 19774 32812 19802
rect 32692 19378 32720 19774
rect 32876 19718 32904 21966
rect 33520 20602 33548 21966
rect 33612 21418 33640 22034
rect 34072 21622 34100 22034
rect 34060 21616 34112 21622
rect 34060 21558 34112 21564
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 33600 21412 33652 21418
rect 33600 21354 33652 21360
rect 33508 20596 33560 20602
rect 33508 20538 33560 20544
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33244 19854 33272 20402
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33520 19922 33548 20334
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32956 19712 33008 19718
rect 32956 19654 33008 19660
rect 32680 19372 32732 19378
rect 32680 19314 32732 19320
rect 32680 18964 32732 18970
rect 32680 18906 32732 18912
rect 32496 18828 32548 18834
rect 32496 18770 32548 18776
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32220 18624 32272 18630
rect 32220 18566 32272 18572
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32048 16952 32168 16980
rect 31944 16584 31996 16590
rect 31944 16526 31996 16532
rect 32036 16448 32088 16454
rect 32036 16390 32088 16396
rect 32048 16182 32076 16390
rect 32036 16176 32088 16182
rect 32036 16118 32088 16124
rect 31760 16040 31812 16046
rect 31760 15982 31812 15988
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 32140 15314 32168 16952
rect 32232 15502 32260 18566
rect 32508 17746 32536 18770
rect 32692 18698 32720 18906
rect 32876 18714 32904 19654
rect 32968 19446 32996 19654
rect 32956 19440 33008 19446
rect 32956 19382 33008 19388
rect 33048 18760 33100 18766
rect 32876 18708 33048 18714
rect 32876 18702 33100 18708
rect 33138 18728 33194 18737
rect 32680 18692 32732 18698
rect 32680 18634 32732 18640
rect 32876 18686 33088 18702
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32312 17604 32364 17610
rect 32312 17546 32364 17552
rect 32324 16590 32352 17546
rect 32312 16584 32364 16590
rect 32312 16526 32364 16532
rect 32496 16584 32548 16590
rect 32496 16526 32548 16532
rect 32508 16250 32536 16526
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32600 16114 32628 17614
rect 32876 17610 32904 18686
rect 33138 18663 33140 18672
rect 33192 18663 33194 18672
rect 33140 18634 33192 18640
rect 33244 18426 33272 19790
rect 33520 19514 33548 19858
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33704 19446 33732 21422
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33692 19440 33744 19446
rect 33692 19382 33744 19388
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33508 19372 33560 19378
rect 33508 19314 33560 19320
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 33336 18086 33364 19314
rect 33520 18970 33548 19314
rect 33600 19168 33652 19174
rect 33600 19110 33652 19116
rect 33508 18964 33560 18970
rect 33508 18906 33560 18912
rect 33612 18358 33640 19110
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 33324 18080 33376 18086
rect 33324 18022 33376 18028
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32588 16108 32640 16114
rect 32588 16050 32640 16056
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 32600 15366 32628 16050
rect 32968 15910 32996 17818
rect 33048 17604 33100 17610
rect 33048 17546 33100 17552
rect 33060 17202 33088 17546
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 33520 16590 33548 18226
rect 33612 16658 33640 18294
rect 33692 17332 33744 17338
rect 33692 17274 33744 17280
rect 33600 16652 33652 16658
rect 33600 16594 33652 16600
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33048 16448 33100 16454
rect 33048 16390 33100 16396
rect 33060 16114 33088 16390
rect 33520 16250 33548 16526
rect 33508 16244 33560 16250
rect 33508 16186 33560 16192
rect 33704 16114 33732 17274
rect 33876 16652 33928 16658
rect 33876 16594 33928 16600
rect 33782 16144 33838 16153
rect 33048 16108 33100 16114
rect 33048 16050 33100 16056
rect 33692 16108 33744 16114
rect 33782 16079 33838 16088
rect 33692 16050 33744 16056
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 32876 15366 32904 15846
rect 32588 15360 32640 15366
rect 31772 15162 31800 15302
rect 32140 15286 32260 15314
rect 32588 15302 32640 15308
rect 32864 15360 32916 15366
rect 32864 15302 32916 15308
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 32232 14958 32260 15286
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31680 11558 31708 12106
rect 32232 12102 32260 14894
rect 32968 14550 32996 15846
rect 32956 14544 33008 14550
rect 32876 14492 32956 14498
rect 32876 14486 33008 14492
rect 32876 14470 32996 14486
rect 33060 14482 33088 16050
rect 33416 14952 33468 14958
rect 33416 14894 33468 14900
rect 33048 14476 33100 14482
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 12434 32352 13806
rect 32876 13394 32904 14470
rect 33048 14418 33100 14424
rect 33060 14362 33088 14418
rect 32968 14334 33088 14362
rect 32968 13462 32996 14334
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33244 13530 33272 13874
rect 33428 13841 33456 14894
rect 33704 14362 33732 16050
rect 33796 15910 33824 16079
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33888 15094 33916 16594
rect 33876 15088 33928 15094
rect 33876 15030 33928 15036
rect 33980 14890 34008 20334
rect 34164 19242 34192 23734
rect 34532 23730 34560 24103
rect 34612 23792 34664 23798
rect 34612 23734 34664 23740
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34532 21010 34560 22986
rect 34624 21622 34652 23734
rect 34716 23662 34744 24262
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34704 23656 34756 23662
rect 34704 23598 34756 23604
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34612 21616 34664 21622
rect 34612 21558 34664 21564
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 34624 20058 34652 21558
rect 34716 20942 34744 23122
rect 34808 21554 34836 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34612 20052 34664 20058
rect 34612 19994 34664 20000
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 34440 19378 34468 19858
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34152 19236 34204 19242
rect 34152 19178 34204 19184
rect 34716 17320 34744 20878
rect 34808 19854 34836 21490
rect 35360 21418 35388 23666
rect 35636 23526 35664 32302
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 35728 23066 35756 32438
rect 36004 31890 36032 32728
rect 35992 31884 36044 31890
rect 35992 31826 36044 31832
rect 36004 31754 36032 31826
rect 36280 31822 36308 32846
rect 36372 31890 36400 32914
rect 36544 32020 36596 32026
rect 36544 31962 36596 31968
rect 36360 31884 36412 31890
rect 36360 31826 36412 31832
rect 36268 31816 36320 31822
rect 36268 31758 36320 31764
rect 36004 31726 36124 31754
rect 35900 31680 35952 31686
rect 35900 31622 35952 31628
rect 35912 31346 35940 31622
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35992 31136 36044 31142
rect 35992 31078 36044 31084
rect 35900 30388 35952 30394
rect 35900 30330 35952 30336
rect 35912 28558 35940 30330
rect 36004 30258 36032 31078
rect 35992 30252 36044 30258
rect 35992 30194 36044 30200
rect 36096 30138 36124 31726
rect 36280 30258 36308 31758
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 36004 30122 36124 30138
rect 35992 30116 36124 30122
rect 36044 30110 36124 30116
rect 35992 30058 36044 30064
rect 36004 28694 36032 30058
rect 36280 29850 36308 30194
rect 36268 29844 36320 29850
rect 36268 29786 36320 29792
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 35992 28688 36044 28694
rect 35992 28630 36044 28636
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35808 26852 35860 26858
rect 35808 26794 35860 26800
rect 35820 23594 35848 26794
rect 35992 24608 36044 24614
rect 35992 24550 36044 24556
rect 36004 23730 36032 24550
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 35808 23588 35860 23594
rect 35808 23530 35860 23536
rect 35452 23038 35756 23066
rect 35452 21486 35480 23038
rect 35624 22976 35676 22982
rect 35624 22918 35676 22924
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 35544 21690 35572 21966
rect 35532 21684 35584 21690
rect 35532 21626 35584 21632
rect 35440 21480 35492 21486
rect 35440 21422 35492 21428
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35164 20052 35216 20058
rect 35164 19994 35216 20000
rect 35072 19916 35124 19922
rect 35072 19858 35124 19864
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 34808 18290 34836 19790
rect 35084 19174 35112 19858
rect 35176 19786 35204 19994
rect 35360 19854 35388 21354
rect 35636 20942 35664 22918
rect 35716 22228 35768 22234
rect 35716 22170 35768 22176
rect 35728 22098 35756 22170
rect 35716 22094 35768 22098
rect 35820 22094 35848 23530
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35716 22092 35848 22094
rect 35768 22066 35848 22092
rect 35716 22034 35768 22040
rect 35728 21026 35756 22034
rect 35808 22024 35860 22030
rect 35808 21966 35860 21972
rect 35820 21146 35848 21966
rect 35912 21894 35940 23462
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 35900 21888 35952 21894
rect 35900 21830 35952 21836
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35912 21078 35940 21830
rect 36004 21622 36032 21898
rect 35992 21616 36044 21622
rect 35992 21558 36044 21564
rect 35900 21072 35952 21078
rect 35728 20998 35848 21026
rect 35900 21014 35952 21020
rect 35624 20936 35676 20942
rect 35624 20878 35676 20884
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 35440 20460 35492 20466
rect 35440 20402 35492 20408
rect 35624 20460 35676 20466
rect 35624 20402 35676 20408
rect 35256 19848 35308 19854
rect 35254 19816 35256 19825
rect 35348 19848 35400 19854
rect 35308 19816 35310 19825
rect 35164 19780 35216 19786
rect 35348 19790 35400 19796
rect 35254 19751 35310 19760
rect 35164 19722 35216 19728
rect 35176 19281 35204 19722
rect 35452 19514 35480 20402
rect 35636 20058 35664 20402
rect 35624 20052 35676 20058
rect 35624 19994 35676 20000
rect 35622 19952 35678 19961
rect 35728 19938 35756 20810
rect 35820 20262 35848 20998
rect 35808 20256 35860 20262
rect 35808 20198 35860 20204
rect 35678 19910 35756 19938
rect 35622 19887 35678 19896
rect 35440 19508 35492 19514
rect 35440 19450 35492 19456
rect 35162 19272 35218 19281
rect 35218 19230 35388 19258
rect 35162 19207 35218 19216
rect 35072 19168 35124 19174
rect 35072 19110 35124 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18714 35388 19230
rect 35440 19168 35492 19174
rect 35440 19110 35492 19116
rect 35268 18686 35388 18714
rect 35268 18358 35296 18686
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35360 18358 35388 18566
rect 35256 18352 35308 18358
rect 35256 18294 35308 18300
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 34796 18284 34848 18290
rect 34796 18226 34848 18232
rect 35072 18284 35124 18290
rect 35072 18226 35124 18232
rect 35084 18193 35112 18226
rect 35070 18184 35126 18193
rect 35070 18119 35126 18128
rect 35268 18034 35296 18294
rect 35452 18290 35480 19110
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 35440 18148 35492 18154
rect 35440 18090 35492 18096
rect 35268 18006 35388 18034
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34440 17292 34744 17320
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33612 14334 33732 14362
rect 33612 13870 33640 14334
rect 33692 14272 33744 14278
rect 33692 14214 33744 14220
rect 33600 13864 33652 13870
rect 33414 13832 33470 13841
rect 33600 13806 33652 13812
rect 33414 13767 33470 13776
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 32956 13456 33008 13462
rect 32956 13398 33008 13404
rect 32864 13388 32916 13394
rect 32864 13330 32916 13336
rect 33244 13326 33272 13466
rect 33232 13320 33284 13326
rect 33232 13262 33284 13268
rect 33140 12844 33192 12850
rect 33140 12786 33192 12792
rect 33152 12434 33180 12786
rect 32324 12406 32444 12434
rect 32220 12096 32272 12102
rect 32220 12038 32272 12044
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 32324 11830 32352 12038
rect 32312 11824 32364 11830
rect 32312 11766 32364 11772
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31680 11218 31708 11494
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 31484 11008 31536 11014
rect 31484 10950 31536 10956
rect 31496 9654 31524 10950
rect 32232 10266 32260 11086
rect 32220 10260 32272 10266
rect 32220 10202 32272 10208
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32048 9722 32076 9998
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 31484 9648 31536 9654
rect 31484 9590 31536 9596
rect 32048 9110 32076 9658
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 31300 8560 31352 8566
rect 31300 8502 31352 8508
rect 31312 8106 31340 8502
rect 32140 8362 32168 9998
rect 32128 8356 32180 8362
rect 32128 8298 32180 8304
rect 31220 8090 31340 8106
rect 32416 8090 32444 12406
rect 33060 12406 33180 12434
rect 32772 12300 32824 12306
rect 32824 12260 32904 12288
rect 32772 12242 32824 12248
rect 32876 12170 32904 12260
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 32680 12096 32732 12102
rect 32680 12038 32732 12044
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 32692 11898 32720 12038
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 32784 9518 32812 12038
rect 33060 11558 33088 12406
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33060 10062 33088 11494
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 33152 11150 33180 11290
rect 33428 11286 33456 13767
rect 33704 13326 33732 14214
rect 33692 13320 33744 13326
rect 33692 13262 33744 13268
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 33796 12850 33824 13126
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33416 11280 33468 11286
rect 33416 11222 33468 11228
rect 33520 11150 33548 11834
rect 33140 11144 33192 11150
rect 33140 11086 33192 11092
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32968 9518 32996 9862
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32864 9512 32916 9518
rect 32864 9454 32916 9460
rect 32956 9512 33008 9518
rect 32956 9454 33008 9460
rect 31208 8084 31340 8090
rect 31260 8078 31340 8084
rect 32404 8084 32456 8090
rect 31208 8026 31260 8032
rect 32404 8026 32456 8032
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30760 5574 30788 6258
rect 30840 6248 30892 6254
rect 30840 6190 30892 6196
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30760 5370 30788 5510
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30852 4826 30880 6190
rect 32416 5778 32444 8026
rect 32784 7818 32812 9454
rect 32876 9178 32904 9454
rect 32864 9172 32916 9178
rect 32864 9114 32916 9120
rect 32968 8838 32996 9454
rect 33060 9042 33088 9998
rect 33152 9654 33180 11086
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 33968 10600 34020 10606
rect 33968 10542 34020 10548
rect 33784 10464 33836 10470
rect 33784 10406 33836 10412
rect 33796 10062 33824 10406
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33876 9988 33928 9994
rect 33876 9930 33928 9936
rect 33140 9648 33192 9654
rect 33140 9590 33192 9596
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 32956 8832 33008 8838
rect 32956 8774 33008 8780
rect 33796 8566 33824 8910
rect 33784 8560 33836 8566
rect 33784 8502 33836 8508
rect 32956 8492 33008 8498
rect 32956 8434 33008 8440
rect 32968 7886 32996 8434
rect 33048 8288 33100 8294
rect 33048 8230 33100 8236
rect 33060 8022 33088 8230
rect 33888 8090 33916 9930
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 32772 7812 32824 7818
rect 32772 7754 32824 7760
rect 32968 7426 32996 7822
rect 32784 7410 32996 7426
rect 32772 7404 32996 7410
rect 32824 7398 32996 7404
rect 32772 7346 32824 7352
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31772 5302 31800 5646
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 31760 5296 31812 5302
rect 31760 5238 31812 5244
rect 32600 5234 32628 5510
rect 32968 5302 32996 7398
rect 33060 6882 33088 7958
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33152 7002 33180 7414
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 33060 6866 33180 6882
rect 33060 6860 33192 6866
rect 33060 6854 33140 6860
rect 33140 6802 33192 6808
rect 33152 5778 33180 6802
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 32956 5296 33008 5302
rect 32956 5238 33008 5244
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 31208 5160 31260 5166
rect 31208 5102 31260 5108
rect 31220 4826 31248 5102
rect 30840 4820 30892 4826
rect 30840 4762 30892 4768
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 30852 4282 30880 4762
rect 32968 4690 32996 5238
rect 32956 4684 33008 4690
rect 32956 4626 33008 4632
rect 30840 4276 30892 4282
rect 30840 4218 30892 4224
rect 30564 4208 30616 4214
rect 30564 4150 30616 4156
rect 33152 4010 33180 5714
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33704 5370 33732 5646
rect 33692 5364 33744 5370
rect 33692 5306 33744 5312
rect 33416 4548 33468 4554
rect 33416 4490 33468 4496
rect 33428 4282 33456 4490
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33980 4162 34008 10542
rect 34164 10198 34192 10610
rect 34440 10198 34468 17292
rect 34900 17202 34928 17478
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34888 17196 34940 17202
rect 34888 17138 34940 17144
rect 34532 16182 34560 17138
rect 34716 16590 34744 17138
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 16794 34836 17070
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34704 16584 34756 16590
rect 34704 16526 34756 16532
rect 35072 16584 35124 16590
rect 35072 16526 35124 16532
rect 34612 16448 34664 16454
rect 34612 16390 34664 16396
rect 34520 16176 34572 16182
rect 34520 16118 34572 16124
rect 34520 14816 34572 14822
rect 34624 14804 34652 16390
rect 34716 15706 34744 16526
rect 34978 16416 35034 16425
rect 34978 16351 35034 16360
rect 34992 16046 35020 16351
rect 35084 16250 35112 16526
rect 35256 16516 35308 16522
rect 35360 16504 35388 18006
rect 35308 16476 35388 16504
rect 35256 16458 35308 16464
rect 35072 16244 35124 16250
rect 35072 16186 35124 16192
rect 35360 16114 35388 16476
rect 35452 16454 35480 18090
rect 35440 16448 35492 16454
rect 35438 16416 35440 16425
rect 35492 16416 35494 16425
rect 35438 16351 35494 16360
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 34980 16040 35032 16046
rect 34980 15982 35032 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34572 14776 34652 14804
rect 34520 14758 34572 14764
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34532 11898 34560 14486
rect 34612 13388 34664 13394
rect 34612 13330 34664 13336
rect 34624 12918 34652 13330
rect 34716 12986 34744 15642
rect 35438 15600 35494 15609
rect 35438 15535 35440 15544
rect 35492 15535 35494 15544
rect 35440 15506 35492 15512
rect 35348 15496 35400 15502
rect 35070 15464 35126 15473
rect 34980 15428 35032 15434
rect 35348 15438 35400 15444
rect 35070 15399 35072 15408
rect 34980 15370 35032 15376
rect 35124 15399 35126 15408
rect 35072 15370 35124 15376
rect 34992 15162 35020 15370
rect 34980 15156 35032 15162
rect 34980 15098 35032 15104
rect 35360 15026 35388 15438
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14414 35388 14962
rect 35452 14482 35480 15098
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 35544 14346 35572 18702
rect 35636 14550 35664 19887
rect 35820 18086 35848 20198
rect 36096 18902 36124 29582
rect 36176 29164 36228 29170
rect 36176 29106 36228 29112
rect 36188 28422 36216 29106
rect 36280 28558 36308 29786
rect 36372 29714 36400 31826
rect 36556 31482 36584 31962
rect 36544 31476 36596 31482
rect 36544 31418 36596 31424
rect 36740 30938 36768 35634
rect 37464 35012 37516 35018
rect 37464 34954 37516 34960
rect 37476 34746 37504 34954
rect 37464 34740 37516 34746
rect 37464 34682 37516 34688
rect 37660 34202 37688 35634
rect 37936 35630 37964 36722
rect 39028 36712 39080 36718
rect 39028 36654 39080 36660
rect 37924 35624 37976 35630
rect 37924 35566 37976 35572
rect 38016 35624 38068 35630
rect 39040 35601 39068 36654
rect 38016 35566 38068 35572
rect 39026 35592 39082 35601
rect 37740 34944 37792 34950
rect 37740 34886 37792 34892
rect 37752 34610 37780 34886
rect 37740 34604 37792 34610
rect 37740 34546 37792 34552
rect 37648 34196 37700 34202
rect 37648 34138 37700 34144
rect 37752 33454 37780 34546
rect 37832 34468 37884 34474
rect 37832 34410 37884 34416
rect 37844 33998 37872 34410
rect 37832 33992 37884 33998
rect 37832 33934 37884 33940
rect 37844 33658 37872 33934
rect 37832 33652 37884 33658
rect 37832 33594 37884 33600
rect 37936 33590 37964 35566
rect 38028 34542 38056 35566
rect 39026 35527 39082 35536
rect 38016 34536 38068 34542
rect 38016 34478 38068 34484
rect 37924 33584 37976 33590
rect 37924 33526 37976 33532
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 37740 33448 37792 33454
rect 37740 33390 37792 33396
rect 37096 33312 37148 33318
rect 37096 33254 37148 33260
rect 37108 32910 37136 33254
rect 37844 33114 37872 33458
rect 38028 33454 38056 34478
rect 38106 34232 38162 34241
rect 38106 34167 38162 34176
rect 38120 34066 38148 34167
rect 38108 34060 38160 34066
rect 38108 34002 38160 34008
rect 37924 33448 37976 33454
rect 37924 33390 37976 33396
rect 38016 33448 38068 33454
rect 38016 33390 38068 33396
rect 37832 33108 37884 33114
rect 37832 33050 37884 33056
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 37936 32774 37964 33390
rect 37924 32768 37976 32774
rect 37924 32710 37976 32716
rect 37936 32434 37964 32710
rect 37924 32428 37976 32434
rect 37924 32370 37976 32376
rect 36912 31748 36964 31754
rect 36912 31690 36964 31696
rect 36924 31482 36952 31690
rect 36912 31476 36964 31482
rect 36912 31418 36964 31424
rect 38028 31278 38056 33390
rect 38106 32872 38162 32881
rect 38106 32807 38162 32816
rect 38120 32502 38148 32807
rect 38108 32496 38160 32502
rect 38108 32438 38160 32444
rect 38106 31512 38162 31521
rect 38106 31447 38162 31456
rect 38120 31414 38148 31447
rect 38108 31408 38160 31414
rect 38108 31350 38160 31356
rect 38016 31272 38068 31278
rect 38016 31214 38068 31220
rect 36728 30932 36780 30938
rect 36728 30874 36780 30880
rect 37832 30728 37884 30734
rect 37832 30670 37884 30676
rect 37844 30122 37872 30670
rect 38028 30190 38056 31214
rect 39028 30660 39080 30666
rect 39028 30602 39080 30608
rect 38200 30320 38252 30326
rect 38200 30262 38252 30268
rect 38016 30184 38068 30190
rect 38016 30126 38068 30132
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 36360 29708 36412 29714
rect 36360 29650 36412 29656
rect 36372 28626 36400 29650
rect 37476 29646 37504 29990
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 38028 29238 38056 30126
rect 38212 29850 38240 30262
rect 39040 30161 39068 30602
rect 39026 30152 39082 30161
rect 39026 30087 39082 30096
rect 38200 29844 38252 29850
rect 38200 29786 38252 29792
rect 38016 29232 38068 29238
rect 38016 29174 38068 29180
rect 37556 29164 37608 29170
rect 37556 29106 37608 29112
rect 36360 28620 36412 28626
rect 36360 28562 36412 28568
rect 36268 28552 36320 28558
rect 36268 28494 36320 28500
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36188 28150 36216 28358
rect 36176 28144 36228 28150
rect 36176 28086 36228 28092
rect 36372 27062 36400 28562
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 37476 28218 37504 28426
rect 37464 28212 37516 28218
rect 37464 28154 37516 28160
rect 37568 27130 37596 29106
rect 37832 28416 37884 28422
rect 37832 28358 37884 28364
rect 37844 28218 37872 28358
rect 37832 28212 37884 28218
rect 37832 28154 37884 28160
rect 38028 28014 38056 29174
rect 39028 29096 39080 29102
rect 39028 29038 39080 29044
rect 39040 28801 39068 29038
rect 39026 28792 39082 28801
rect 39026 28727 39082 28736
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 38936 27532 38988 27538
rect 38936 27474 38988 27480
rect 38948 27441 38976 27474
rect 38934 27432 38990 27441
rect 37924 27396 37976 27402
rect 38934 27367 38990 27376
rect 39028 27396 39080 27402
rect 37924 27338 37976 27344
rect 39028 27338 39080 27344
rect 37936 27130 37964 27338
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 37924 27124 37976 27130
rect 37924 27066 37976 27072
rect 36360 27056 36412 27062
rect 36360 26998 36412 27004
rect 36268 26784 36320 26790
rect 36268 26726 36320 26732
rect 36280 25974 36308 26726
rect 36372 26450 36400 26998
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 36820 26784 36872 26790
rect 36820 26726 36872 26732
rect 36360 26444 36412 26450
rect 36360 26386 36412 26392
rect 36832 26382 36860 26726
rect 37844 26586 37872 26930
rect 38108 26920 38160 26926
rect 38108 26862 38160 26868
rect 37832 26580 37884 26586
rect 37832 26522 37884 26528
rect 36820 26376 36872 26382
rect 36820 26318 36872 26324
rect 36268 25968 36320 25974
rect 36268 25910 36320 25916
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 36728 25832 36780 25838
rect 36728 25774 36780 25780
rect 36740 25294 36768 25774
rect 36728 25288 36780 25294
rect 36728 25230 36780 25236
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36280 23322 36308 23666
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 36740 23118 36768 25230
rect 37464 25220 37516 25226
rect 37464 25162 37516 25168
rect 37476 24954 37504 25162
rect 37464 24948 37516 24954
rect 37464 24890 37516 24896
rect 37936 24750 37964 25842
rect 38016 25152 38068 25158
rect 38016 25094 38068 25100
rect 38028 24886 38056 25094
rect 38016 24880 38068 24886
rect 38016 24822 38068 24828
rect 38120 24750 38148 26862
rect 39040 26081 39068 27338
rect 39026 26072 39082 26081
rect 39026 26007 39082 26016
rect 39028 25832 39080 25838
rect 39028 25774 39080 25780
rect 37924 24744 37976 24750
rect 37924 24686 37976 24692
rect 38108 24744 38160 24750
rect 39040 24721 39068 25774
rect 38108 24686 38160 24692
rect 39026 24712 39082 24721
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37844 23866 37872 24142
rect 37936 24070 37964 24686
rect 37924 24064 37976 24070
rect 37924 24006 37976 24012
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 38120 23662 38148 24686
rect 39026 24647 39082 24656
rect 39028 24132 39080 24138
rect 39028 24074 39080 24080
rect 38200 23724 38252 23730
rect 38200 23666 38252 23672
rect 38108 23656 38160 23662
rect 38108 23598 38160 23604
rect 37096 23520 37148 23526
rect 37096 23462 37148 23468
rect 37108 23118 37136 23462
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 37096 23112 37148 23118
rect 37096 23054 37148 23060
rect 36740 22030 36768 23054
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36728 22024 36780 22030
rect 36728 21966 36780 21972
rect 36280 21690 36308 21966
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 36740 19854 36768 21966
rect 37464 21956 37516 21962
rect 37464 21898 37516 21904
rect 37476 21690 37504 21898
rect 37752 21894 37780 22578
rect 38120 22094 38148 23598
rect 38212 23322 38240 23666
rect 39040 23361 39068 24074
rect 39026 23352 39082 23361
rect 38200 23316 38252 23322
rect 39026 23287 39082 23296
rect 38200 23258 38252 23264
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 38028 22066 38148 22094
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37924 21888 37976 21894
rect 37924 21830 37976 21836
rect 37936 21690 37964 21830
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37924 21684 37976 21690
rect 37924 21626 37976 21632
rect 38028 21486 38056 22066
rect 39040 22001 39068 22510
rect 39026 21992 39082 22001
rect 39026 21927 39082 21936
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 38212 21622 38240 21830
rect 38200 21616 38252 21622
rect 38200 21558 38252 21564
rect 38016 21480 38068 21486
rect 38016 21422 38068 21428
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37752 20534 37780 20878
rect 37740 20528 37792 20534
rect 37740 20470 37792 20476
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37464 20256 37516 20262
rect 37464 20198 37516 20204
rect 37476 19854 37504 20198
rect 36728 19848 36780 19854
rect 36728 19790 36780 19796
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 36740 19446 36768 19790
rect 37844 19718 37872 20402
rect 38028 20398 38056 21422
rect 39028 20868 39080 20874
rect 39028 20810 39080 20816
rect 39040 20641 39068 20810
rect 39026 20632 39082 20641
rect 39026 20567 39082 20576
rect 38016 20392 38068 20398
rect 38016 20334 38068 20340
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 36728 19440 36780 19446
rect 36728 19382 36780 19388
rect 36084 18896 36136 18902
rect 36084 18838 36136 18844
rect 35900 18284 35952 18290
rect 35900 18226 35952 18232
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 35808 18080 35860 18086
rect 35808 18022 35860 18028
rect 35716 17196 35768 17202
rect 35716 17138 35768 17144
rect 35728 16998 35756 17138
rect 35820 17066 35848 18022
rect 35808 17060 35860 17066
rect 35808 17002 35860 17008
rect 35716 16992 35768 16998
rect 35716 16934 35768 16940
rect 35728 15858 35756 16934
rect 35728 15830 35848 15858
rect 35716 15360 35768 15366
rect 35716 15302 35768 15308
rect 35728 15026 35756 15302
rect 35716 15020 35768 15026
rect 35716 14962 35768 14968
rect 35716 14816 35768 14822
rect 35716 14758 35768 14764
rect 35624 14544 35676 14550
rect 35624 14486 35676 14492
rect 35728 14482 35756 14758
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35532 14340 35584 14346
rect 35532 14282 35584 14288
rect 35624 14340 35676 14346
rect 35624 14282 35676 14288
rect 35636 14006 35664 14282
rect 35624 14000 35676 14006
rect 35624 13942 35676 13948
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 34808 13326 34836 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34612 12912 34664 12918
rect 34612 12854 34664 12860
rect 34624 12238 34652 12854
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34624 11218 34652 12174
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 35360 11082 35388 12038
rect 35452 11694 35480 12038
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35452 11506 35480 11630
rect 35452 11478 35572 11506
rect 35544 11354 35572 11478
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35348 11076 35400 11082
rect 35348 11018 35400 11024
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 34532 10606 34560 10950
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34152 10192 34204 10198
rect 34152 10134 34204 10140
rect 34428 10192 34480 10198
rect 34428 10134 34480 10140
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 34520 9580 34572 9586
rect 34520 9522 34572 9528
rect 34244 8424 34296 8430
rect 34244 8366 34296 8372
rect 34256 7886 34284 8366
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 34072 6730 34100 7142
rect 34060 6724 34112 6730
rect 34060 6666 34112 6672
rect 34072 6390 34100 6666
rect 34060 6384 34112 6390
rect 34060 6326 34112 6332
rect 34256 6322 34284 7822
rect 34532 6390 34560 9522
rect 34704 9512 34756 9518
rect 34704 9454 34756 9460
rect 34716 8514 34744 9454
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34808 8634 34836 8774
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34716 8486 34836 8514
rect 34808 7410 34836 8486
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 35268 8242 35296 8434
rect 35268 8214 35388 8242
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 8090 35388 8214
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34612 7336 34664 7342
rect 34612 7278 34664 7284
rect 34520 6384 34572 6390
rect 34520 6326 34572 6332
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 5642 34284 6258
rect 34532 5642 34560 6326
rect 34624 6254 34652 7278
rect 34716 6458 34744 7346
rect 34808 6882 34836 7346
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34808 6854 34928 6882
rect 34704 6452 34756 6458
rect 34704 6394 34756 6400
rect 34900 6322 34928 6854
rect 35452 6458 35480 9998
rect 35636 9110 35664 13942
rect 35728 13394 35756 14418
rect 35716 13388 35768 13394
rect 35716 13330 35768 13336
rect 35820 13190 35848 15830
rect 35912 14804 35940 18226
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36004 15706 36032 17138
rect 36096 16250 36124 17138
rect 36084 16244 36136 16250
rect 36084 16186 36136 16192
rect 35992 15700 36044 15706
rect 35992 15642 36044 15648
rect 35992 14816 36044 14822
rect 35912 14776 35992 14804
rect 35992 14758 36044 14764
rect 36004 14618 36032 14758
rect 36372 14618 36400 18226
rect 36740 17678 36768 19382
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37568 18630 37596 19314
rect 38028 18834 38056 20334
rect 39028 19372 39080 19378
rect 39028 19314 39080 19320
rect 39040 19281 39068 19314
rect 39026 19272 39082 19281
rect 39026 19207 39082 19216
rect 38016 18828 38068 18834
rect 38016 18770 38068 18776
rect 37004 18624 37056 18630
rect 37004 18566 37056 18572
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37016 17678 37044 18566
rect 37568 18426 37596 18566
rect 37556 18420 37608 18426
rect 37556 18362 37608 18368
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 36728 17672 36780 17678
rect 36728 17614 36780 17620
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 36740 16658 36768 17614
rect 37740 17264 37792 17270
rect 37740 17206 37792 17212
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 37556 16584 37608 16590
rect 37556 16526 37608 16532
rect 37464 16516 37516 16522
rect 37464 16458 37516 16464
rect 37476 16250 37504 16458
rect 37464 16244 37516 16250
rect 37464 16186 37516 16192
rect 37568 15434 37596 16526
rect 37752 15570 37780 17206
rect 37844 17066 37872 18226
rect 37832 17060 37884 17066
rect 37832 17002 37884 17008
rect 37844 16250 37872 17002
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 38028 16046 38056 18770
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38120 17882 38148 18634
rect 39028 18216 39080 18222
rect 39028 18158 39080 18164
rect 39040 17921 39068 18158
rect 39026 17912 39082 17921
rect 38108 17876 38160 17882
rect 39026 17847 39082 17856
rect 38108 17818 38160 17824
rect 39028 17128 39080 17134
rect 39028 17070 39080 17076
rect 39040 16561 39068 17070
rect 39026 16552 39082 16561
rect 39026 16487 39082 16496
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 38120 16114 38148 16390
rect 38108 16108 38160 16114
rect 38108 16050 38160 16056
rect 38016 16040 38068 16046
rect 38016 15982 38068 15988
rect 38028 15638 38056 15982
rect 38016 15632 38068 15638
rect 38016 15574 38068 15580
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 37556 15428 37608 15434
rect 37556 15370 37608 15376
rect 37188 15360 37240 15366
rect 37188 15302 37240 15308
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 36360 14612 36412 14618
rect 36360 14554 36412 14560
rect 37200 14414 37228 15302
rect 37568 14618 37596 15370
rect 38106 15192 38162 15201
rect 38106 15127 38162 15136
rect 38120 15094 38148 15127
rect 38108 15088 38160 15094
rect 38108 15030 38160 15036
rect 37556 14612 37608 14618
rect 37556 14554 37608 14560
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 38292 13864 38344 13870
rect 38290 13832 38292 13841
rect 38344 13832 38346 13841
rect 38290 13767 38346 13776
rect 35808 13184 35860 13190
rect 35808 13126 35860 13132
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 38304 12481 38332 12582
rect 38290 12472 38346 12481
rect 38016 12436 38068 12442
rect 38290 12407 38346 12416
rect 38016 12378 38068 12384
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 35716 11756 35768 11762
rect 35716 11698 35768 11704
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35440 6452 35492 6458
rect 35440 6394 35492 6400
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34888 6316 34940 6322
rect 34888 6258 34940 6264
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34244 5636 34296 5642
rect 34244 5578 34296 5584
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34256 5302 34284 5578
rect 34808 5370 34836 6258
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35544 5914 35572 8910
rect 35728 7478 35756 11698
rect 35820 10606 35848 12242
rect 37924 12232 37976 12238
rect 37924 12174 37976 12180
rect 37464 12164 37516 12170
rect 37464 12106 37516 12112
rect 37476 11898 37504 12106
rect 37832 12096 37884 12102
rect 37832 12038 37884 12044
rect 37844 11898 37872 12038
rect 37936 11898 37964 12174
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 37924 11892 37976 11898
rect 37924 11834 37976 11840
rect 35992 11756 36044 11762
rect 35992 11698 36044 11704
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35820 7954 35848 10542
rect 36004 10062 36032 11698
rect 36268 11688 36320 11694
rect 36268 11630 36320 11636
rect 36280 11082 36308 11630
rect 36268 11076 36320 11082
rect 36268 11018 36320 11024
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 36280 10130 36308 11018
rect 37476 10810 37504 11018
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 37648 10736 37700 10742
rect 37648 10678 37700 10684
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37384 10130 37412 10610
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 37372 10124 37424 10130
rect 37372 10066 37424 10072
rect 35992 10056 36044 10062
rect 35992 9998 36044 10004
rect 36280 9178 36308 10066
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 36372 9654 36400 9998
rect 36360 9648 36412 9654
rect 36360 9590 36412 9596
rect 36268 9172 36320 9178
rect 36268 9114 36320 9120
rect 36268 9036 36320 9042
rect 36268 8978 36320 8984
rect 36280 8634 36308 8978
rect 36372 8974 36400 9590
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 36004 8022 36032 8366
rect 35992 8016 36044 8022
rect 35992 7958 36044 7964
rect 35808 7948 35860 7954
rect 35808 7890 35860 7896
rect 35716 7472 35768 7478
rect 35716 7414 35768 7420
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 34244 5296 34296 5302
rect 34244 5238 34296 5244
rect 34336 5228 34388 5234
rect 34336 5170 34388 5176
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 34348 4826 34376 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4826 35388 5170
rect 34336 4820 34388 4826
rect 34336 4762 34388 4768
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 34348 4282 34376 4762
rect 36004 4554 36032 7958
rect 36280 7886 36308 8570
rect 36820 8560 36872 8566
rect 36820 8502 36872 8508
rect 36832 7886 36860 8502
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37200 7886 37228 8298
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 36820 7880 36872 7886
rect 36820 7822 36872 7828
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 36832 6798 36860 7822
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36464 5370 36492 5646
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36464 4622 36492 5306
rect 36832 5302 36860 6734
rect 37464 6724 37516 6730
rect 37464 6666 37516 6672
rect 37476 6458 37504 6666
rect 37464 6452 37516 6458
rect 37464 6394 37516 6400
rect 37660 5302 37688 10678
rect 37830 10160 37886 10169
rect 37830 10095 37886 10104
rect 37844 10062 37872 10095
rect 37832 10056 37884 10062
rect 37832 9998 37884 10004
rect 37740 8900 37792 8906
rect 37740 8842 37792 8848
rect 37752 8634 37780 8842
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 37752 8106 37780 8570
rect 37752 8090 37872 8106
rect 37752 8084 37884 8090
rect 37752 8078 37832 8084
rect 37832 8026 37884 8032
rect 37740 7404 37792 7410
rect 37740 7346 37792 7352
rect 37752 7002 37780 7346
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37752 6458 37780 6938
rect 37936 6662 37964 11834
rect 38028 11694 38056 12378
rect 38016 11688 38068 11694
rect 38016 11630 38068 11636
rect 38028 10606 38056 11630
rect 39026 11112 39082 11121
rect 39026 11047 39082 11056
rect 38200 11008 38252 11014
rect 38200 10950 38252 10956
rect 38212 10674 38240 10950
rect 38200 10668 38252 10674
rect 38200 10610 38252 10616
rect 38016 10600 38068 10606
rect 38016 10542 38068 10548
rect 38028 8430 38056 10542
rect 39040 10130 39068 11047
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 39026 9752 39082 9761
rect 39026 9687 39082 9696
rect 39040 9654 39068 9687
rect 39028 9648 39080 9654
rect 39028 9590 39080 9596
rect 38108 8900 38160 8906
rect 38108 8842 38160 8848
rect 38016 8424 38068 8430
rect 38120 8401 38148 8842
rect 38016 8366 38068 8372
rect 38106 8392 38162 8401
rect 38106 8327 38162 8336
rect 38108 7336 38160 7342
rect 38108 7278 38160 7284
rect 38120 7041 38148 7278
rect 38106 7032 38162 7041
rect 38106 6967 38162 6976
rect 37924 6656 37976 6662
rect 37924 6598 37976 6604
rect 37936 6458 37964 6598
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37924 6452 37976 6458
rect 37924 6394 37976 6400
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 37752 5370 37780 6258
rect 38016 6248 38068 6254
rect 38016 6190 38068 6196
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 37844 5710 37872 6054
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 37740 5364 37792 5370
rect 37740 5306 37792 5312
rect 36820 5296 36872 5302
rect 36820 5238 36872 5244
rect 37648 5296 37700 5302
rect 37648 5238 37700 5244
rect 36832 4690 36860 5238
rect 37556 5092 37608 5098
rect 37556 5034 37608 5040
rect 37464 5024 37516 5030
rect 37464 4966 37516 4972
rect 36820 4684 36872 4690
rect 36820 4626 36872 4632
rect 37476 4622 37504 4966
rect 37568 4826 37596 5034
rect 37752 4826 37780 5306
rect 38028 5166 38056 6190
rect 38106 5672 38162 5681
rect 38106 5607 38108 5616
rect 38160 5607 38162 5616
rect 38108 5578 38160 5584
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 37556 4820 37608 4826
rect 37556 4762 37608 4768
rect 37740 4820 37792 4826
rect 37740 4762 37792 4768
rect 36452 4616 36504 4622
rect 36452 4558 36504 4564
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 35992 4548 36044 4554
rect 35992 4490 36044 4496
rect 39026 4312 39082 4321
rect 34336 4276 34388 4282
rect 39026 4247 39082 4256
rect 34336 4218 34388 4224
rect 33888 4146 34008 4162
rect 39040 4146 39068 4247
rect 33876 4140 34008 4146
rect 33928 4134 34008 4140
rect 39028 4140 39080 4146
rect 33876 4082 33928 4088
rect 39028 4082 39080 4088
rect 37830 4040 37886 4049
rect 33140 4004 33192 4010
rect 37830 3975 37886 3984
rect 33140 3946 33192 3952
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37844 3058 37872 3975
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 38108 2984 38160 2990
rect 38106 2952 38108 2961
rect 38160 2952 38162 2961
rect 38106 2887 38162 2896
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 38120 1601 38148 2314
rect 38106 1592 38162 1601
rect 38106 1527 38162 1536
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 5538 35944 5594 36000
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4986 28872 5042 28928
rect 4894 28600 4950 28656
rect 4710 27784 4766 27840
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 5630 27784 5686 27840
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 7102 27784 7158 27840
rect 8206 31356 8208 31376
rect 8208 31356 8260 31376
rect 8260 31356 8262 31376
rect 8206 31320 8262 31356
rect 8758 31320 8814 31376
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 12438 31864 12494 31920
rect 13726 32272 13782 32328
rect 13634 31340 13690 31376
rect 13634 31320 13636 31340
rect 13636 31320 13688 31340
rect 13688 31320 13690 31340
rect 13174 29144 13230 29200
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 15106 30096 15162 30152
rect 14646 20868 14702 20904
rect 14646 20848 14648 20868
rect 14648 20848 14700 20868
rect 14700 20848 14702 20868
rect 15198 26152 15254 26208
rect 16302 32428 16358 32464
rect 16302 32408 16304 32428
rect 16304 32408 16356 32428
rect 16356 32408 16358 32428
rect 15842 31864 15898 31920
rect 15290 20460 15346 20496
rect 15290 20440 15292 20460
rect 15292 20440 15344 20460
rect 15344 20440 15346 20460
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 16486 26152 16542 26208
rect 17314 30368 17370 30424
rect 17774 30116 17830 30152
rect 17774 30096 17776 30116
rect 17776 30096 17828 30116
rect 17828 30096 17830 30116
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 18786 33904 18842 33960
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 18970 31728 19026 31784
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19706 33360 19762 33416
rect 19614 33224 19670 33280
rect 19430 32716 19432 32736
rect 19432 32716 19484 32736
rect 19484 32716 19486 32736
rect 19430 32680 19486 32716
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19798 32000 19854 32056
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19522 31320 19578 31376
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20258 32972 20314 33008
rect 20258 32952 20260 32972
rect 20260 32952 20312 32972
rect 20312 32952 20314 32972
rect 20534 32952 20590 33008
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19614 26968 19670 27024
rect 19430 26288 19486 26344
rect 17866 24656 17922 24712
rect 18418 24556 18420 24576
rect 18420 24556 18472 24576
rect 18472 24556 18474 24576
rect 18418 24520 18474 24556
rect 17590 20848 17646 20904
rect 18326 20032 18382 20088
rect 18234 19388 18236 19408
rect 18236 19388 18288 19408
rect 18288 19388 18290 19408
rect 18234 19352 18290 19388
rect 16118 13268 16120 13288
rect 16120 13268 16172 13288
rect 16172 13268 16174 13288
rect 16118 13232 16174 13268
rect 17498 13268 17500 13288
rect 17500 13268 17552 13288
rect 17552 13268 17554 13288
rect 17498 13232 17554 13268
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20166 26288 20222 26344
rect 19246 20324 19302 20360
rect 19246 20304 19248 20324
rect 19248 20304 19300 20324
rect 19300 20304 19302 20324
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20994 31728 21050 31784
rect 20810 29008 20866 29064
rect 20718 28600 20774 28656
rect 21730 33360 21786 33416
rect 21362 31864 21418 31920
rect 21454 29960 21510 30016
rect 21638 29708 21694 29744
rect 21638 29688 21640 29708
rect 21640 29688 21692 29708
rect 21692 29688 21694 29708
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19430 20168 19486 20224
rect 20074 20304 20130 20360
rect 20074 20168 20130 20224
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20166 20032 20222 20088
rect 21454 26152 21510 26208
rect 20350 19352 20406 19408
rect 19246 18944 19302 19000
rect 19614 18844 19616 18864
rect 19616 18844 19668 18864
rect 19668 18844 19670 18864
rect 19614 18808 19670 18844
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20074 18964 20130 19000
rect 20074 18944 20076 18964
rect 20076 18944 20128 18964
rect 20128 18944 20130 18964
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20534 15444 20536 15464
rect 20536 15444 20588 15464
rect 20588 15444 20590 15464
rect 20534 15408 20590 15444
rect 20442 15000 20498 15056
rect 21178 19372 21234 19408
rect 21178 19352 21180 19372
rect 21180 19352 21232 19372
rect 21232 19352 21234 19372
rect 21638 26560 21694 26616
rect 21822 26424 21878 26480
rect 21638 26016 21694 26072
rect 21362 16088 21418 16144
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 22006 26696 22062 26752
rect 22006 26424 22062 26480
rect 22098 26016 22154 26072
rect 24858 36216 24914 36272
rect 22742 32716 22744 32736
rect 22744 32716 22796 32736
rect 22796 32716 22798 32736
rect 22742 32680 22798 32716
rect 22834 30540 22836 30560
rect 22836 30540 22888 30560
rect 22888 30540 22890 30560
rect 22834 30504 22890 30540
rect 23294 30640 23350 30696
rect 22374 21936 22430 21992
rect 22006 19796 22008 19816
rect 22008 19796 22060 19816
rect 22060 19796 22062 19816
rect 22006 19760 22062 19796
rect 22098 18128 22154 18184
rect 22742 29416 22798 29472
rect 22926 29280 22982 29336
rect 23110 28600 23166 28656
rect 23570 29960 23626 30016
rect 23018 26152 23074 26208
rect 23110 24812 23166 24848
rect 23110 24792 23112 24812
rect 23112 24792 23164 24812
rect 23164 24792 23166 24812
rect 22006 16088 22062 16144
rect 22006 14456 22062 14512
rect 21730 14356 21732 14376
rect 21732 14356 21784 14376
rect 21784 14356 21786 14376
rect 21730 14320 21786 14356
rect 23478 29008 23534 29064
rect 23754 31728 23810 31784
rect 24030 31728 24086 31784
rect 23662 26580 23718 26616
rect 23662 26560 23664 26580
rect 23664 26560 23716 26580
rect 23716 26560 23718 26580
rect 23478 24656 23534 24712
rect 23202 22072 23258 22128
rect 23478 23432 23534 23488
rect 24950 34992 25006 35048
rect 24306 29688 24362 29744
rect 25962 34992 26018 35048
rect 25410 33224 25466 33280
rect 25686 32272 25742 32328
rect 25042 29044 25044 29064
rect 25044 29044 25096 29064
rect 25096 29044 25098 29064
rect 25042 29008 25098 29044
rect 25226 29044 25228 29064
rect 25228 29044 25280 29064
rect 25280 29044 25282 29064
rect 25226 29008 25282 29044
rect 24950 26696 25006 26752
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 23386 20576 23442 20632
rect 24766 21120 24822 21176
rect 25410 26968 25466 27024
rect 25226 21972 25228 21992
rect 25228 21972 25280 21992
rect 25280 21972 25282 21992
rect 25226 21936 25282 21972
rect 24398 16224 24454 16280
rect 24306 16088 24362 16144
rect 23570 13912 23626 13968
rect 24122 15020 24178 15056
rect 24122 15000 24124 15020
rect 24124 15000 24176 15020
rect 24176 15000 24178 15020
rect 22098 6160 22154 6216
rect 26514 29280 26570 29336
rect 25502 20168 25558 20224
rect 25318 14320 25374 14376
rect 25594 13948 25596 13968
rect 25596 13948 25648 13968
rect 25648 13948 25650 13968
rect 25594 13912 25650 13948
rect 24950 11328 25006 11384
rect 25686 11348 25742 11384
rect 25686 11328 25688 11348
rect 25688 11328 25740 11348
rect 25740 11328 25742 11348
rect 26238 24928 26294 24984
rect 26422 20884 26424 20904
rect 26424 20884 26476 20904
rect 26476 20884 26478 20904
rect 26422 20848 26478 20884
rect 27250 31864 27306 31920
rect 27066 29452 27068 29472
rect 27068 29452 27120 29472
rect 27120 29452 27122 29472
rect 27066 29416 27122 29452
rect 27710 32408 27766 32464
rect 27618 27648 27674 27704
rect 27710 26968 27766 27024
rect 27526 24928 27582 24984
rect 26146 18808 26202 18864
rect 26054 15136 26110 15192
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 27526 23432 27582 23488
rect 27526 19896 27582 19952
rect 27986 26324 27988 26344
rect 27988 26324 28040 26344
rect 28040 26324 28042 26344
rect 27986 26288 28042 26324
rect 28262 30676 28264 30696
rect 28264 30676 28316 30696
rect 28316 30676 28318 30696
rect 28262 30640 28318 30676
rect 28262 29180 28264 29200
rect 28264 29180 28316 29200
rect 28316 29180 28318 29200
rect 28262 29144 28318 29180
rect 27894 24520 27950 24576
rect 28262 26288 28318 26344
rect 28170 24792 28226 24848
rect 27986 23296 28042 23352
rect 27986 21256 28042 21312
rect 30930 35028 30932 35048
rect 30932 35028 30984 35048
rect 30984 35028 30986 35048
rect 29826 33496 29882 33552
rect 29918 33088 29974 33144
rect 30102 33768 30158 33824
rect 28630 23976 28686 24032
rect 28998 24928 29054 24984
rect 28906 23976 28962 24032
rect 28262 21256 28318 21312
rect 28078 19896 28134 19952
rect 27894 19624 27950 19680
rect 28538 20712 28594 20768
rect 28722 22108 28724 22128
rect 28724 22108 28776 22128
rect 28776 22108 28778 22128
rect 28722 22072 28778 22108
rect 27618 12280 27674 12336
rect 27526 12044 27528 12064
rect 27528 12044 27580 12064
rect 27580 12044 27582 12064
rect 27526 12008 27582 12044
rect 28630 19896 28686 19952
rect 28446 19488 28502 19544
rect 28722 19624 28778 19680
rect 28630 19352 28686 19408
rect 28538 19080 28594 19136
rect 29090 20304 29146 20360
rect 29734 27512 29790 27568
rect 29642 20984 29698 21040
rect 29274 20032 29330 20088
rect 29090 19916 29146 19952
rect 29090 19896 29092 19916
rect 29092 19896 29144 19916
rect 29144 19896 29146 19916
rect 28998 19624 29054 19680
rect 29182 19660 29184 19680
rect 29184 19660 29236 19680
rect 29236 19660 29238 19680
rect 29182 19624 29238 19660
rect 28906 19488 28962 19544
rect 29090 19488 29146 19544
rect 29090 19388 29092 19408
rect 29092 19388 29144 19408
rect 29144 19388 29146 19408
rect 29090 19352 29146 19388
rect 27986 15136 28042 15192
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 28446 15136 28502 15192
rect 28354 15020 28410 15056
rect 28354 15000 28356 15020
rect 28356 15000 28408 15020
rect 28408 15000 28410 15020
rect 29274 19352 29330 19408
rect 29182 15544 29238 15600
rect 28998 13932 29054 13968
rect 28998 13912 29000 13932
rect 29000 13912 29052 13932
rect 29052 13912 29054 13932
rect 30102 30116 30158 30152
rect 30102 30096 30104 30116
rect 30104 30096 30156 30116
rect 30156 30096 30158 30116
rect 30102 29008 30158 29064
rect 30930 34992 30986 35028
rect 30470 31592 30526 31648
rect 30470 30776 30526 30832
rect 30746 31184 30802 31240
rect 30378 26288 30434 26344
rect 30010 22752 30066 22808
rect 30746 25744 30802 25800
rect 30378 21972 30380 21992
rect 30380 21972 30432 21992
rect 30432 21972 30434 21992
rect 30378 21936 30434 21972
rect 29734 20032 29790 20088
rect 30010 21120 30066 21176
rect 29734 13912 29790 13968
rect 29734 13812 29736 13832
rect 29736 13812 29788 13832
rect 29788 13812 29790 13832
rect 29734 13776 29790 13812
rect 30010 19624 30066 19680
rect 30102 19352 30158 19408
rect 30102 13932 30158 13968
rect 30102 13912 30104 13932
rect 30104 13912 30156 13932
rect 30156 13912 30158 13932
rect 31666 33768 31722 33824
rect 30930 29008 30986 29064
rect 31298 31048 31354 31104
rect 31206 29144 31262 29200
rect 31482 29452 31484 29472
rect 31484 29452 31536 29472
rect 31536 29452 31538 29472
rect 31482 29416 31538 29452
rect 31206 24148 31208 24168
rect 31208 24148 31260 24168
rect 31260 24148 31262 24168
rect 31206 24112 31262 24148
rect 30746 20848 30802 20904
rect 30654 20168 30710 20224
rect 30286 16652 30342 16688
rect 31022 19780 31078 19816
rect 31022 19760 31024 19780
rect 31024 19760 31076 19780
rect 31076 19760 31078 19780
rect 30286 16632 30288 16652
rect 30288 16632 30340 16652
rect 30340 16632 30342 16652
rect 30378 16360 30434 16416
rect 30930 16224 30986 16280
rect 30654 15408 30710 15464
rect 31114 14456 31170 14512
rect 31482 19216 31538 19272
rect 33138 33088 33194 33144
rect 33138 26424 33194 26480
rect 32678 23432 32734 23488
rect 33046 23724 33102 23760
rect 33046 23704 33048 23724
rect 33048 23704 33100 23724
rect 33100 23704 33102 23724
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 39026 38256 39082 38312
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34794 35128 34850 35184
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34334 31592 34390 31648
rect 33506 29008 33562 29064
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35530 33768 35586 33824
rect 39026 36896 39082 36952
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35162 29144 35218 29200
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35254 26324 35256 26344
rect 35256 26324 35308 26344
rect 35308 26324 35310 26344
rect 35254 26288 35310 26324
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34518 24112 34574 24168
rect 32402 19796 32404 19816
rect 32404 19796 32456 19816
rect 32456 19796 32458 19816
rect 32402 19760 32458 19796
rect 33138 18692 33194 18728
rect 33138 18672 33140 18692
rect 33140 18672 33192 18692
rect 33192 18672 33194 18692
rect 33782 16088 33838 16144
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35254 19796 35256 19816
rect 35256 19796 35308 19816
rect 35308 19796 35310 19816
rect 35254 19760 35310 19796
rect 35622 19896 35678 19952
rect 35162 19216 35218 19272
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35070 18128 35126 18184
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 33414 13776 33470 13832
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34978 16360 35034 16416
rect 35438 16396 35440 16416
rect 35440 16396 35492 16416
rect 35492 16396 35494 16416
rect 35438 16360 35494 16396
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35438 15564 35494 15600
rect 35438 15544 35440 15564
rect 35440 15544 35492 15564
rect 35492 15544 35494 15564
rect 35070 15428 35126 15464
rect 35070 15408 35072 15428
rect 35072 15408 35124 15428
rect 35124 15408 35126 15428
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 39026 35536 39082 35592
rect 38106 34176 38162 34232
rect 38106 32816 38162 32872
rect 38106 31456 38162 31512
rect 39026 30096 39082 30152
rect 39026 28736 39082 28792
rect 38934 27376 38990 27432
rect 39026 26016 39082 26072
rect 39026 24656 39082 24712
rect 39026 23296 39082 23352
rect 39026 21936 39082 21992
rect 39026 20576 39082 20632
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 39026 19216 39082 19272
rect 39026 17856 39082 17912
rect 39026 16496 39082 16552
rect 38106 15136 38162 15192
rect 38290 13812 38292 13832
rect 38292 13812 38344 13832
rect 38344 13812 38346 13832
rect 38290 13776 38346 13812
rect 38290 12416 38346 12472
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37830 10104 37886 10160
rect 39026 11056 39082 11112
rect 39026 9696 39082 9752
rect 38106 8336 38162 8392
rect 38106 6976 38162 7032
rect 38106 5636 38162 5672
rect 38106 5616 38108 5636
rect 38108 5616 38160 5636
rect 38160 5616 38162 5636
rect 39026 4256 39082 4312
rect 37830 3984 37886 4040
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38106 2932 38108 2952
rect 38108 2932 38160 2952
rect 38160 2932 38162 2952
rect 38106 2896 38162 2932
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38106 1536 38162 1592
<< metal3 >>
rect 39021 38314 39087 38317
rect 39200 38314 40000 38344
rect 39021 38312 40000 38314
rect 39021 38256 39026 38312
rect 39082 38256 40000 38312
rect 39021 38254 40000 38256
rect 39021 38251 39087 38254
rect 39200 38224 40000 38254
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 39021 36954 39087 36957
rect 39200 36954 40000 36984
rect 39021 36952 40000 36954
rect 39021 36896 39026 36952
rect 39082 36896 40000 36952
rect 39021 36894 40000 36896
rect 39021 36891 39087 36894
rect 39200 36864 40000 36894
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 20110 36212 20116 36276
rect 20180 36274 20186 36276
rect 24853 36274 24919 36277
rect 20180 36272 24919 36274
rect 20180 36216 24858 36272
rect 24914 36216 24919 36272
rect 20180 36214 24919 36216
rect 20180 36212 20186 36214
rect 24853 36211 24919 36214
rect 5533 36004 5599 36005
rect 5533 36000 5580 36004
rect 5644 36002 5650 36004
rect 5533 35944 5538 36000
rect 5533 35940 5580 35944
rect 5644 35942 5690 36002
rect 5644 35940 5650 35942
rect 5533 35939 5599 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 39021 35594 39087 35597
rect 39200 35594 40000 35624
rect 39021 35592 40000 35594
rect 39021 35536 39026 35592
rect 39082 35536 40000 35592
rect 39021 35534 40000 35536
rect 39021 35531 39087 35534
rect 39200 35504 40000 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 22502 35124 22508 35188
rect 22572 35186 22578 35188
rect 34789 35186 34855 35189
rect 22572 35184 34855 35186
rect 22572 35128 34794 35184
rect 34850 35128 34855 35184
rect 22572 35126 34855 35128
rect 22572 35124 22578 35126
rect 34789 35123 34855 35126
rect 24945 35050 25011 35053
rect 25262 35050 25268 35052
rect 24945 35048 25268 35050
rect 24945 34992 24950 35048
rect 25006 34992 25268 35048
rect 24945 34990 25268 34992
rect 24945 34987 25011 34990
rect 25262 34988 25268 34990
rect 25332 35050 25338 35052
rect 25957 35050 26023 35053
rect 30925 35052 30991 35053
rect 30925 35050 30972 35052
rect 25332 35048 26023 35050
rect 25332 34992 25962 35048
rect 26018 34992 26023 35048
rect 25332 34990 26023 34992
rect 30880 35048 30972 35050
rect 30880 34992 30930 35048
rect 30880 34990 30972 34992
rect 25332 34988 25338 34990
rect 25957 34987 26023 34990
rect 30925 34988 30972 34990
rect 31036 34988 31042 35052
rect 30925 34987 30991 34988
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 38101 34234 38167 34237
rect 39200 34234 40000 34264
rect 38101 34232 40000 34234
rect 38101 34176 38106 34232
rect 38162 34176 40000 34232
rect 38101 34174 40000 34176
rect 38101 34171 38167 34174
rect 39200 34144 40000 34174
rect 18781 33962 18847 33965
rect 18781 33960 31770 33962
rect 18781 33904 18786 33960
rect 18842 33904 31770 33960
rect 18781 33902 31770 33904
rect 18781 33899 18847 33902
rect 31710 33829 31770 33902
rect 30097 33828 30163 33829
rect 30046 33764 30052 33828
rect 30116 33826 30163 33828
rect 31661 33826 31770 33829
rect 35525 33826 35591 33829
rect 30116 33824 30208 33826
rect 30158 33768 30208 33824
rect 30116 33766 30208 33768
rect 31661 33824 35591 33826
rect 31661 33768 31666 33824
rect 31722 33768 35530 33824
rect 35586 33768 35591 33824
rect 31661 33766 35591 33768
rect 30116 33764 30163 33766
rect 30097 33763 30163 33764
rect 31661 33763 31727 33766
rect 35525 33763 35591 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 28390 33492 28396 33556
rect 28460 33554 28466 33556
rect 29821 33554 29887 33557
rect 28460 33552 29887 33554
rect 28460 33496 29826 33552
rect 29882 33496 29887 33552
rect 28460 33494 29887 33496
rect 28460 33492 28466 33494
rect 29821 33491 29887 33494
rect 19701 33418 19767 33421
rect 21725 33418 21791 33421
rect 19701 33416 21791 33418
rect 19701 33360 19706 33416
rect 19762 33360 21730 33416
rect 21786 33360 21791 33416
rect 19701 33358 21791 33360
rect 19701 33355 19767 33358
rect 21725 33355 21791 33358
rect 19609 33282 19675 33285
rect 25405 33282 25471 33285
rect 19609 33280 25471 33282
rect 19609 33224 19614 33280
rect 19670 33224 25410 33280
rect 25466 33224 25471 33280
rect 19609 33222 25471 33224
rect 19609 33219 19675 33222
rect 25405 33219 25471 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 29913 33146 29979 33149
rect 33133 33146 33199 33149
rect 29913 33144 33199 33146
rect 29913 33088 29918 33144
rect 29974 33088 33138 33144
rect 33194 33088 33199 33144
rect 29913 33086 33199 33088
rect 29913 33083 29979 33086
rect 33133 33083 33199 33086
rect 20253 33010 20319 33013
rect 20529 33010 20595 33013
rect 20253 33008 20595 33010
rect 20253 32952 20258 33008
rect 20314 32952 20534 33008
rect 20590 32952 20595 33008
rect 20253 32950 20595 32952
rect 20253 32947 20319 32950
rect 20529 32947 20595 32950
rect 38101 32874 38167 32877
rect 39200 32874 40000 32904
rect 38101 32872 40000 32874
rect 38101 32816 38106 32872
rect 38162 32816 40000 32872
rect 38101 32814 40000 32816
rect 38101 32811 38167 32814
rect 39200 32784 40000 32814
rect 19425 32740 19491 32741
rect 19374 32738 19380 32740
rect 19334 32678 19380 32738
rect 19444 32736 19491 32740
rect 19486 32680 19491 32736
rect 19374 32676 19380 32678
rect 19444 32676 19491 32680
rect 19425 32675 19491 32676
rect 22737 32738 22803 32741
rect 22870 32738 22876 32740
rect 22737 32736 22876 32738
rect 22737 32680 22742 32736
rect 22798 32680 22876 32736
rect 22737 32678 22876 32680
rect 22737 32675 22803 32678
rect 22870 32676 22876 32678
rect 22940 32676 22946 32740
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 16297 32466 16363 32469
rect 16430 32466 16436 32468
rect 16297 32464 16436 32466
rect 16297 32408 16302 32464
rect 16358 32408 16436 32464
rect 16297 32406 16436 32408
rect 16297 32403 16363 32406
rect 16430 32404 16436 32406
rect 16500 32466 16506 32468
rect 27705 32466 27771 32469
rect 27838 32466 27844 32468
rect 16500 32464 27844 32466
rect 16500 32408 27710 32464
rect 27766 32408 27844 32464
rect 16500 32406 27844 32408
rect 16500 32404 16506 32406
rect 27705 32403 27771 32406
rect 27838 32404 27844 32406
rect 27908 32404 27914 32468
rect 13721 32330 13787 32333
rect 25681 32330 25747 32333
rect 13721 32328 25747 32330
rect 13721 32272 13726 32328
rect 13782 32272 25686 32328
rect 25742 32272 25747 32328
rect 13721 32270 25747 32272
rect 13721 32267 13787 32270
rect 25681 32267 25747 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19793 32058 19859 32061
rect 20110 32058 20116 32060
rect 19793 32056 20116 32058
rect 19793 32000 19798 32056
rect 19854 32000 20116 32056
rect 19793 31998 20116 32000
rect 19793 31995 19859 31998
rect 20110 31996 20116 31998
rect 20180 31996 20186 32060
rect 12433 31922 12499 31925
rect 15837 31922 15903 31925
rect 12433 31920 15903 31922
rect 12433 31864 12438 31920
rect 12494 31864 15842 31920
rect 15898 31864 15903 31920
rect 12433 31862 15903 31864
rect 12433 31859 12499 31862
rect 15837 31859 15903 31862
rect 21357 31922 21423 31925
rect 27245 31922 27311 31925
rect 21357 31920 27311 31922
rect 21357 31864 21362 31920
rect 21418 31864 27250 31920
rect 27306 31864 27311 31920
rect 21357 31862 27311 31864
rect 21357 31859 21423 31862
rect 27245 31859 27311 31862
rect 18965 31786 19031 31789
rect 20989 31786 21055 31789
rect 18965 31784 21055 31786
rect 18965 31728 18970 31784
rect 19026 31728 20994 31784
rect 21050 31728 21055 31784
rect 18965 31726 21055 31728
rect 18965 31723 19031 31726
rect 20989 31723 21055 31726
rect 23749 31786 23815 31789
rect 24025 31786 24091 31789
rect 23749 31784 24091 31786
rect 23749 31728 23754 31784
rect 23810 31728 24030 31784
rect 24086 31728 24091 31784
rect 23749 31726 24091 31728
rect 23749 31723 23815 31726
rect 24025 31723 24091 31726
rect 30465 31650 30531 31653
rect 34329 31650 34395 31653
rect 30465 31648 34395 31650
rect 30465 31592 30470 31648
rect 30526 31592 34334 31648
rect 34390 31592 34395 31648
rect 30465 31590 34395 31592
rect 30465 31587 30531 31590
rect 34329 31587 34395 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 38101 31514 38167 31517
rect 39200 31514 40000 31544
rect 38101 31512 40000 31514
rect 38101 31456 38106 31512
rect 38162 31456 40000 31512
rect 38101 31454 40000 31456
rect 38101 31451 38167 31454
rect 39200 31424 40000 31454
rect 8201 31378 8267 31381
rect 8753 31378 8819 31381
rect 13629 31378 13695 31381
rect 8201 31376 13695 31378
rect 8201 31320 8206 31376
rect 8262 31320 8758 31376
rect 8814 31320 13634 31376
rect 13690 31320 13695 31376
rect 8201 31318 13695 31320
rect 8201 31315 8267 31318
rect 8753 31315 8819 31318
rect 13629 31315 13695 31318
rect 19374 31316 19380 31380
rect 19444 31378 19450 31380
rect 19517 31378 19583 31381
rect 19444 31376 19583 31378
rect 19444 31320 19522 31376
rect 19578 31320 19583 31376
rect 19444 31318 19583 31320
rect 19444 31316 19450 31318
rect 19517 31315 19583 31318
rect 30741 31244 30807 31245
rect 30741 31242 30788 31244
rect 30696 31240 30788 31242
rect 30696 31184 30746 31240
rect 30696 31182 30788 31184
rect 30741 31180 30788 31182
rect 30852 31180 30858 31244
rect 30741 31179 30807 31180
rect 31150 31044 31156 31108
rect 31220 31106 31226 31108
rect 31293 31106 31359 31109
rect 31220 31104 31359 31106
rect 31220 31048 31298 31104
rect 31354 31048 31359 31104
rect 31220 31046 31359 31048
rect 31220 31044 31226 31046
rect 31293 31043 31359 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 28574 30772 28580 30836
rect 28644 30834 28650 30836
rect 30465 30834 30531 30837
rect 28644 30832 30531 30834
rect 28644 30776 30470 30832
rect 30526 30776 30531 30832
rect 28644 30774 30531 30776
rect 28644 30772 28650 30774
rect 30465 30771 30531 30774
rect 23289 30698 23355 30701
rect 28257 30698 28323 30701
rect 23289 30696 28323 30698
rect 23289 30640 23294 30696
rect 23350 30640 28262 30696
rect 28318 30640 28323 30696
rect 23289 30638 28323 30640
rect 23289 30635 23355 30638
rect 28257 30635 28323 30638
rect 22829 30562 22895 30565
rect 23054 30562 23060 30564
rect 22829 30560 23060 30562
rect 22829 30504 22834 30560
rect 22890 30504 23060 30560
rect 22829 30502 23060 30504
rect 22829 30499 22895 30502
rect 23054 30500 23060 30502
rect 23124 30500 23130 30564
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 17309 30426 17375 30429
rect 17534 30426 17540 30428
rect 17309 30424 17540 30426
rect 17309 30368 17314 30424
rect 17370 30368 17540 30424
rect 17309 30366 17540 30368
rect 17309 30363 17375 30366
rect 17534 30364 17540 30366
rect 17604 30364 17610 30428
rect 15101 30154 15167 30157
rect 17769 30154 17835 30157
rect 15101 30152 17835 30154
rect 15101 30096 15106 30152
rect 15162 30096 17774 30152
rect 17830 30096 17835 30152
rect 15101 30094 17835 30096
rect 15101 30091 15167 30094
rect 17769 30091 17835 30094
rect 30097 30154 30163 30157
rect 30230 30154 30236 30156
rect 30097 30152 30236 30154
rect 30097 30096 30102 30152
rect 30158 30096 30236 30152
rect 30097 30094 30236 30096
rect 30097 30091 30163 30094
rect 30230 30092 30236 30094
rect 30300 30092 30306 30156
rect 39021 30154 39087 30157
rect 39200 30154 40000 30184
rect 39021 30152 40000 30154
rect 39021 30096 39026 30152
rect 39082 30096 40000 30152
rect 39021 30094 40000 30096
rect 39021 30091 39087 30094
rect 39200 30064 40000 30094
rect 21449 30018 21515 30021
rect 23565 30018 23631 30021
rect 21449 30016 23631 30018
rect 21449 29960 21454 30016
rect 21510 29960 23570 30016
rect 23626 29960 23631 30016
rect 21449 29958 23631 29960
rect 21449 29955 21515 29958
rect 23565 29955 23631 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 21633 29746 21699 29749
rect 24301 29746 24367 29749
rect 21633 29744 24367 29746
rect 21633 29688 21638 29744
rect 21694 29688 24306 29744
rect 24362 29688 24367 29744
rect 21633 29686 24367 29688
rect 21633 29683 21699 29686
rect 24301 29683 24367 29686
rect 22737 29474 22803 29477
rect 27061 29474 27127 29477
rect 31477 29476 31543 29477
rect 31477 29474 31524 29476
rect 22737 29472 27127 29474
rect 22737 29416 22742 29472
rect 22798 29416 27066 29472
rect 27122 29416 27127 29472
rect 22737 29414 27127 29416
rect 31432 29472 31524 29474
rect 31432 29416 31482 29472
rect 31432 29414 31524 29416
rect 22737 29411 22803 29414
rect 27061 29411 27127 29414
rect 31477 29412 31524 29414
rect 31588 29412 31594 29476
rect 31477 29411 31543 29412
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 22921 29338 22987 29341
rect 26509 29338 26575 29341
rect 22921 29336 26575 29338
rect 22921 29280 22926 29336
rect 22982 29280 26514 29336
rect 26570 29280 26575 29336
rect 22921 29278 26575 29280
rect 22921 29275 22987 29278
rect 26509 29275 26575 29278
rect 13169 29202 13235 29205
rect 28257 29202 28323 29205
rect 31201 29202 31267 29205
rect 35157 29202 35223 29205
rect 13169 29200 35223 29202
rect 13169 29144 13174 29200
rect 13230 29144 28262 29200
rect 28318 29144 31206 29200
rect 31262 29144 35162 29200
rect 35218 29144 35223 29200
rect 13169 29142 35223 29144
rect 13169 29139 13235 29142
rect 28257 29139 28323 29142
rect 31201 29139 31267 29142
rect 35157 29139 35223 29142
rect 20805 29066 20871 29069
rect 23473 29066 23539 29069
rect 20805 29064 23539 29066
rect 20805 29008 20810 29064
rect 20866 29008 23478 29064
rect 23534 29008 23539 29064
rect 20805 29006 23539 29008
rect 20805 29003 20871 29006
rect 23473 29003 23539 29006
rect 25037 29066 25103 29069
rect 25221 29066 25287 29069
rect 25037 29064 25287 29066
rect 25037 29008 25042 29064
rect 25098 29008 25226 29064
rect 25282 29008 25287 29064
rect 25037 29006 25287 29008
rect 25037 29003 25103 29006
rect 25221 29003 25287 29006
rect 29862 29004 29868 29068
rect 29932 29066 29938 29068
rect 30097 29066 30163 29069
rect 29932 29064 30163 29066
rect 29932 29008 30102 29064
rect 30158 29008 30163 29064
rect 29932 29006 30163 29008
rect 29932 29004 29938 29006
rect 30097 29003 30163 29006
rect 30925 29066 30991 29069
rect 33501 29066 33567 29069
rect 30925 29064 33567 29066
rect 30925 29008 30930 29064
rect 30986 29008 33506 29064
rect 33562 29008 33567 29064
rect 30925 29006 33567 29008
rect 30925 29003 30991 29006
rect 33501 29003 33567 29006
rect 4981 28930 5047 28933
rect 4981 28928 5090 28930
rect 4981 28872 4986 28928
rect 5042 28872 5090 28928
rect 4981 28867 5090 28872
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4889 28658 4955 28661
rect 5030 28658 5090 28867
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 39021 28794 39087 28797
rect 39200 28794 40000 28824
rect 39021 28792 40000 28794
rect 39021 28736 39026 28792
rect 39082 28736 40000 28792
rect 39021 28734 40000 28736
rect 39021 28731 39087 28734
rect 39200 28704 40000 28734
rect 4889 28656 5090 28658
rect 4889 28600 4894 28656
rect 4950 28600 5090 28656
rect 4889 28598 5090 28600
rect 20713 28658 20779 28661
rect 22870 28658 22876 28660
rect 20713 28656 22876 28658
rect 20713 28600 20718 28656
rect 20774 28600 22876 28656
rect 20713 28598 22876 28600
rect 4889 28595 4955 28598
rect 20713 28595 20779 28598
rect 22870 28596 22876 28598
rect 22940 28658 22946 28660
rect 23105 28658 23171 28661
rect 22940 28656 23171 28658
rect 22940 28600 23110 28656
rect 23166 28600 23171 28656
rect 22940 28598 23171 28600
rect 22940 28596 22946 28598
rect 23105 28595 23171 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4705 27842 4771 27845
rect 5625 27842 5691 27845
rect 7097 27842 7163 27845
rect 4705 27840 7163 27842
rect 4705 27784 4710 27840
rect 4766 27784 5630 27840
rect 5686 27784 7102 27840
rect 7158 27784 7163 27840
rect 4705 27782 7163 27784
rect 4705 27779 4771 27782
rect 5625 27779 5691 27782
rect 7097 27779 7163 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 25998 27644 26004 27708
rect 26068 27706 26074 27708
rect 27613 27706 27679 27709
rect 26068 27704 27679 27706
rect 26068 27648 27618 27704
rect 27674 27648 27679 27704
rect 26068 27646 27679 27648
rect 26068 27644 26074 27646
rect 27613 27643 27679 27646
rect 27838 27508 27844 27572
rect 27908 27570 27914 27572
rect 29729 27570 29795 27573
rect 27908 27568 29795 27570
rect 27908 27512 29734 27568
rect 29790 27512 29795 27568
rect 27908 27510 29795 27512
rect 27908 27508 27914 27510
rect 29729 27507 29795 27510
rect 38929 27434 38995 27437
rect 39200 27434 40000 27464
rect 38929 27432 40000 27434
rect 38929 27376 38934 27432
rect 38990 27376 40000 27432
rect 38929 27374 40000 27376
rect 38929 27371 38995 27374
rect 39200 27344 40000 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 19609 27026 19675 27029
rect 25405 27026 25471 27029
rect 27705 27026 27771 27029
rect 19609 27024 27771 27026
rect 19609 26968 19614 27024
rect 19670 26968 25410 27024
rect 25466 26968 27710 27024
rect 27766 26968 27771 27024
rect 19609 26966 27771 26968
rect 19609 26963 19675 26966
rect 25405 26963 25471 26966
rect 27705 26963 27771 26966
rect 22001 26754 22067 26757
rect 24945 26754 25011 26757
rect 22001 26752 25011 26754
rect 22001 26696 22006 26752
rect 22062 26696 24950 26752
rect 25006 26696 25011 26752
rect 22001 26694 25011 26696
rect 22001 26691 22067 26694
rect 24945 26691 25011 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 21633 26618 21699 26621
rect 23657 26618 23723 26621
rect 21633 26616 23723 26618
rect 21633 26560 21638 26616
rect 21694 26560 23662 26616
rect 23718 26560 23723 26616
rect 21633 26558 23723 26560
rect 21633 26555 21699 26558
rect 23657 26555 23723 26558
rect 21817 26482 21883 26485
rect 22001 26482 22067 26485
rect 31518 26482 31524 26484
rect 21817 26480 22067 26482
rect 21817 26424 21822 26480
rect 21878 26424 22006 26480
rect 22062 26424 22067 26480
rect 21817 26422 22067 26424
rect 21817 26419 21883 26422
rect 22001 26419 22067 26422
rect 28030 26422 31524 26482
rect 28030 26349 28090 26422
rect 31518 26420 31524 26422
rect 31588 26482 31594 26484
rect 33133 26482 33199 26485
rect 31588 26480 33199 26482
rect 31588 26424 33138 26480
rect 33194 26424 33199 26480
rect 31588 26422 33199 26424
rect 31588 26420 31594 26422
rect 33133 26419 33199 26422
rect 19425 26346 19491 26349
rect 20161 26346 20227 26349
rect 27981 26346 28090 26349
rect 19425 26344 28090 26346
rect 19425 26288 19430 26344
rect 19486 26288 20166 26344
rect 20222 26288 27986 26344
rect 28042 26288 28090 26344
rect 19425 26286 28090 26288
rect 28257 26346 28323 26349
rect 28390 26346 28396 26348
rect 28257 26344 28396 26346
rect 28257 26288 28262 26344
rect 28318 26288 28396 26344
rect 28257 26286 28396 26288
rect 19425 26283 19491 26286
rect 20161 26283 20227 26286
rect 27981 26283 28047 26286
rect 28257 26283 28323 26286
rect 28390 26284 28396 26286
rect 28460 26284 28466 26348
rect 30373 26346 30439 26349
rect 35249 26346 35315 26349
rect 30373 26344 35315 26346
rect 30373 26288 30378 26344
rect 30434 26288 35254 26344
rect 35310 26288 35315 26344
rect 30373 26286 35315 26288
rect 30373 26283 30439 26286
rect 35249 26283 35315 26286
rect 15193 26210 15259 26213
rect 16481 26212 16547 26213
rect 16430 26210 16436 26212
rect 15193 26208 16436 26210
rect 16500 26210 16547 26212
rect 21449 26210 21515 26213
rect 23013 26210 23079 26213
rect 16500 26208 16628 26210
rect 15193 26152 15198 26208
rect 15254 26152 16436 26208
rect 16542 26152 16628 26208
rect 15193 26150 16436 26152
rect 15193 26147 15259 26150
rect 16430 26148 16436 26150
rect 16500 26150 16628 26152
rect 21449 26208 23079 26210
rect 21449 26152 21454 26208
rect 21510 26152 23018 26208
rect 23074 26152 23079 26208
rect 21449 26150 23079 26152
rect 16500 26148 16547 26150
rect 16481 26147 16547 26148
rect 21449 26147 21515 26150
rect 23013 26147 23079 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 21633 26074 21699 26077
rect 22093 26074 22159 26077
rect 21633 26072 22159 26074
rect 21633 26016 21638 26072
rect 21694 26016 22098 26072
rect 22154 26016 22159 26072
rect 21633 26014 22159 26016
rect 21633 26011 21699 26014
rect 22093 26011 22159 26014
rect 39021 26074 39087 26077
rect 39200 26074 40000 26104
rect 39021 26072 40000 26074
rect 39021 26016 39026 26072
rect 39082 26016 40000 26072
rect 39021 26014 40000 26016
rect 39021 26011 39087 26014
rect 39200 25984 40000 26014
rect 30741 25802 30807 25805
rect 31150 25802 31156 25804
rect 30741 25800 31156 25802
rect 30741 25744 30746 25800
rect 30802 25744 31156 25800
rect 30741 25742 31156 25744
rect 30741 25739 30807 25742
rect 31150 25740 31156 25742
rect 31220 25740 31226 25804
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 26233 24986 26299 24989
rect 27521 24988 27587 24989
rect 26366 24986 26372 24988
rect 26233 24984 26372 24986
rect 26233 24928 26238 24984
rect 26294 24928 26372 24984
rect 26233 24926 26372 24928
rect 26233 24923 26299 24926
rect 26366 24924 26372 24926
rect 26436 24924 26442 24988
rect 27470 24986 27476 24988
rect 27430 24926 27476 24986
rect 27540 24984 27587 24988
rect 27582 24928 27587 24984
rect 27470 24924 27476 24926
rect 27540 24924 27587 24928
rect 28758 24924 28764 24988
rect 28828 24986 28834 24988
rect 28993 24986 29059 24989
rect 28828 24984 29059 24986
rect 28828 24928 28998 24984
rect 29054 24928 29059 24984
rect 28828 24926 29059 24928
rect 28828 24924 28834 24926
rect 27521 24923 27587 24924
rect 28993 24923 29059 24926
rect 17534 24788 17540 24852
rect 17604 24850 17610 24852
rect 23105 24850 23171 24853
rect 17604 24848 23171 24850
rect 17604 24792 23110 24848
rect 23166 24792 23171 24848
rect 17604 24790 23171 24792
rect 17604 24788 17610 24790
rect 23105 24787 23171 24790
rect 28165 24852 28231 24853
rect 28165 24848 28212 24852
rect 28276 24850 28282 24852
rect 28165 24792 28170 24848
rect 28165 24788 28212 24792
rect 28276 24790 28322 24850
rect 28276 24788 28282 24790
rect 28165 24787 28231 24788
rect 17861 24714 17927 24717
rect 23473 24714 23539 24717
rect 17861 24712 23539 24714
rect 17861 24656 17866 24712
rect 17922 24656 23478 24712
rect 23534 24656 23539 24712
rect 17861 24654 23539 24656
rect 17861 24651 17927 24654
rect 23473 24651 23539 24654
rect 39021 24714 39087 24717
rect 39200 24714 40000 24744
rect 39021 24712 40000 24714
rect 39021 24656 39026 24712
rect 39082 24656 40000 24712
rect 39021 24654 40000 24656
rect 39021 24651 39087 24654
rect 39200 24624 40000 24654
rect 18413 24578 18479 24581
rect 21214 24578 21220 24580
rect 18413 24576 21220 24578
rect 18413 24520 18418 24576
rect 18474 24520 21220 24576
rect 18413 24518 21220 24520
rect 18413 24515 18479 24518
rect 21214 24516 21220 24518
rect 21284 24516 21290 24580
rect 23238 24516 23244 24580
rect 23308 24578 23314 24580
rect 27889 24578 27955 24581
rect 28574 24578 28580 24580
rect 23308 24576 28580 24578
rect 23308 24520 27894 24576
rect 27950 24520 28580 24576
rect 23308 24518 28580 24520
rect 23308 24516 23314 24518
rect 27889 24515 27955 24518
rect 28574 24516 28580 24518
rect 28644 24516 28650 24580
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 31201 24170 31267 24173
rect 34513 24170 34579 24173
rect 31201 24168 34579 24170
rect 31201 24112 31206 24168
rect 31262 24112 34518 24168
rect 34574 24112 34579 24168
rect 31201 24110 34579 24112
rect 31201 24107 31267 24110
rect 34513 24107 34579 24110
rect 28625 24034 28691 24037
rect 28901 24034 28967 24037
rect 28625 24032 28967 24034
rect 28625 23976 28630 24032
rect 28686 23976 28906 24032
rect 28962 23976 28967 24032
rect 28625 23974 28967 23976
rect 28625 23971 28691 23974
rect 28901 23971 28967 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 30046 23700 30052 23764
rect 30116 23762 30122 23764
rect 33041 23762 33107 23765
rect 30116 23760 33107 23762
rect 30116 23704 33046 23760
rect 33102 23704 33107 23760
rect 30116 23702 33107 23704
rect 30116 23700 30122 23702
rect 33041 23699 33107 23702
rect 23473 23492 23539 23493
rect 23422 23428 23428 23492
rect 23492 23490 23539 23492
rect 27521 23490 27587 23493
rect 32673 23490 32739 23493
rect 23492 23488 23584 23490
rect 23534 23432 23584 23488
rect 23492 23430 23584 23432
rect 27521 23488 32739 23490
rect 27521 23432 27526 23488
rect 27582 23432 32678 23488
rect 32734 23432 32739 23488
rect 27521 23430 32739 23432
rect 23492 23428 23539 23430
rect 23473 23427 23539 23428
rect 27521 23427 27587 23430
rect 32673 23427 32739 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 27981 23356 28047 23357
rect 27981 23352 28028 23356
rect 28092 23354 28098 23356
rect 39021 23354 39087 23357
rect 39200 23354 40000 23384
rect 27981 23296 27986 23352
rect 27981 23292 28028 23296
rect 28092 23294 28138 23354
rect 39021 23352 40000 23354
rect 39021 23296 39026 23352
rect 39082 23296 40000 23352
rect 39021 23294 40000 23296
rect 28092 23292 28098 23294
rect 27981 23291 28047 23292
rect 39021 23291 39087 23294
rect 39200 23264 40000 23294
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 30005 22812 30071 22813
rect 30005 22810 30052 22812
rect 29960 22808 30052 22810
rect 29960 22752 30010 22808
rect 29960 22750 30052 22752
rect 30005 22748 30052 22750
rect 30116 22748 30122 22812
rect 30005 22747 30071 22748
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 23197 22130 23263 22133
rect 28717 22130 28783 22133
rect 23197 22128 28783 22130
rect 23197 22072 23202 22128
rect 23258 22072 28722 22128
rect 28778 22072 28783 22128
rect 23197 22070 28783 22072
rect 23197 22067 23263 22070
rect 28717 22067 28783 22070
rect 22369 21994 22435 21997
rect 25221 21996 25287 21997
rect 22502 21994 22508 21996
rect 22369 21992 22508 21994
rect 22369 21936 22374 21992
rect 22430 21936 22508 21992
rect 22369 21934 22508 21936
rect 22369 21931 22435 21934
rect 22502 21932 22508 21934
rect 22572 21932 22578 21996
rect 25221 21994 25268 21996
rect 25176 21992 25268 21994
rect 25176 21936 25226 21992
rect 25176 21934 25268 21936
rect 25221 21932 25268 21934
rect 25332 21932 25338 21996
rect 29862 21932 29868 21996
rect 29932 21994 29938 21996
rect 30373 21994 30439 21997
rect 29932 21992 30439 21994
rect 29932 21936 30378 21992
rect 30434 21936 30439 21992
rect 29932 21934 30439 21936
rect 29932 21932 29938 21934
rect 25221 21931 25287 21932
rect 30373 21931 30439 21934
rect 39021 21994 39087 21997
rect 39200 21994 40000 22024
rect 39021 21992 40000 21994
rect 39021 21936 39026 21992
rect 39082 21936 40000 21992
rect 39021 21934 40000 21936
rect 39021 21931 39087 21934
rect 39200 21904 40000 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 27981 21314 28047 21317
rect 28257 21314 28323 21317
rect 27981 21312 28323 21314
rect 27981 21256 27986 21312
rect 28042 21256 28262 21312
rect 28318 21256 28323 21312
rect 27981 21254 28323 21256
rect 27981 21251 28047 21254
rect 28257 21251 28323 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 24761 21178 24827 21181
rect 30005 21178 30071 21181
rect 24761 21176 30071 21178
rect 24761 21120 24766 21176
rect 24822 21120 30010 21176
rect 30066 21120 30071 21176
rect 24761 21118 30071 21120
rect 24761 21115 24827 21118
rect 30005 21115 30071 21118
rect 29637 21042 29703 21045
rect 30966 21042 30972 21044
rect 29637 21040 30972 21042
rect 29637 20984 29642 21040
rect 29698 20984 30972 21040
rect 29637 20982 30972 20984
rect 29637 20979 29703 20982
rect 30966 20980 30972 20982
rect 31036 20980 31042 21044
rect 14641 20906 14707 20909
rect 17585 20906 17651 20909
rect 14641 20904 17651 20906
rect 14641 20848 14646 20904
rect 14702 20848 17590 20904
rect 17646 20848 17651 20904
rect 14641 20846 17651 20848
rect 14641 20843 14707 20846
rect 17585 20843 17651 20846
rect 26417 20906 26483 20909
rect 30741 20906 30807 20909
rect 26417 20904 30807 20906
rect 26417 20848 26422 20904
rect 26478 20848 30746 20904
rect 30802 20848 30807 20904
rect 26417 20846 30807 20848
rect 26417 20843 26483 20846
rect 30741 20843 30807 20846
rect 28533 20772 28599 20773
rect 28533 20768 28580 20772
rect 28644 20770 28650 20772
rect 28533 20712 28538 20768
rect 28533 20708 28580 20712
rect 28644 20710 28690 20770
rect 28644 20708 28650 20710
rect 28533 20707 28599 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 23381 20636 23447 20637
rect 23381 20632 23428 20636
rect 23492 20634 23498 20636
rect 39021 20634 39087 20637
rect 39200 20634 40000 20664
rect 23381 20576 23386 20632
rect 23381 20572 23428 20576
rect 23492 20574 23538 20634
rect 39021 20632 40000 20634
rect 39021 20576 39026 20632
rect 39082 20576 40000 20632
rect 39021 20574 40000 20576
rect 23492 20572 23498 20574
rect 23381 20571 23447 20572
rect 39021 20571 39087 20574
rect 39200 20544 40000 20574
rect 5574 20436 5580 20500
rect 5644 20498 5650 20500
rect 15285 20498 15351 20501
rect 5644 20496 15351 20498
rect 5644 20440 15290 20496
rect 15346 20440 15351 20496
rect 5644 20438 15351 20440
rect 5644 20436 5650 20438
rect 15285 20435 15351 20438
rect 19241 20362 19307 20365
rect 20069 20362 20135 20365
rect 19241 20360 20135 20362
rect 19241 20304 19246 20360
rect 19302 20304 20074 20360
rect 20130 20304 20135 20360
rect 19241 20302 20135 20304
rect 19241 20299 19307 20302
rect 20069 20299 20135 20302
rect 29085 20364 29151 20365
rect 29085 20360 29132 20364
rect 29196 20362 29202 20364
rect 29085 20304 29090 20360
rect 29085 20300 29132 20304
rect 29196 20302 29242 20362
rect 29196 20300 29202 20302
rect 29085 20299 29151 20300
rect 19425 20226 19491 20229
rect 20069 20226 20135 20229
rect 19425 20224 20135 20226
rect 19425 20168 19430 20224
rect 19486 20168 20074 20224
rect 20130 20168 20135 20224
rect 19425 20166 20135 20168
rect 19425 20163 19491 20166
rect 20069 20163 20135 20166
rect 25497 20226 25563 20229
rect 30649 20226 30715 20229
rect 25497 20224 30715 20226
rect 25497 20168 25502 20224
rect 25558 20168 30654 20224
rect 30710 20168 30715 20224
rect 25497 20166 30715 20168
rect 25497 20163 25563 20166
rect 30649 20163 30715 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 18321 20090 18387 20093
rect 20161 20090 20227 20093
rect 18321 20088 20227 20090
rect 18321 20032 18326 20088
rect 18382 20032 20166 20088
rect 20222 20032 20227 20088
rect 18321 20030 20227 20032
rect 18321 20027 18387 20030
rect 20161 20027 20227 20030
rect 29269 20090 29335 20093
rect 29729 20090 29795 20093
rect 29269 20088 29795 20090
rect 29269 20032 29274 20088
rect 29330 20032 29734 20088
rect 29790 20032 29795 20088
rect 29269 20030 29795 20032
rect 29269 20027 29335 20030
rect 29729 20027 29795 20030
rect 27521 19954 27587 19957
rect 28073 19954 28139 19957
rect 28625 19954 28691 19957
rect 27521 19952 28691 19954
rect 27521 19896 27526 19952
rect 27582 19896 28078 19952
rect 28134 19896 28630 19952
rect 28686 19896 28691 19952
rect 27521 19894 28691 19896
rect 27521 19891 27587 19894
rect 28073 19891 28139 19894
rect 28625 19891 28691 19894
rect 29085 19954 29151 19957
rect 35617 19954 35683 19957
rect 29085 19952 35683 19954
rect 29085 19896 29090 19952
rect 29146 19896 35622 19952
rect 35678 19896 35683 19952
rect 29085 19894 35683 19896
rect 29085 19891 29151 19894
rect 35617 19891 35683 19894
rect 22001 19818 22067 19821
rect 31017 19818 31083 19821
rect 22001 19816 31083 19818
rect 22001 19760 22006 19816
rect 22062 19760 31022 19816
rect 31078 19760 31083 19816
rect 22001 19758 31083 19760
rect 22001 19755 22067 19758
rect 31017 19755 31083 19758
rect 32397 19818 32463 19821
rect 35249 19818 35315 19821
rect 32397 19816 35315 19818
rect 32397 19760 32402 19816
rect 32458 19760 35254 19816
rect 35310 19760 35315 19816
rect 32397 19758 35315 19760
rect 32397 19755 32463 19758
rect 35249 19755 35315 19758
rect 27889 19682 27955 19685
rect 28717 19682 28783 19685
rect 28993 19682 29059 19685
rect 27889 19680 29059 19682
rect 27889 19624 27894 19680
rect 27950 19624 28722 19680
rect 28778 19624 28998 19680
rect 29054 19624 29059 19680
rect 27889 19622 29059 19624
rect 27889 19619 27955 19622
rect 28717 19619 28783 19622
rect 28993 19619 29059 19622
rect 29177 19682 29243 19685
rect 30005 19682 30071 19685
rect 29177 19680 30071 19682
rect 29177 19624 29182 19680
rect 29238 19624 30010 19680
rect 30066 19624 30071 19680
rect 29177 19622 30071 19624
rect 29177 19619 29243 19622
rect 30005 19619 30071 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 28441 19546 28507 19549
rect 28901 19546 28967 19549
rect 28441 19544 28967 19546
rect 28441 19488 28446 19544
rect 28502 19488 28906 19544
rect 28962 19488 28967 19544
rect 28441 19486 28967 19488
rect 28441 19483 28507 19486
rect 28901 19483 28967 19486
rect 29085 19548 29151 19549
rect 29085 19544 29132 19548
rect 29196 19546 29202 19548
rect 29085 19488 29090 19544
rect 29085 19484 29132 19488
rect 29196 19486 29242 19546
rect 29196 19484 29202 19486
rect 29085 19483 29151 19484
rect 18229 19410 18295 19413
rect 20345 19410 20411 19413
rect 21173 19410 21239 19413
rect 18229 19408 21239 19410
rect 18229 19352 18234 19408
rect 18290 19352 20350 19408
rect 20406 19352 21178 19408
rect 21234 19352 21239 19408
rect 18229 19350 21239 19352
rect 18229 19347 18295 19350
rect 20345 19347 20411 19350
rect 21173 19347 21239 19350
rect 28625 19410 28691 19413
rect 29085 19410 29151 19413
rect 28625 19408 29151 19410
rect 28625 19352 28630 19408
rect 28686 19352 29090 19408
rect 29146 19352 29151 19408
rect 28625 19350 29151 19352
rect 28625 19347 28691 19350
rect 29085 19347 29151 19350
rect 29269 19410 29335 19413
rect 30097 19410 30163 19413
rect 29269 19408 30163 19410
rect 29269 19352 29274 19408
rect 29330 19352 30102 19408
rect 30158 19352 30163 19408
rect 29269 19350 30163 19352
rect 29269 19347 29335 19350
rect 30097 19347 30163 19350
rect 31477 19274 31543 19277
rect 35157 19274 35223 19277
rect 31477 19272 35223 19274
rect 31477 19216 31482 19272
rect 31538 19216 35162 19272
rect 35218 19216 35223 19272
rect 31477 19214 35223 19216
rect 31477 19211 31543 19214
rect 35157 19211 35223 19214
rect 39021 19274 39087 19277
rect 39200 19274 40000 19304
rect 39021 19272 40000 19274
rect 39021 19216 39026 19272
rect 39082 19216 40000 19272
rect 39021 19214 40000 19216
rect 39021 19211 39087 19214
rect 39200 19184 40000 19214
rect 28533 19138 28599 19141
rect 30782 19138 30788 19140
rect 28533 19136 30788 19138
rect 28533 19080 28538 19136
rect 28594 19080 30788 19136
rect 28533 19078 30788 19080
rect 28533 19075 28599 19078
rect 30782 19076 30788 19078
rect 30852 19076 30858 19140
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19241 19002 19307 19005
rect 20069 19002 20135 19005
rect 19241 19000 20135 19002
rect 19241 18944 19246 19000
rect 19302 18944 20074 19000
rect 20130 18944 20135 19000
rect 19241 18942 20135 18944
rect 19241 18939 19307 18942
rect 20069 18939 20135 18942
rect 19609 18866 19675 18869
rect 26141 18866 26207 18869
rect 19609 18864 26207 18866
rect 19609 18808 19614 18864
rect 19670 18808 26146 18864
rect 26202 18808 26207 18864
rect 19609 18806 26207 18808
rect 19609 18803 19675 18806
rect 26141 18803 26207 18806
rect 30230 18668 30236 18732
rect 30300 18730 30306 18732
rect 33133 18730 33199 18733
rect 30300 18728 33199 18730
rect 30300 18672 33138 18728
rect 33194 18672 33199 18728
rect 30300 18670 33199 18672
rect 30300 18668 30306 18670
rect 33133 18667 33199 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 22093 18188 22159 18189
rect 22093 18184 22140 18188
rect 22204 18186 22210 18188
rect 23238 18186 23244 18188
rect 22093 18128 22098 18184
rect 22093 18124 22140 18128
rect 22204 18126 23244 18186
rect 22204 18124 22210 18126
rect 23238 18124 23244 18126
rect 23308 18124 23314 18188
rect 34462 18124 34468 18188
rect 34532 18186 34538 18188
rect 35065 18186 35131 18189
rect 34532 18184 35131 18186
rect 34532 18128 35070 18184
rect 35126 18128 35131 18184
rect 34532 18126 35131 18128
rect 34532 18124 34538 18126
rect 22093 18123 22159 18124
rect 35065 18123 35131 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 39021 17914 39087 17917
rect 39200 17914 40000 17944
rect 39021 17912 40000 17914
rect 39021 17856 39026 17912
rect 39082 17856 40000 17912
rect 39021 17854 40000 17856
rect 39021 17851 39087 17854
rect 39200 17824 40000 17854
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 30281 16692 30347 16693
rect 30230 16690 30236 16692
rect 30190 16630 30236 16690
rect 30300 16688 30347 16692
rect 30342 16632 30347 16688
rect 30230 16628 30236 16630
rect 30300 16628 30347 16632
rect 30281 16627 30347 16628
rect 39021 16554 39087 16557
rect 39200 16554 40000 16584
rect 39021 16552 40000 16554
rect 39021 16496 39026 16552
rect 39082 16496 40000 16552
rect 39021 16494 40000 16496
rect 39021 16491 39087 16494
rect 39200 16464 40000 16494
rect 30373 16418 30439 16421
rect 34973 16418 35039 16421
rect 35433 16418 35499 16421
rect 30373 16416 35499 16418
rect 30373 16360 30378 16416
rect 30434 16360 34978 16416
rect 35034 16360 35438 16416
rect 35494 16360 35499 16416
rect 30373 16358 35499 16360
rect 30373 16355 30439 16358
rect 34973 16355 35039 16358
rect 35433 16355 35499 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 24393 16282 24459 16285
rect 26366 16282 26372 16284
rect 24393 16280 26372 16282
rect 24393 16224 24398 16280
rect 24454 16224 26372 16280
rect 24393 16222 26372 16224
rect 24393 16219 24459 16222
rect 26366 16220 26372 16222
rect 26436 16282 26442 16284
rect 30925 16282 30991 16285
rect 26436 16280 30991 16282
rect 26436 16224 30930 16280
rect 30986 16224 30991 16280
rect 26436 16222 30991 16224
rect 26436 16220 26442 16222
rect 30925 16219 30991 16222
rect 21357 16146 21423 16149
rect 22001 16146 22067 16149
rect 24301 16146 24367 16149
rect 33777 16146 33843 16149
rect 21357 16144 33843 16146
rect 21357 16088 21362 16144
rect 21418 16088 22006 16144
rect 22062 16088 24306 16144
rect 24362 16088 33782 16144
rect 33838 16088 33843 16144
rect 21357 16086 33843 16088
rect 21357 16083 21423 16086
rect 22001 16083 22067 16086
rect 24301 16083 24367 16086
rect 33777 16083 33843 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 29177 15602 29243 15605
rect 35433 15602 35499 15605
rect 29177 15600 35499 15602
rect 29177 15544 29182 15600
rect 29238 15544 35438 15600
rect 35494 15544 35499 15600
rect 29177 15542 35499 15544
rect 29177 15539 29243 15542
rect 35433 15539 35499 15542
rect 20529 15466 20595 15469
rect 23054 15466 23060 15468
rect 20529 15464 23060 15466
rect 20529 15408 20534 15464
rect 20590 15408 23060 15464
rect 20529 15406 23060 15408
rect 20529 15403 20595 15406
rect 23054 15404 23060 15406
rect 23124 15404 23130 15468
rect 30649 15466 30715 15469
rect 35065 15466 35131 15469
rect 30649 15464 35131 15466
rect 30649 15408 30654 15464
rect 30710 15408 35070 15464
rect 35126 15408 35131 15464
rect 30649 15406 35131 15408
rect 30649 15403 30715 15406
rect 35065 15403 35131 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 26049 15196 26115 15197
rect 25998 15194 26004 15196
rect 25958 15134 26004 15194
rect 26068 15192 26115 15196
rect 26110 15136 26115 15192
rect 25998 15132 26004 15134
rect 26068 15132 26115 15136
rect 26049 15131 26115 15132
rect 27981 15194 28047 15197
rect 28206 15194 28212 15196
rect 27981 15192 28212 15194
rect 27981 15136 27986 15192
rect 28042 15136 28212 15192
rect 27981 15134 28212 15136
rect 27981 15131 28047 15134
rect 28206 15132 28212 15134
rect 28276 15132 28282 15196
rect 28441 15194 28507 15197
rect 28758 15194 28764 15196
rect 28441 15192 28764 15194
rect 28441 15136 28446 15192
rect 28502 15136 28764 15192
rect 28441 15134 28764 15136
rect 28441 15131 28507 15134
rect 28758 15132 28764 15134
rect 28828 15132 28834 15196
rect 38101 15194 38167 15197
rect 39200 15194 40000 15224
rect 38101 15192 40000 15194
rect 38101 15136 38106 15192
rect 38162 15136 40000 15192
rect 38101 15134 40000 15136
rect 38101 15131 38167 15134
rect 39200 15104 40000 15134
rect 20437 15058 20503 15061
rect 24117 15058 24183 15061
rect 28349 15060 28415 15061
rect 28349 15058 28396 15060
rect 20437 15056 24183 15058
rect 20437 15000 20442 15056
rect 20498 15000 24122 15056
rect 24178 15000 24183 15056
rect 20437 14998 24183 15000
rect 28304 15056 28396 15058
rect 28304 15000 28354 15056
rect 28304 14998 28396 15000
rect 20437 14995 20503 14998
rect 24117 14995 24183 14998
rect 28349 14996 28396 14998
rect 28460 14996 28466 15060
rect 28349 14995 28415 14996
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 22001 14514 22067 14517
rect 31109 14514 31175 14517
rect 22001 14512 31770 14514
rect 22001 14456 22006 14512
rect 22062 14456 31114 14512
rect 31170 14456 31770 14512
rect 22001 14454 31770 14456
rect 22001 14451 22067 14454
rect 31109 14451 31175 14454
rect 21725 14378 21791 14381
rect 25313 14378 25379 14381
rect 21725 14376 25379 14378
rect 21725 14320 21730 14376
rect 21786 14320 25318 14376
rect 25374 14320 25379 14376
rect 21725 14318 25379 14320
rect 21725 14315 21791 14318
rect 25313 14315 25379 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 23565 13970 23631 13973
rect 25589 13970 25655 13973
rect 23565 13968 25655 13970
rect 23565 13912 23570 13968
rect 23626 13912 25594 13968
rect 25650 13912 25655 13968
rect 23565 13910 25655 13912
rect 23565 13907 23631 13910
rect 25589 13907 25655 13910
rect 28993 13970 29059 13973
rect 29729 13970 29795 13973
rect 30097 13970 30163 13973
rect 28993 13968 30163 13970
rect 28993 13912 28998 13968
rect 29054 13912 29734 13968
rect 29790 13912 30102 13968
rect 30158 13912 30163 13968
rect 28993 13910 30163 13912
rect 31710 13970 31770 14454
rect 34462 13970 34468 13972
rect 31710 13910 34468 13970
rect 28993 13907 29059 13910
rect 29729 13907 29795 13910
rect 30097 13907 30163 13910
rect 34462 13908 34468 13910
rect 34532 13908 34538 13972
rect 29729 13834 29795 13837
rect 33409 13834 33475 13837
rect 29729 13832 33475 13834
rect 29729 13776 29734 13832
rect 29790 13776 33414 13832
rect 33470 13776 33475 13832
rect 29729 13774 33475 13776
rect 29729 13771 29795 13774
rect 33409 13771 33475 13774
rect 38285 13834 38351 13837
rect 39200 13834 40000 13864
rect 38285 13832 40000 13834
rect 38285 13776 38290 13832
rect 38346 13776 40000 13832
rect 38285 13774 40000 13776
rect 38285 13771 38351 13774
rect 39200 13744 40000 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 16113 13290 16179 13293
rect 17493 13290 17559 13293
rect 16113 13288 17559 13290
rect 16113 13232 16118 13288
rect 16174 13232 17498 13288
rect 17554 13232 17559 13288
rect 16113 13230 17559 13232
rect 16113 13227 16179 13230
rect 17493 13227 17559 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38285 12474 38351 12477
rect 39200 12474 40000 12504
rect 38285 12472 40000 12474
rect 38285 12416 38290 12472
rect 38346 12416 40000 12472
rect 38285 12414 40000 12416
rect 38285 12411 38351 12414
rect 39200 12384 40000 12414
rect 27470 12276 27476 12340
rect 27540 12338 27546 12340
rect 27613 12338 27679 12341
rect 27540 12336 27679 12338
rect 27540 12280 27618 12336
rect 27674 12280 27679 12336
rect 27540 12278 27679 12280
rect 27540 12276 27546 12278
rect 27613 12275 27679 12278
rect 22134 12004 22140 12068
rect 22204 12066 22210 12068
rect 27521 12066 27587 12069
rect 22204 12064 27587 12066
rect 22204 12008 27526 12064
rect 27582 12008 27587 12064
rect 22204 12006 27587 12008
rect 22204 12004 22210 12006
rect 27521 12003 27587 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 21214 11324 21220 11388
rect 21284 11386 21290 11388
rect 24945 11386 25011 11389
rect 25681 11386 25747 11389
rect 21284 11384 25747 11386
rect 21284 11328 24950 11384
rect 25006 11328 25686 11384
rect 25742 11328 25747 11384
rect 21284 11326 25747 11328
rect 21284 11324 21290 11326
rect 24945 11323 25011 11326
rect 25681 11323 25747 11326
rect 39021 11114 39087 11117
rect 39200 11114 40000 11144
rect 39021 11112 40000 11114
rect 39021 11056 39026 11112
rect 39082 11056 40000 11112
rect 39021 11054 40000 11056
rect 39021 11051 39087 11054
rect 39200 11024 40000 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 28574 10100 28580 10164
rect 28644 10162 28650 10164
rect 37825 10162 37891 10165
rect 28644 10160 37891 10162
rect 28644 10104 37830 10160
rect 37886 10104 37891 10160
rect 28644 10102 37891 10104
rect 28644 10100 28650 10102
rect 37825 10099 37891 10102
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 39021 9754 39087 9757
rect 39200 9754 40000 9784
rect 39021 9752 40000 9754
rect 39021 9696 39026 9752
rect 39082 9696 40000 9752
rect 39021 9694 40000 9696
rect 39021 9691 39087 9694
rect 39200 9664 40000 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 38101 8394 38167 8397
rect 39200 8394 40000 8424
rect 38101 8392 40000 8394
rect 38101 8336 38106 8392
rect 38162 8336 40000 8392
rect 38101 8334 40000 8336
rect 38101 8331 38167 8334
rect 39200 8304 40000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 38101 7034 38167 7037
rect 39200 7034 40000 7064
rect 38101 7032 40000 7034
rect 38101 6976 38106 7032
rect 38162 6976 40000 7032
rect 38101 6974 40000 6976
rect 38101 6971 38167 6974
rect 39200 6944 40000 6974
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 22093 6220 22159 6221
rect 22093 6216 22140 6220
rect 22204 6218 22210 6220
rect 22093 6160 22098 6216
rect 22093 6156 22140 6160
rect 22204 6158 22250 6218
rect 22204 6156 22210 6158
rect 22093 6155 22159 6156
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38101 5674 38167 5677
rect 39200 5674 40000 5704
rect 38101 5672 40000 5674
rect 38101 5616 38106 5672
rect 38162 5616 40000 5672
rect 38101 5614 40000 5616
rect 38101 5611 38167 5614
rect 39200 5584 40000 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 39021 4314 39087 4317
rect 39200 4314 40000 4344
rect 39021 4312 40000 4314
rect 39021 4256 39026 4312
rect 39082 4256 40000 4312
rect 39021 4254 40000 4256
rect 39021 4251 39087 4254
rect 39200 4224 40000 4254
rect 30230 3980 30236 4044
rect 30300 4042 30306 4044
rect 37825 4042 37891 4045
rect 30300 4040 37891 4042
rect 30300 3984 37830 4040
rect 37886 3984 37891 4040
rect 30300 3982 37891 3984
rect 30300 3980 30306 3982
rect 37825 3979 37891 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 38101 2954 38167 2957
rect 39200 2954 40000 2984
rect 38101 2952 40000 2954
rect 38101 2896 38106 2952
rect 38162 2896 40000 2952
rect 38101 2894 40000 2896
rect 38101 2891 38167 2894
rect 39200 2864 40000 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 38101 1594 38167 1597
rect 39200 1594 40000 1624
rect 38101 1592 40000 1594
rect 38101 1536 38106 1592
rect 38162 1536 40000 1592
rect 38101 1534 40000 1536
rect 38101 1531 38167 1534
rect 39200 1504 40000 1534
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 20116 36212 20180 36276
rect 5580 36000 5644 36004
rect 5580 35944 5594 36000
rect 5594 35944 5644 36000
rect 5580 35940 5644 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 22508 35124 22572 35188
rect 25268 34988 25332 35052
rect 30972 35048 31036 35052
rect 30972 34992 30986 35048
rect 30986 34992 31036 35048
rect 30972 34988 31036 34992
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 30052 33824 30116 33828
rect 30052 33768 30102 33824
rect 30102 33768 30116 33824
rect 30052 33764 30116 33768
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 28396 33492 28460 33556
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19380 32736 19444 32740
rect 19380 32680 19430 32736
rect 19430 32680 19444 32736
rect 19380 32676 19444 32680
rect 22876 32676 22940 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 16436 32404 16500 32468
rect 27844 32404 27908 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 20116 31996 20180 32060
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 19380 31316 19444 31380
rect 30788 31240 30852 31244
rect 30788 31184 30802 31240
rect 30802 31184 30852 31240
rect 30788 31180 30852 31184
rect 31156 31044 31220 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 28580 30772 28644 30836
rect 23060 30500 23124 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 17540 30364 17604 30428
rect 30236 30092 30300 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 31524 29472 31588 29476
rect 31524 29416 31538 29472
rect 31538 29416 31588 29472
rect 31524 29412 31588 29416
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 29868 29004 29932 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 22876 28596 22940 28660
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 26004 27644 26068 27708
rect 27844 27508 27908 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 31524 26420 31588 26484
rect 28396 26284 28460 26348
rect 16436 26208 16500 26212
rect 16436 26152 16486 26208
rect 16486 26152 16500 26208
rect 16436 26148 16500 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 31156 25740 31220 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 26372 24924 26436 24988
rect 27476 24984 27540 24988
rect 27476 24928 27526 24984
rect 27526 24928 27540 24984
rect 27476 24924 27540 24928
rect 28764 24924 28828 24988
rect 17540 24788 17604 24852
rect 28212 24848 28276 24852
rect 28212 24792 28226 24848
rect 28226 24792 28276 24848
rect 28212 24788 28276 24792
rect 21220 24516 21284 24580
rect 23244 24516 23308 24580
rect 28580 24516 28644 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 30052 23700 30116 23764
rect 23428 23488 23492 23492
rect 23428 23432 23478 23488
rect 23478 23432 23492 23488
rect 23428 23428 23492 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 28028 23352 28092 23356
rect 28028 23296 28042 23352
rect 28042 23296 28092 23352
rect 28028 23292 28092 23296
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 30052 22808 30116 22812
rect 30052 22752 30066 22808
rect 30066 22752 30116 22808
rect 30052 22748 30116 22752
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 22508 21932 22572 21996
rect 25268 21992 25332 21996
rect 25268 21936 25282 21992
rect 25282 21936 25332 21992
rect 25268 21932 25332 21936
rect 29868 21932 29932 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 30972 20980 31036 21044
rect 28580 20768 28644 20772
rect 28580 20712 28594 20768
rect 28594 20712 28644 20768
rect 28580 20708 28644 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 23428 20632 23492 20636
rect 23428 20576 23442 20632
rect 23442 20576 23492 20632
rect 23428 20572 23492 20576
rect 5580 20436 5644 20500
rect 29132 20360 29196 20364
rect 29132 20304 29146 20360
rect 29146 20304 29196 20360
rect 29132 20300 29196 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 29132 19544 29196 19548
rect 29132 19488 29146 19544
rect 29146 19488 29196 19544
rect 29132 19484 29196 19488
rect 30788 19076 30852 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 30236 18668 30300 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 22140 18184 22204 18188
rect 22140 18128 22154 18184
rect 22154 18128 22204 18184
rect 22140 18124 22204 18128
rect 23244 18124 23308 18188
rect 34468 18124 34532 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 30236 16688 30300 16692
rect 30236 16632 30286 16688
rect 30286 16632 30300 16688
rect 30236 16628 30300 16632
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 26372 16220 26436 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 23060 15404 23124 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 26004 15192 26068 15196
rect 26004 15136 26054 15192
rect 26054 15136 26068 15192
rect 26004 15132 26068 15136
rect 28212 15132 28276 15196
rect 28764 15132 28828 15196
rect 28396 15056 28460 15060
rect 28396 15000 28410 15056
rect 28410 15000 28460 15056
rect 28396 14996 28460 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 34468 13908 34532 13972
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 27476 12276 27540 12340
rect 22140 12004 22204 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 21220 11324 21284 11388
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 28580 10100 28644 10164
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 22140 6216 22204 6220
rect 22140 6160 22154 6216
rect 22154 6160 22204 6216
rect 22140 6156 22204 6160
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 30236 3980 30300 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 5579 36004 5645 36005
rect 5579 35940 5580 36004
rect 5644 35940 5645 36004
rect 5579 35939 5645 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 5582 20501 5642 35939
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 20115 36276 20181 36277
rect 20115 36212 20116 36276
rect 20180 36212 20181 36276
rect 20115 36211 20181 36212
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19379 32740 19445 32741
rect 19379 32676 19380 32740
rect 19444 32676 19445 32740
rect 19379 32675 19445 32676
rect 16435 32468 16501 32469
rect 16435 32404 16436 32468
rect 16500 32404 16501 32468
rect 16435 32403 16501 32404
rect 16438 26213 16498 32403
rect 19382 31381 19442 32675
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 20118 32061 20178 36211
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 22507 35188 22573 35189
rect 22507 35124 22508 35188
rect 22572 35124 22573 35188
rect 22507 35123 22573 35124
rect 20115 32060 20181 32061
rect 20115 31996 20116 32060
rect 20180 31996 20181 32060
rect 20115 31995 20181 31996
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19379 31380 19445 31381
rect 19379 31316 19380 31380
rect 19444 31316 19445 31380
rect 19379 31315 19445 31316
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 17539 30428 17605 30429
rect 17539 30364 17540 30428
rect 17604 30364 17605 30428
rect 17539 30363 17605 30364
rect 16435 26212 16501 26213
rect 16435 26148 16436 26212
rect 16500 26148 16501 26212
rect 16435 26147 16501 26148
rect 17542 24853 17602 30363
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 17539 24852 17605 24853
rect 17539 24788 17540 24852
rect 17604 24788 17605 24852
rect 17539 24787 17605 24788
rect 19568 23968 19888 24992
rect 21219 24580 21285 24581
rect 21219 24516 21220 24580
rect 21284 24516 21285 24580
rect 21219 24515 21285 24516
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 5579 20500 5645 20501
rect 5579 20436 5580 20500
rect 5644 20436 5645 20500
rect 5579 20435 5645 20436
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 21222 11389 21282 24515
rect 22510 21997 22570 35123
rect 25267 35052 25333 35053
rect 25267 34988 25268 35052
rect 25332 34988 25333 35052
rect 25267 34987 25333 34988
rect 30971 35052 31037 35053
rect 30971 34988 30972 35052
rect 31036 34988 31037 35052
rect 30971 34987 31037 34988
rect 22875 32740 22941 32741
rect 22875 32676 22876 32740
rect 22940 32676 22941 32740
rect 22875 32675 22941 32676
rect 22878 28661 22938 32675
rect 23059 30564 23125 30565
rect 23059 30500 23060 30564
rect 23124 30500 23125 30564
rect 23059 30499 23125 30500
rect 22875 28660 22941 28661
rect 22875 28596 22876 28660
rect 22940 28596 22941 28660
rect 22875 28595 22941 28596
rect 22507 21996 22573 21997
rect 22507 21932 22508 21996
rect 22572 21932 22573 21996
rect 22507 21931 22573 21932
rect 22139 18188 22205 18189
rect 22139 18124 22140 18188
rect 22204 18124 22205 18188
rect 22139 18123 22205 18124
rect 22142 12069 22202 18123
rect 23062 15469 23122 30499
rect 23243 24580 23309 24581
rect 23243 24516 23244 24580
rect 23308 24516 23309 24580
rect 23243 24515 23309 24516
rect 23246 18189 23306 24515
rect 23427 23492 23493 23493
rect 23427 23428 23428 23492
rect 23492 23428 23493 23492
rect 23427 23427 23493 23428
rect 23430 20637 23490 23427
rect 25270 21997 25330 34987
rect 30051 33828 30117 33829
rect 30051 33764 30052 33828
rect 30116 33764 30117 33828
rect 30051 33763 30117 33764
rect 28395 33556 28461 33557
rect 28395 33492 28396 33556
rect 28460 33492 28461 33556
rect 28395 33491 28461 33492
rect 27843 32468 27909 32469
rect 27843 32404 27844 32468
rect 27908 32404 27909 32468
rect 27843 32403 27909 32404
rect 26003 27708 26069 27709
rect 26003 27644 26004 27708
rect 26068 27644 26069 27708
rect 26003 27643 26069 27644
rect 25267 21996 25333 21997
rect 25267 21932 25268 21996
rect 25332 21932 25333 21996
rect 25267 21931 25333 21932
rect 23427 20636 23493 20637
rect 23427 20572 23428 20636
rect 23492 20572 23493 20636
rect 23427 20571 23493 20572
rect 23243 18188 23309 18189
rect 23243 18124 23244 18188
rect 23308 18124 23309 18188
rect 23243 18123 23309 18124
rect 23059 15468 23125 15469
rect 23059 15404 23060 15468
rect 23124 15404 23125 15468
rect 23059 15403 23125 15404
rect 26006 15197 26066 27643
rect 27846 27573 27906 32403
rect 28398 31770 28458 33491
rect 28030 31710 28458 31770
rect 27843 27572 27909 27573
rect 27843 27508 27844 27572
rect 27908 27508 27909 27572
rect 27843 27507 27909 27508
rect 26371 24988 26437 24989
rect 26371 24924 26372 24988
rect 26436 24924 26437 24988
rect 26371 24923 26437 24924
rect 27475 24988 27541 24989
rect 27475 24924 27476 24988
rect 27540 24924 27541 24988
rect 27475 24923 27541 24924
rect 26374 16285 26434 24923
rect 26371 16284 26437 16285
rect 26371 16220 26372 16284
rect 26436 16220 26437 16284
rect 26371 16219 26437 16220
rect 26003 15196 26069 15197
rect 26003 15132 26004 15196
rect 26068 15132 26069 15196
rect 26003 15131 26069 15132
rect 27478 12341 27538 24923
rect 28030 23357 28090 31710
rect 28579 30836 28645 30837
rect 28579 30772 28580 30836
rect 28644 30772 28645 30836
rect 28579 30771 28645 30772
rect 28395 26348 28461 26349
rect 28395 26284 28396 26348
rect 28460 26284 28461 26348
rect 28395 26283 28461 26284
rect 28211 24852 28277 24853
rect 28211 24788 28212 24852
rect 28276 24788 28277 24852
rect 28211 24787 28277 24788
rect 28027 23356 28093 23357
rect 28027 23292 28028 23356
rect 28092 23292 28093 23356
rect 28027 23291 28093 23292
rect 28214 15197 28274 24787
rect 28211 15196 28277 15197
rect 28211 15132 28212 15196
rect 28276 15132 28277 15196
rect 28211 15131 28277 15132
rect 28398 15061 28458 26283
rect 28582 24581 28642 30771
rect 29867 29068 29933 29069
rect 29867 29004 29868 29068
rect 29932 29004 29933 29068
rect 29867 29003 29933 29004
rect 28763 24988 28829 24989
rect 28763 24924 28764 24988
rect 28828 24924 28829 24988
rect 28763 24923 28829 24924
rect 28579 24580 28645 24581
rect 28579 24516 28580 24580
rect 28644 24516 28645 24580
rect 28579 24515 28645 24516
rect 28579 20772 28645 20773
rect 28579 20708 28580 20772
rect 28644 20708 28645 20772
rect 28579 20707 28645 20708
rect 28395 15060 28461 15061
rect 28395 14996 28396 15060
rect 28460 14996 28461 15060
rect 28395 14995 28461 14996
rect 27475 12340 27541 12341
rect 27475 12276 27476 12340
rect 27540 12276 27541 12340
rect 27475 12275 27541 12276
rect 22139 12068 22205 12069
rect 22139 12004 22140 12068
rect 22204 12004 22205 12068
rect 22139 12003 22205 12004
rect 21219 11388 21285 11389
rect 21219 11324 21220 11388
rect 21284 11324 21285 11388
rect 21219 11323 21285 11324
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 22142 6221 22202 12003
rect 28582 10165 28642 20707
rect 28766 15197 28826 24923
rect 29870 21997 29930 29003
rect 30054 23765 30114 33763
rect 30787 31244 30853 31245
rect 30787 31180 30788 31244
rect 30852 31180 30853 31244
rect 30787 31179 30853 31180
rect 30235 30156 30301 30157
rect 30235 30092 30236 30156
rect 30300 30092 30301 30156
rect 30235 30091 30301 30092
rect 30051 23764 30117 23765
rect 30051 23700 30052 23764
rect 30116 23700 30117 23764
rect 30051 23699 30117 23700
rect 30054 22813 30114 23699
rect 30051 22812 30117 22813
rect 30051 22748 30052 22812
rect 30116 22748 30117 22812
rect 30051 22747 30117 22748
rect 29867 21996 29933 21997
rect 29867 21932 29868 21996
rect 29932 21932 29933 21996
rect 29867 21931 29933 21932
rect 29131 20364 29197 20365
rect 29131 20300 29132 20364
rect 29196 20300 29197 20364
rect 29131 20299 29197 20300
rect 29134 19549 29194 20299
rect 29131 19548 29197 19549
rect 29131 19484 29132 19548
rect 29196 19484 29197 19548
rect 29131 19483 29197 19484
rect 30238 18733 30298 30091
rect 30790 19141 30850 31179
rect 30974 21045 31034 34987
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 31155 31108 31221 31109
rect 31155 31044 31156 31108
rect 31220 31044 31221 31108
rect 31155 31043 31221 31044
rect 31158 25805 31218 31043
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 31523 29476 31589 29477
rect 31523 29412 31524 29476
rect 31588 29412 31589 29476
rect 31523 29411 31589 29412
rect 31526 26485 31586 29411
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 31523 26484 31589 26485
rect 31523 26420 31524 26484
rect 31588 26420 31589 26484
rect 31523 26419 31589 26420
rect 31155 25804 31221 25805
rect 31155 25740 31156 25804
rect 31220 25740 31221 25804
rect 31155 25739 31221 25740
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 30971 21044 31037 21045
rect 30971 20980 30972 21044
rect 31036 20980 31037 21044
rect 30971 20979 31037 20980
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 30787 19140 30853 19141
rect 30787 19076 30788 19140
rect 30852 19076 30853 19140
rect 30787 19075 30853 19076
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 30235 18732 30301 18733
rect 30235 18668 30236 18732
rect 30300 18668 30301 18732
rect 30235 18667 30301 18668
rect 34467 18188 34533 18189
rect 34467 18124 34468 18188
rect 34532 18124 34533 18188
rect 34467 18123 34533 18124
rect 30235 16692 30301 16693
rect 30235 16628 30236 16692
rect 30300 16628 30301 16692
rect 30235 16627 30301 16628
rect 28763 15196 28829 15197
rect 28763 15132 28764 15196
rect 28828 15132 28829 15196
rect 28763 15131 28829 15132
rect 28579 10164 28645 10165
rect 28579 10100 28580 10164
rect 28644 10100 28645 10164
rect 28579 10099 28645 10100
rect 22139 6220 22205 6221
rect 22139 6156 22140 6220
rect 22204 6156 22205 6220
rect 22139 6155 22205 6156
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 30238 4045 30298 16627
rect 34470 13973 34530 18123
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34467 13972 34533 13973
rect 34467 13908 34468 13972
rect 34532 13908 34533 13972
rect 34467 13907 34533 13908
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 30235 4044 30301 4045
rect 30235 3980 30236 4044
rect 30300 3980 30301 4044
rect 30235 3979 30301 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_267
timestamp 1676037725
transform 1 0 25668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1676037725
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_303
timestamp 1676037725
transform 1 0 28980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_324
timestamp 1676037725
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_360
timestamp 1676037725
transform 1 0 34224 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_372
timestamp 1676037725
transform 1 0 35328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_161
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_183
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1676037725
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1676037725
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1676037725
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1676037725
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_327
timestamp 1676037725
transform 1 0 31188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_339
timestamp 1676037725
transform 1 0 32292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1676037725
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_373
timestamp 1676037725
transform 1 0 35420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_383
timestamp 1676037725
transform 1 0 36340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_387
timestamp 1676037725
transform 1 0 36708 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1676037725
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1676037725
transform 1 0 23644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp 1676037725
transform 1 0 24380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_263
timestamp 1676037725
transform 1 0 25300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1676037725
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1676037725
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_355
timestamp 1676037725
transform 1 0 33764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_364
timestamp 1676037725
transform 1 0 34592 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_368
timestamp 1676037725
transform 1 0 34960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_404
timestamp 1676037725
transform 1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1676037725
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_232
timestamp 1676037725
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1676037725
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_261
timestamp 1676037725
transform 1 0 25116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_266
timestamp 1676037725
transform 1 0 25576 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_278
timestamp 1676037725
transform 1 0 26680 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_290
timestamp 1676037725
transform 1 0 27784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_300
timestamp 1676037725
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_315
timestamp 1676037725
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_332
timestamp 1676037725
transform 1 0 31648 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_340
timestamp 1676037725
transform 1 0 32384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_351
timestamp 1676037725
transform 1 0 33396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1676037725
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_375
timestamp 1676037725
transform 1 0 35604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_387
timestamp 1676037725
transform 1 0 36708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1676037725
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_177
timestamp 1676037725
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1676037725
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1676037725
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_230
timestamp 1676037725
transform 1 0 22264 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_238
timestamp 1676037725
transform 1 0 23000 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_265
timestamp 1676037725
transform 1 0 25484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1676037725
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1676037725
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1676037725
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_327
timestamp 1676037725
transform 1 0 31188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_362
timestamp 1676037725
transform 1 0 34408 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_374
timestamp 1676037725
transform 1 0 35512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1676037725
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_404
timestamp 1676037725
transform 1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_169
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1676037725
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_224
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1676037725
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_264
timestamp 1676037725
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_288
timestamp 1676037725
transform 1 0 27600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp 1676037725
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_323
timestamp 1676037725
transform 1 0 30820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_335
timestamp 1676037725
transform 1 0 31924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_347
timestamp 1676037725
transform 1 0 33028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_385
timestamp 1676037725
transform 1 0 36524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1676037725
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_122
timestamp 1676037725
transform 1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_130
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_150
timestamp 1676037725
transform 1 0 14904 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1676037725
transform 1 0 15272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1676037725
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_198
timestamp 1676037725
transform 1 0 19320 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_212
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_230
timestamp 1676037725
transform 1 0 22264 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_242
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_292
timestamp 1676037725
transform 1 0 27968 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_304
timestamp 1676037725
transform 1 0 29072 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_316
timestamp 1676037725
transform 1 0 30176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1676037725
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_359
timestamp 1676037725
transform 1 0 34132 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_162
timestamp 1676037725
transform 1 0 16008 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1676037725
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_238
timestamp 1676037725
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1676037725
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1676037725
transform 1 0 25668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1676037725
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_300
timestamp 1676037725
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_318
timestamp 1676037725
transform 1 0 30360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_322
timestamp 1676037725
transform 1 0 30728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_339
timestamp 1676037725
transform 1 0 32292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_352
timestamp 1676037725
transform 1 0 33488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1676037725
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_380
timestamp 1676037725
transform 1 0 36064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_388
timestamp 1676037725
transform 1 0 36800 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1676037725
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_128
timestamp 1676037725
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_136
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_146
timestamp 1676037725
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1676037725
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_194
timestamp 1676037725
transform 1 0 18952 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_200
timestamp 1676037725
transform 1 0 19504 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1676037725
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_268
timestamp 1676037725
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_296
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_309
timestamp 1676037725
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_356
timestamp 1676037725
transform 1 0 33856 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1676037725
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_149
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_180
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_206
timestamp 1676037725
transform 1 0 20056 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_212
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_222
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_234
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1676037725
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1676037725
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_264
timestamp 1676037725
transform 1 0 25392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_279
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_294
timestamp 1676037725
transform 1 0 28152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_320
timestamp 1676037725
transform 1 0 30544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_340
timestamp 1676037725
transform 1 0 32384 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_373
timestamp 1676037725
transform 1 0 35420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1676037725
transform 1 0 37444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1676037725
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1676037725
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1676037725
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_174
timestamp 1676037725
transform 1 0 17112 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_186
timestamp 1676037725
transform 1 0 18216 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_262
timestamp 1676037725
transform 1 0 25208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_270
timestamp 1676037725
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_299
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_322
timestamp 1676037725
transform 1 0 30728 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_348
timestamp 1676037725
transform 1 0 33120 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_370
timestamp 1676037725
transform 1 0 35144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1676037725
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1676037725
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_220
timestamp 1676037725
transform 1 0 21344 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_227
timestamp 1676037725
transform 1 0 21988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_239
timestamp 1676037725
transform 1 0 23092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_266
timestamp 1676037725
transform 1 0 25576 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_278
timestamp 1676037725
transform 1 0 26680 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_290
timestamp 1676037725
transform 1 0 27784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_302
timestamp 1676037725
transform 1 0 28888 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1676037725
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_390
timestamp 1676037725
transform 1 0 36984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_398
timestamp 1676037725
transform 1 0 37720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1676037725
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_151
timestamp 1676037725
transform 1 0 14996 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_206
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_212
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_246
timestamp 1676037725
transform 1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_252
timestamp 1676037725
transform 1 0 24288 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_324
timestamp 1676037725
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_364
timestamp 1676037725
transform 1 0 34592 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1676037725
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_404
timestamp 1676037725
transform 1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_106
timestamp 1676037725
transform 1 0 10856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_114
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1676037725
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1676037725
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_185
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1676037725
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_212
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_220
timestamp 1676037725
transform 1 0 21344 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_270
timestamp 1676037725
transform 1 0 25944 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_292
timestamp 1676037725
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_296
timestamp 1676037725
transform 1 0 28336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_332
timestamp 1676037725
transform 1 0 31648 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1676037725
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1676037725
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_387
timestamp 1676037725
transform 1 0 36708 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_404
timestamp 1676037725
transform 1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_86
timestamp 1676037725
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_98
timestamp 1676037725
transform 1 0 10120 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_130
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1676037725
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1676037725
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_266
timestamp 1676037725
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1676037725
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_355
timestamp 1676037725
transform 1 0 33764 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_367
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1676037725
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1676037725
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1676037725
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1676037725
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_228
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_261
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_284
timestamp 1676037725
transform 1 0 27232 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_290
timestamp 1676037725
transform 1 0 27784 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1676037725
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_331
timestamp 1676037725
transform 1 0 31556 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_348
timestamp 1676037725
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1676037725
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_378
timestamp 1676037725
transform 1 0 35880 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_386
timestamp 1676037725
transform 1 0 36616 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1676037725
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_65
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1676037725
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_136
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1676037725
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_241
timestamp 1676037725
transform 1 0 23276 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_246
timestamp 1676037725
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_262
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_300
timestamp 1676037725
transform 1 0 28704 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_312
timestamp 1676037725
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_324
timestamp 1676037725
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_353
timestamp 1676037725
transform 1 0 33580 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_371
timestamp 1676037725
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_383
timestamp 1676037725
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1676037725
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_103
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_183
timestamp 1676037725
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_225
timestamp 1676037725
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_259
timestamp 1676037725
transform 1 0 24932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1676037725
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_329
timestamp 1676037725
transform 1 0 31372 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_341
timestamp 1676037725
transform 1 0 32476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_348
timestamp 1676037725
transform 1 0 33120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_355
timestamp 1676037725
transform 1 0 33764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_373
timestamp 1676037725
transform 1 0 35420 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_393
timestamp 1676037725
transform 1 0 37260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1676037725
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_89
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1676037725
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_185
timestamp 1676037725
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1676037725
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1676037725
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_304
timestamp 1676037725
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_321
timestamp 1676037725
transform 1 0 30636 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_345
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_354
timestamp 1676037725
transform 1 0 33672 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_366
timestamp 1676037725
transform 1 0 34776 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_378
timestamp 1676037725
transform 1 0 35880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 1676037725
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_149
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_157
timestamp 1676037725
transform 1 0 15548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_169
timestamp 1676037725
transform 1 0 16652 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_184
timestamp 1676037725
transform 1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_190
timestamp 1676037725
transform 1 0 18584 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_210
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1676037725
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_228
timestamp 1676037725
transform 1 0 22080 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1676037725
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_263
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_275
timestamp 1676037725
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_281
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_285
timestamp 1676037725
transform 1 0 27324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1676037725
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_341
timestamp 1676037725
transform 1 0 32476 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_349
timestamp 1676037725
transform 1 0 33212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1676037725
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_381
timestamp 1676037725
transform 1 0 36156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1676037725
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1676037725
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_100
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_140
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1676037725
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_203
timestamp 1676037725
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_254
timestamp 1676037725
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_262
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1676037725
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1676037725
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_300
timestamp 1676037725
transform 1 0 28704 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_312
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_357
timestamp 1676037725
transform 1 0 33948 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_363
timestamp 1676037725
transform 1 0 34500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_381
timestamp 1676037725
transform 1 0 36156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1676037725
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1676037725
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_107
timestamp 1676037725
transform 1 0 10948 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_120
timestamp 1676037725
transform 1 0 12144 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_212
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1676037725
transform 1 0 22816 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 1676037725
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_273
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_281
timestamp 1676037725
transform 1 0 26956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_285
timestamp 1676037725
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_334
timestamp 1676037725
transform 1 0 31832 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_346
timestamp 1676037725
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1676037725
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_376
timestamp 1676037725
transform 1 0 35696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_388
timestamp 1676037725
transform 1 0 36800 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1676037725
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1676037725
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_87
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_201
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_239
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_271
timestamp 1676037725
transform 1 0 26036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_291
timestamp 1676037725
transform 1 0 27876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_299
timestamp 1676037725
transform 1 0 28612 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_308
timestamp 1676037725
transform 1 0 29440 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1676037725
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_346
timestamp 1676037725
transform 1 0 32936 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_357
timestamp 1676037725
transform 1 0 33948 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_369
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_378
timestamp 1676037725
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_404
timestamp 1676037725
transform 1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1676037725
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1676037725
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1676037725
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_176
timestamp 1676037725
transform 1 0 17296 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1676037725
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_217
timestamp 1676037725
transform 1 0 21068 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_235
timestamp 1676037725
transform 1 0 22724 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1676037725
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_279
timestamp 1676037725
transform 1 0 26772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_290
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_319
timestamp 1676037725
transform 1 0 30452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_323
timestamp 1676037725
transform 1 0 30820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_331
timestamp 1676037725
transform 1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_335
timestamp 1676037725
transform 1 0 31924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_344
timestamp 1676037725
transform 1 0 32752 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_375
timestamp 1676037725
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1676037725
transform 1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1676037725
transform 1 0 8188 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_122
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_142
timestamp 1676037725
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1676037725
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1676037725
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_208
timestamp 1676037725
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1676037725
transform 1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_304
timestamp 1676037725
transform 1 0 29072 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_318
timestamp 1676037725
transform 1 0 30360 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_326
timestamp 1676037725
transform 1 0 31096 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_359
timestamp 1676037725
transform 1 0 34132 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1676037725
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_371
timestamp 1676037725
transform 1 0 35236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1676037725
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1676037725
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_130
timestamp 1676037725
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_178
timestamp 1676037725
transform 1 0 17480 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1676037725
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_229
timestamp 1676037725
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_262
timestamp 1676037725
transform 1 0 25208 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_270
timestamp 1676037725
transform 1 0 25944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_290
timestamp 1676037725
transform 1 0 27784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_298
timestamp 1676037725
transform 1 0 28520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1676037725
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_328
timestamp 1676037725
transform 1 0 31280 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_339
timestamp 1676037725
transform 1 0 32292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_351
timestamp 1676037725
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_385
timestamp 1676037725
transform 1 0 36524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1676037725
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_77
timestamp 1676037725
transform 1 0 8188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_182
timestamp 1676037725
transform 1 0 17848 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1676037725
transform 1 0 20608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_233
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_267
timestamp 1676037725
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_289
timestamp 1676037725
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_297
timestamp 1676037725
transform 1 0 28428 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_314
timestamp 1676037725
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_354
timestamp 1676037725
transform 1 0 33672 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_366
timestamp 1676037725
transform 1 0 34776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_376
timestamp 1676037725
transform 1 0 35696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1676037725
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_35
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_52
timestamp 1676037725
transform 1 0 5888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1676037725
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_94
timestamp 1676037725
transform 1 0 9752 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1676037725
transform 1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1676037725
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_159
timestamp 1676037725
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_171
timestamp 1676037725
transform 1 0 16836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_218
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_234
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_260
timestamp 1676037725
transform 1 0 25024 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_279
timestamp 1676037725
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_291
timestamp 1676037725
transform 1 0 27876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1676037725
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1676037725
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1676037725
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_400
timestamp 1676037725
transform 1 0 37904 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1676037725
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_65
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_77
timestamp 1676037725
transform 1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_94
timestamp 1676037725
transform 1 0 9752 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1676037725
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_131
timestamp 1676037725
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1676037725
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1676037725
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1676037725
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_247
timestamp 1676037725
transform 1 0 23828 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_292
timestamp 1676037725
transform 1 0 27968 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1676037725
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_302
timestamp 1676037725
transform 1 0 28888 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_314
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1676037725
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_345
timestamp 1676037725
transform 1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_353
timestamp 1676037725
transform 1 0 33580 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_378
timestamp 1676037725
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1676037725
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp 1676037725
transform 1 0 7912 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_103
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_116
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_128
timestamp 1676037725
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_171
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_262
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_270
timestamp 1676037725
transform 1 0 25944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_280
timestamp 1676037725
transform 1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 1676037725
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_317
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_332
timestamp 1676037725
transform 1 0 31648 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_338
timestamp 1676037725
transform 1 0 32200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_347
timestamp 1676037725
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1676037725
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_375
timestamp 1676037725
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1676037725
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_87
timestamp 1676037725
transform 1 0 9108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1676037725
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_190
timestamp 1676037725
transform 1 0 18584 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_248
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_254
timestamp 1676037725
transform 1 0 24472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_268
timestamp 1676037725
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_290
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_302
timestamp 1676037725
transform 1 0 28888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_312
timestamp 1676037725
transform 1 0 29808 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_320
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_345
timestamp 1676037725
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_353
timestamp 1676037725
transform 1 0 33580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_365
timestamp 1676037725
transform 1 0 34684 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_378
timestamp 1676037725
transform 1 0 35880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_404
timestamp 1676037725
transform 1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 1676037725
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_54
timestamp 1676037725
transform 1 0 6072 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_66
timestamp 1676037725
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1676037725
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_107
timestamp 1676037725
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_127
timestamp 1676037725
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_172
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1676037725
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_261
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_284
timestamp 1676037725
transform 1 0 27232 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1676037725
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_325
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_335
timestamp 1676037725
transform 1 0 31924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_347
timestamp 1676037725
transform 1 0 33028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1676037725
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_381
timestamp 1676037725
transform 1 0 36156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_393
timestamp 1676037725
transform 1 0 37260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1676037725
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_38
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_46
timestamp 1676037725
transform 1 0 5336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_66
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_72
timestamp 1676037725
transform 1 0 7728 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_80
timestamp 1676037725
transform 1 0 8464 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_89
timestamp 1676037725
transform 1 0 9292 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_156
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_195
timestamp 1676037725
transform 1 0 19044 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_207
timestamp 1676037725
transform 1 0 20148 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_243
timestamp 1676037725
transform 1 0 23460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_251
timestamp 1676037725
transform 1 0 24196 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1676037725
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_286
timestamp 1676037725
transform 1 0 27416 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_294
timestamp 1676037725
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1676037725
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_346
timestamp 1676037725
transform 1 0 32936 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_383
timestamp 1676037725
transform 1 0 36340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_404
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_40
timestamp 1676037725
transform 1 0 4784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1676037725
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1676037725
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_108
timestamp 1676037725
transform 1 0 11040 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_120
timestamp 1676037725
transform 1 0 12144 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1676037725
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_156
timestamp 1676037725
transform 1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_175
timestamp 1676037725
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1676037725
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_270
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_278
timestamp 1676037725
transform 1 0 26680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_286
timestamp 1676037725
transform 1 0 27416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_293
timestamp 1676037725
transform 1 0 28060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_297
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_339
timestamp 1676037725
transform 1 0 32292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_348
timestamp 1676037725
transform 1 0 33120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1676037725
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_373
timestamp 1676037725
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_381
timestamp 1676037725
transform 1 0 36156 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_387
timestamp 1676037725
transform 1 0 36708 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_404
timestamp 1676037725
transform 1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_73
timestamp 1676037725
transform 1 0 7820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_77
timestamp 1676037725
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_85
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_97
timestamp 1676037725
transform 1 0 10028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1676037725
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_131
timestamp 1676037725
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_152
timestamp 1676037725
transform 1 0 15088 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_185
timestamp 1676037725
transform 1 0 18124 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_212
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_235
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_247
timestamp 1676037725
transform 1 0 23828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_253
timestamp 1676037725
transform 1 0 24380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_257
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1676037725
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_297
timestamp 1676037725
transform 1 0 28428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_309
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_354
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_366
timestamp 1676037725
transform 1 0 34776 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1676037725
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_40
timestamp 1676037725
transform 1 0 4784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_50
timestamp 1676037725
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_63
timestamp 1676037725
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1676037725
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_105
timestamp 1676037725
transform 1 0 10764 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_125
timestamp 1676037725
transform 1 0 12604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1676037725
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1676037725
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_154
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_161
timestamp 1676037725
transform 1 0 15916 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_167
timestamp 1676037725
transform 1 0 16468 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1676037725
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_234
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1676037725
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_266
timestamp 1676037725
transform 1 0 25576 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_272
timestamp 1676037725
transform 1 0 26128 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_288
timestamp 1676037725
transform 1 0 27600 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1676037725
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_324
timestamp 1676037725
transform 1 0 30912 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_336
timestamp 1676037725
transform 1 0 32016 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_348
timestamp 1676037725
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1676037725
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_379
timestamp 1676037725
transform 1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_387
timestamp 1676037725
transform 1 0 36708 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_404
timestamp 1676037725
transform 1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_45
timestamp 1676037725
transform 1 0 5244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1676037725
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_66
timestamp 1676037725
transform 1 0 7176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_78
timestamp 1676037725
transform 1 0 8280 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_96
timestamp 1676037725
transform 1 0 9936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1676037725
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_142
timestamp 1676037725
transform 1 0 14168 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_178
timestamp 1676037725
transform 1 0 17480 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_190
timestamp 1676037725
transform 1 0 18584 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1676037725
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1676037725
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_252
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1676037725
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_304
timestamp 1676037725
transform 1 0 29072 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_351
timestamp 1676037725
transform 1 0 33396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_359
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_375
timestamp 1676037725
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1676037725
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 1676037725
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_56
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_66
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_70
timestamp 1676037725
transform 1 0 7544 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1676037725
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_94
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_102
timestamp 1676037725
transform 1 0 10488 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_119
timestamp 1676037725
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1676037725
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_173
timestamp 1676037725
transform 1 0 17020 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1676037725
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_204
timestamp 1676037725
transform 1 0 19872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1676037725
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_228
timestamp 1676037725
transform 1 0 22080 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_242
timestamp 1676037725
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_272
timestamp 1676037725
transform 1 0 26128 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1676037725
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_290
timestamp 1676037725
transform 1 0 27784 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1676037725
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_335
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_346
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_354
timestamp 1676037725
transform 1 0 33672 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1676037725
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_372
timestamp 1676037725
transform 1 0 35328 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_384
timestamp 1676037725
transform 1 0 36432 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_396
timestamp 1676037725
transform 1 0 37536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_34
timestamp 1676037725
transform 1 0 4232 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1676037725
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1676037725
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_66
timestamp 1676037725
transform 1 0 7176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_78
timestamp 1676037725
transform 1 0 8280 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_84
timestamp 1676037725
transform 1 0 8832 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1676037725
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1676037725
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1676037725
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1676037725
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1676037725
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_199
timestamp 1676037725
transform 1 0 19412 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1676037725
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1676037725
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1676037725
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1676037725
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_294
timestamp 1676037725
transform 1 0 28152 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_304
timestamp 1676037725
transform 1 0 29072 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_311
timestamp 1676037725
transform 1 0 29716 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1676037725
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_360
timestamp 1676037725
transform 1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_364
timestamp 1676037725
transform 1 0 34592 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_382
timestamp 1676037725
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1676037725
transform 1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_37
timestamp 1676037725
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_49
timestamp 1676037725
transform 1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_57
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_66
timestamp 1676037725
transform 1 0 7176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1676037725
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_95
timestamp 1676037725
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_107
timestamp 1676037725
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_119
timestamp 1676037725
transform 1 0 12052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_149
timestamp 1676037725
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_161
timestamp 1676037725
transform 1 0 15916 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_176
timestamp 1676037725
transform 1 0 17296 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_184
timestamp 1676037725
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_219
timestamp 1676037725
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_231
timestamp 1676037725
transform 1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1676037725
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_266
timestamp 1676037725
transform 1 0 25576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_281
timestamp 1676037725
transform 1 0 26956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_287
timestamp 1676037725
transform 1 0 27508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_295
timestamp 1676037725
transform 1 0 28244 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1676037725
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_319
timestamp 1676037725
transform 1 0 30452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_331
timestamp 1676037725
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_343
timestamp 1676037725
transform 1 0 32660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1676037725
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1676037725
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_379
timestamp 1676037725
transform 1 0 35972 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_385
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1676037725
transform 1 0 38088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1676037725
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_63
timestamp 1676037725
transform 1 0 6900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp 1676037725
transform 1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_82
timestamp 1676037725
transform 1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_90
timestamp 1676037725
transform 1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1676037725
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1676037725
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_132
timestamp 1676037725
transform 1 0 13248 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_138
timestamp 1676037725
transform 1 0 13800 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_145
timestamp 1676037725
transform 1 0 14444 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_157
timestamp 1676037725
transform 1 0 15548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1676037725
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_201
timestamp 1676037725
transform 1 0 19596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_234
timestamp 1676037725
transform 1 0 22632 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_245
timestamp 1676037725
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1676037725
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1676037725
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1676037725
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_294
timestamp 1676037725
transform 1 0 28152 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_300
timestamp 1676037725
transform 1 0 28704 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1676037725
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_364
timestamp 1676037725
transform 1 0 34592 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_387
timestamp 1676037725
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_48
timestamp 1676037725
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_55
timestamp 1676037725
transform 1 0 6164 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_67
timestamp 1676037725
transform 1 0 7268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_75
timestamp 1676037725
transform 1 0 8004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1676037725
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_92
timestamp 1676037725
transform 1 0 9568 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1676037725
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_124
timestamp 1676037725
transform 1 0 12512 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1676037725
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1676037725
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1676037725
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_161
timestamp 1676037725
transform 1 0 15916 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1676037725
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1676037725
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_204
timestamp 1676037725
transform 1 0 19872 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_210
timestamp 1676037725
transform 1 0 20424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_218
timestamp 1676037725
transform 1 0 21160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1676037725
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_239
timestamp 1676037725
transform 1 0 23092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_276
timestamp 1676037725
transform 1 0 26496 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_288
timestamp 1676037725
transform 1 0 27600 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_296
timestamp 1676037725
transform 1 0 28336 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_318
timestamp 1676037725
transform 1 0 30360 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_340
timestamp 1676037725
transform 1 0 32384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_353
timestamp 1676037725
transform 1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1676037725
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_375
timestamp 1676037725
transform 1 0 35604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_383
timestamp 1676037725
transform 1 0 36340 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_34
timestamp 1676037725
transform 1 0 4232 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_40
timestamp 1676037725
transform 1 0 4784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1676037725
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_63
timestamp 1676037725
transform 1 0 6900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_70
timestamp 1676037725
transform 1 0 7544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_91
timestamp 1676037725
transform 1 0 9476 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_102
timestamp 1676037725
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1676037725
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_134
timestamp 1676037725
transform 1 0 13432 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1676037725
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1676037725
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_198
timestamp 1676037725
transform 1 0 19320 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1676037725
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_213
timestamp 1676037725
transform 1 0 20700 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_243
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_247
timestamp 1676037725
transform 1 0 23828 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_251
timestamp 1676037725
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_263
timestamp 1676037725
transform 1 0 25300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_271
timestamp 1676037725
transform 1 0 26036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_299
timestamp 1676037725
transform 1 0 28612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_319
timestamp 1676037725
transform 1 0 30452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1676037725
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1676037725
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_353
timestamp 1676037725
transform 1 0 33580 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1676037725
transform 1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_377
timestamp 1676037725
transform 1 0 35788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1676037725
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_404
timestamp 1676037725
transform 1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_39
timestamp 1676037725
transform 1 0 4692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_52
timestamp 1676037725
transform 1 0 5888 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_60
timestamp 1676037725
transform 1 0 6624 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_68
timestamp 1676037725
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1676037725
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_90
timestamp 1676037725
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_98
timestamp 1676037725
transform 1 0 10120 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_105
timestamp 1676037725
transform 1 0 10764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1676037725
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_175
timestamp 1676037725
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_236
timestamp 1676037725
transform 1 0 22816 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_259
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_273
timestamp 1676037725
transform 1 0 26220 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1676037725
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_294
timestamp 1676037725
transform 1 0 28152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1676037725
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_320
timestamp 1676037725
transform 1 0 30544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_324
timestamp 1676037725
transform 1 0 30912 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_332
timestamp 1676037725
transform 1 0 31648 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_338
timestamp 1676037725
transform 1 0 32200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_348
timestamp 1676037725
transform 1 0 33120 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1676037725
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_373
timestamp 1676037725
transform 1 0 35420 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_385
timestamp 1676037725
transform 1 0 36524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1676037725
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1676037725
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1676037725
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_67
timestamp 1676037725
transform 1 0 7268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_79
timestamp 1676037725
transform 1 0 8372 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_87
timestamp 1676037725
transform 1 0 9108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_92
timestamp 1676037725
transform 1 0 9568 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_98
timestamp 1676037725
transform 1 0 10120 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_148
timestamp 1676037725
transform 1 0 14720 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_160
timestamp 1676037725
transform 1 0 15824 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_174
timestamp 1676037725
transform 1 0 17112 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_186
timestamp 1676037725
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_198
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_206
timestamp 1676037725
transform 1 0 20056 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_212
timestamp 1676037725
transform 1 0 20608 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1676037725
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1676037725
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_239
timestamp 1676037725
transform 1 0 23092 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_255
timestamp 1676037725
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_265
timestamp 1676037725
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1676037725
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_291
timestamp 1676037725
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_295
timestamp 1676037725
transform 1 0 28244 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_300
timestamp 1676037725
transform 1 0 28704 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_308
timestamp 1676037725
transform 1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_319
timestamp 1676037725
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1676037725
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_346
timestamp 1676037725
transform 1 0 32936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_358
timestamp 1676037725
transform 1 0 34040 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_376
timestamp 1676037725
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1676037725
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_404
timestamp 1676037725
transform 1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_40
timestamp 1676037725
transform 1 0 4784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_44
timestamp 1676037725
transform 1 0 5152 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_50
timestamp 1676037725
transform 1 0 5704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_58
timestamp 1676037725
transform 1 0 6440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_64
timestamp 1676037725
transform 1 0 6992 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_73
timestamp 1676037725
transform 1 0 7820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1676037725
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1676037725
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_107
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_113
timestamp 1676037725
transform 1 0 11500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_120
timestamp 1676037725
transform 1 0 12144 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_147
timestamp 1676037725
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_154
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_162
timestamp 1676037725
transform 1 0 16008 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_171
timestamp 1676037725
transform 1 0 16836 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_182
timestamp 1676037725
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_204
timestamp 1676037725
transform 1 0 19872 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_216
timestamp 1676037725
transform 1 0 20976 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_226
timestamp 1676037725
transform 1 0 21896 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_232
timestamp 1676037725
transform 1 0 22448 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_266
timestamp 1676037725
transform 1 0 25576 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_278
timestamp 1676037725
transform 1 0 26680 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_286
timestamp 1676037725
transform 1 0 27416 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_292
timestamp 1676037725
transform 1 0 27968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1676037725
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_317
timestamp 1676037725
transform 1 0 30268 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_328
timestamp 1676037725
transform 1 0 31280 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_341
timestamp 1676037725
transform 1 0 32476 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1676037725
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_373
timestamp 1676037725
transform 1 0 35420 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_382
timestamp 1676037725
transform 1 0 36248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_402
timestamp 1676037725
transform 1 0 38088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1676037725
transform 1 0 38456 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_31
timestamp 1676037725
transform 1 0 3956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_49
timestamp 1676037725
transform 1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_64
timestamp 1676037725
transform 1 0 6992 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_72
timestamp 1676037725
transform 1 0 7728 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1676037725
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_84
timestamp 1676037725
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_91
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_106
timestamp 1676037725
transform 1 0 10856 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1676037725
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_121
timestamp 1676037725
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_128
timestamp 1676037725
transform 1 0 12880 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_148
timestamp 1676037725
transform 1 0 14720 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1676037725
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1676037725
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1676037725
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_257
timestamp 1676037725
transform 1 0 24748 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_266
timestamp 1676037725
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1676037725
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_290
timestamp 1676037725
transform 1 0 27784 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_301
timestamp 1676037725
transform 1 0 28796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_311
timestamp 1676037725
transform 1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_324
timestamp 1676037725
transform 1 0 30912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_333
timestamp 1676037725
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_345
timestamp 1676037725
transform 1 0 32844 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_357
timestamp 1676037725
transform 1 0 33948 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_365
timestamp 1676037725
transform 1 0 34684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_374
timestamp 1676037725
transform 1 0 35512 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_382
timestamp 1676037725
transform 1 0 36248 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1676037725
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_401
timestamp 1676037725
transform 1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_19
timestamp 1676037725
transform 1 0 2852 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1676037725
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_40
timestamp 1676037725
transform 1 0 4784 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_54
timestamp 1676037725
transform 1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_62
timestamp 1676037725
transform 1 0 6808 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1676037725
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_107
timestamp 1676037725
transform 1 0 10948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_120
timestamp 1676037725
transform 1 0 12144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1676037725
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_154
timestamp 1676037725
transform 1 0 15272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_166
timestamp 1676037725
transform 1 0 16376 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1676037725
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_174
timestamp 1676037725
transform 1 0 17112 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_181
timestamp 1676037725
transform 1 0 17756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_205
timestamp 1676037725
transform 1 0 19964 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1676037725
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_225
timestamp 1676037725
transform 1 0 21804 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_237
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1676037725
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_274
timestamp 1676037725
transform 1 0 26312 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_280
timestamp 1676037725
transform 1 0 26864 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_290
timestamp 1676037725
transform 1 0 27784 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_296
timestamp 1676037725
transform 1 0 28336 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1676037725
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_319
timestamp 1676037725
transform 1 0 30452 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_341
timestamp 1676037725
transform 1 0 32476 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1676037725
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_374
timestamp 1676037725
transform 1 0 35512 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_384
timestamp 1676037725
transform 1 0 36432 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1676037725
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_35
timestamp 1676037725
transform 1 0 4324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_43
timestamp 1676037725
transform 1 0 5060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1676037725
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_74
timestamp 1676037725
transform 1 0 7912 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_78
timestamp 1676037725
transform 1 0 8280 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_84
timestamp 1676037725
transform 1 0 8832 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_96
timestamp 1676037725
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1676037725
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_120
timestamp 1676037725
transform 1 0 12144 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_128
timestamp 1676037725
transform 1 0 12880 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_133
timestamp 1676037725
transform 1 0 13340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_141
timestamp 1676037725
transform 1 0 14076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_148
timestamp 1676037725
transform 1 0 14720 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_158
timestamp 1676037725
transform 1 0 15640 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1676037725
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_183
timestamp 1676037725
transform 1 0 17940 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_190
timestamp 1676037725
transform 1 0 18584 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_202
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_210
timestamp 1676037725
transform 1 0 20424 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_233
timestamp 1676037725
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_243
timestamp 1676037725
transform 1 0 23460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1676037725
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_254
timestamp 1676037725
transform 1 0 24472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_260
timestamp 1676037725
transform 1 0 25024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1676037725
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_299
timestamp 1676037725
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_306
timestamp 1676037725
transform 1 0 29256 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_310
timestamp 1676037725
transform 1 0 29624 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_319
timestamp 1676037725
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1676037725
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_344
timestamp 1676037725
transform 1 0 32752 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_352
timestamp 1676037725
transform 1 0 33488 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_370
timestamp 1676037725
transform 1 0 35144 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_374
timestamp 1676037725
transform 1 0 35512 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1676037725
transform 1 0 36340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_46
timestamp 1676037725
transform 1 0 5336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_55
timestamp 1676037725
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1676037725
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_103
timestamp 1676037725
transform 1 0 10580 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_124
timestamp 1676037725
transform 1 0 12512 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_132
timestamp 1676037725
transform 1 0 13248 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_149
timestamp 1676037725
transform 1 0 14812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_162
timestamp 1676037725
transform 1 0 16008 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_166
timestamp 1676037725
transform 1 0 16376 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_172
timestamp 1676037725
transform 1 0 16928 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_178
timestamp 1676037725
transform 1 0 17480 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1676037725
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1676037725
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_213
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_238
timestamp 1676037725
transform 1 0 23000 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_246
timestamp 1676037725
transform 1 0 23736 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_259
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_266
timestamp 1676037725
transform 1 0 25576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_275
timestamp 1676037725
transform 1 0 26404 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1676037725
transform 1 0 27232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1676037725
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_300
timestamp 1676037725
transform 1 0 28704 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_316
timestamp 1676037725
transform 1 0 30176 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_331
timestamp 1676037725
transform 1 0 31556 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_344
timestamp 1676037725
transform 1 0 32752 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1676037725
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_397
timestamp 1676037725
transform 1 0 37628 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1676037725
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1676037725
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_66
timestamp 1676037725
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_78
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_88
timestamp 1676037725
transform 1 0 9200 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_103
timestamp 1676037725
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_122
timestamp 1676037725
transform 1 0 12328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_144
timestamp 1676037725
transform 1 0 14352 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_152
timestamp 1676037725
transform 1 0 15088 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_179
timestamp 1676037725
transform 1 0 17572 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_185
timestamp 1676037725
transform 1 0 18124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1676037725
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_198
timestamp 1676037725
transform 1 0 19320 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_206
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_218
timestamp 1676037725
transform 1 0 21160 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_236
timestamp 1676037725
transform 1 0 22816 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1676037725
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1676037725
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_301
timestamp 1676037725
transform 1 0 28796 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_308
timestamp 1676037725
transform 1 0 29440 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_320
timestamp 1676037725
transform 1 0 30544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_345
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_357
timestamp 1676037725
transform 1 0 33948 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_368
timestamp 1676037725
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_380
timestamp 1676037725
transform 1 0 36064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1676037725
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_36
timestamp 1676037725
transform 1 0 4416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_47
timestamp 1676037725
transform 1 0 5428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_56
timestamp 1676037725
transform 1 0 6256 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_67
timestamp 1676037725
transform 1 0 7268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_71
timestamp 1676037725
transform 1 0 7636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1676037725
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_106
timestamp 1676037725
transform 1 0 10856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_130
timestamp 1676037725
transform 1 0 13064 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_147
timestamp 1676037725
transform 1 0 14628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1676037725
transform 1 0 15272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_163
timestamp 1676037725
transform 1 0 16100 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_204
timestamp 1676037725
transform 1 0 19872 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_216
timestamp 1676037725
transform 1 0 20976 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_225
timestamp 1676037725
transform 1 0 21804 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_238
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_242
timestamp 1676037725
transform 1 0 23368 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_258
timestamp 1676037725
transform 1 0 24840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_271
timestamp 1676037725
transform 1 0 26036 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_279
timestamp 1676037725
transform 1 0 26772 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1676037725
transform 1 0 27416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_314
timestamp 1676037725
transform 1 0 29992 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_326
timestamp 1676037725
transform 1 0 31096 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_334
timestamp 1676037725
transform 1 0 31832 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_340
timestamp 1676037725
transform 1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_347
timestamp 1676037725
transform 1 0 33028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1676037725
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_379
timestamp 1676037725
transform 1 0 35972 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_400
timestamp 1676037725
transform 1 0 37904 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1676037725
transform 1 0 38456 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_41
timestamp 1676037725
transform 1 0 4876 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1676037725
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_64
timestamp 1676037725
transform 1 0 6992 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_72
timestamp 1676037725
transform 1 0 7728 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_84
timestamp 1676037725
transform 1 0 8832 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_92
timestamp 1676037725
transform 1 0 9568 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_103
timestamp 1676037725
transform 1 0 10580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_124
timestamp 1676037725
transform 1 0 12512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_136
timestamp 1676037725
transform 1 0 13616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_142
timestamp 1676037725
transform 1 0 14168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_158
timestamp 1676037725
transform 1 0 15640 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_179
timestamp 1676037725
transform 1 0 17572 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_191
timestamp 1676037725
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_203
timestamp 1676037725
transform 1 0 19780 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_207
timestamp 1676037725
transform 1 0 20148 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_213
timestamp 1676037725
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1676037725
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_232
timestamp 1676037725
transform 1 0 22448 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_240
timestamp 1676037725
transform 1 0 23184 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_262
timestamp 1676037725
transform 1 0 25208 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1676037725
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 1676037725
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_304
timestamp 1676037725
transform 1 0 29072 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_312
timestamp 1676037725
transform 1 0 29808 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_323
timestamp 1676037725
transform 1 0 30820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_343
timestamp 1676037725
transform 1 0 32660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1676037725
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_51
timestamp 1676037725
transform 1 0 5796 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_59
timestamp 1676037725
transform 1 0 6532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_73
timestamp 1676037725
transform 1 0 7820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1676037725
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1676037725
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1676037725
transform 1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_112
timestamp 1676037725
transform 1 0 11408 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_127
timestamp 1676037725
transform 1 0 12788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1676037725
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_150
timestamp 1676037725
transform 1 0 14904 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_159
timestamp 1676037725
transform 1 0 15732 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_171
timestamp 1676037725
transform 1 0 16836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_175
timestamp 1676037725
transform 1 0 17204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_182
timestamp 1676037725
transform 1 0 17848 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1676037725
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_204
timestamp 1676037725
transform 1 0 19872 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_216
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_228
timestamp 1676037725
transform 1 0 22080 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1676037725
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1676037725
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_266
timestamp 1676037725
transform 1 0 25576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_286
timestamp 1676037725
transform 1 0 27416 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_303
timestamp 1676037725
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_319
timestamp 1676037725
transform 1 0 30452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_331
timestamp 1676037725
transform 1 0 31556 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1676037725
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1676037725
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1676037725
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_373
timestamp 1676037725
transform 1 0 35420 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_384
timestamp 1676037725
transform 1 0 36432 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1676037725
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_63
timestamp 1676037725
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_70
timestamp 1676037725
transform 1 0 7544 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_76
timestamp 1676037725
transform 1 0 8096 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_84
timestamp 1676037725
transform 1 0 8832 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_94
timestamp 1676037725
transform 1 0 9752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1676037725
transform 1 0 10948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_119
timestamp 1676037725
transform 1 0 12052 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_123
timestamp 1676037725
transform 1 0 12420 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1676037725
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_175
timestamp 1676037725
transform 1 0 17204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_188
timestamp 1676037725
transform 1 0 18400 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_203
timestamp 1676037725
transform 1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_213
timestamp 1676037725
transform 1 0 20700 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_233
timestamp 1676037725
transform 1 0 22540 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_246
timestamp 1676037725
transform 1 0 23736 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_267
timestamp 1676037725
transform 1 0 25668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1676037725
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1676037725
transform 1 0 28152 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_307
timestamp 1676037725
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_320
timestamp 1676037725
transform 1 0 30544 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_324
timestamp 1676037725
transform 1 0 30912 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_345
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_355
timestamp 1676037725
transform 1 0 33764 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_370
timestamp 1676037725
transform 1 0 35144 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1676037725
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1676037725
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_404
timestamp 1676037725
transform 1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_45
timestamp 1676037725
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_55
timestamp 1676037725
transform 1 0 6164 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_63
timestamp 1676037725
transform 1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_92
timestamp 1676037725
transform 1 0 9568 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_100
timestamp 1676037725
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_108
timestamp 1676037725
transform 1 0 11040 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_116
timestamp 1676037725
transform 1 0 11776 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_158
timestamp 1676037725
transform 1 0 15640 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_170
timestamp 1676037725
transform 1 0 16744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_174
timestamp 1676037725
transform 1 0 17112 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_184
timestamp 1676037725
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_191
timestamp 1676037725
transform 1 0 18676 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_202
timestamp 1676037725
transform 1 0 19688 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_211
timestamp 1676037725
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_215
timestamp 1676037725
transform 1 0 20884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_224
timestamp 1676037725
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_236
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_271
timestamp 1676037725
transform 1 0 26036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_292
timestamp 1676037725
transform 1 0 27968 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1676037725
transform 1 0 28520 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1676037725
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_319
timestamp 1676037725
transform 1 0 30452 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_335
timestamp 1676037725
transform 1 0 31924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_347
timestamp 1676037725
transform 1 0 33028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1676037725
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_397
timestamp 1676037725
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1676037725
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_65
timestamp 1676037725
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_78
timestamp 1676037725
transform 1 0 8280 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_90
timestamp 1676037725
transform 1 0 9384 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_100
timestamp 1676037725
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_154
timestamp 1676037725
transform 1 0 15272 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_201
timestamp 1676037725
transform 1 0 19596 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_211
timestamp 1676037725
transform 1 0 20516 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1676037725
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 1676037725
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1676037725
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_251
timestamp 1676037725
transform 1 0 24196 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_257
timestamp 1676037725
transform 1 0 24748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1676037725
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_295
timestamp 1676037725
transform 1 0 28244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_303
timestamp 1676037725
transform 1 0 28980 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_310
timestamp 1676037725
transform 1 0 29624 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_344
timestamp 1676037725
transform 1 0 32752 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_355
timestamp 1676037725
transform 1 0 33764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_359
timestamp 1676037725
transform 1 0 34132 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_377
timestamp 1676037725
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1676037725
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_404
timestamp 1676037725
transform 1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_103
timestamp 1676037725
transform 1 0 10580 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_119
timestamp 1676037725
transform 1 0 12052 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 1676037725
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_178
timestamp 1676037725
transform 1 0 17480 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_205
timestamp 1676037725
transform 1 0 19964 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_218
timestamp 1676037725
transform 1 0 21160 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_226
timestamp 1676037725
transform 1 0 21896 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_234
timestamp 1676037725
transform 1 0 22632 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_269
timestamp 1676037725
transform 1 0 25852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_281
timestamp 1676037725
transform 1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_290
timestamp 1676037725
transform 1 0 27784 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1676037725
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_331
timestamp 1676037725
transform 1 0 31556 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_347
timestamp 1676037725
transform 1 0 33028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_359
timestamp 1676037725
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_400
timestamp 1676037725
transform 1 0 37904 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1676037725
transform 1 0 38456 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_74
timestamp 1676037725
transform 1 0 7912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_86
timestamp 1676037725
transform 1 0 9016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_90
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1676037725
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_124
timestamp 1676037725
transform 1 0 12512 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_136
timestamp 1676037725
transform 1 0 13616 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1676037725
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1676037725
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_174
timestamp 1676037725
transform 1 0 17112 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1676037725
transform 1 0 17848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_202
timestamp 1676037725
transform 1 0 19688 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_210
timestamp 1676037725
transform 1 0 20424 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1676037725
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_248
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_254
timestamp 1676037725
transform 1 0 24472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_267
timestamp 1676037725
transform 1 0 25668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1676037725
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_292
timestamp 1676037725
transform 1 0 27968 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_300
timestamp 1676037725
transform 1 0 28704 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_318
timestamp 1676037725
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1676037725
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_344
timestamp 1676037725
transform 1 0 32752 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_353
timestamp 1676037725
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_365
timestamp 1676037725
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_377
timestamp 1676037725
transform 1 0 35788 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1676037725
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_404
timestamp 1676037725
transform 1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_54
timestamp 1676037725
transform 1 0 6072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_74
timestamp 1676037725
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_118
timestamp 1676037725
transform 1 0 11960 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_135
timestamp 1676037725
transform 1 0 13524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_149
timestamp 1676037725
transform 1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_155
timestamp 1676037725
transform 1 0 15364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_180
timestamp 1676037725
transform 1 0 17664 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1676037725
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_205
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_214
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1676037725
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_261
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_268
timestamp 1676037725
transform 1 0 25760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_291
timestamp 1676037725
transform 1 0 27876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_320
timestamp 1676037725
transform 1 0 30544 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_328
timestamp 1676037725
transform 1 0 31280 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_336
timestamp 1676037725
transform 1 0 32016 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_349
timestamp 1676037725
transform 1 0 33212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_358
timestamp 1676037725
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_384
timestamp 1676037725
transform 1 0 36432 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1676037725
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_35
timestamp 1676037725
transform 1 0 4324 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1676037725
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1676037725
transform 1 0 13524 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1676037725
transform 1 0 16100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1676037725
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_180
timestamp 1676037725
transform 1 0 17664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1676037725
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1676037725
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_244
timestamp 1676037725
transform 1 0 23552 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_248
timestamp 1676037725
transform 1 0 23920 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_270
timestamp 1676037725
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1676037725
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_303
timestamp 1676037725
transform 1 0 28980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_309
timestamp 1676037725
transform 1 0 29532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_326
timestamp 1676037725
transform 1 0 31096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1676037725
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_356
timestamp 1676037725
transform 1 0 33856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_360
timestamp 1676037725
transform 1 0 34224 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_378
timestamp 1676037725
transform 1 0 35880 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1676037725
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1676037725
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_17
timestamp 1676037725
transform 1 0 2668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1676037725
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1676037725
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_68
timestamp 1676037725
transform 1 0 7360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_72
timestamp 1676037725
transform 1 0 7728 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_96
timestamp 1676037725
transform 1 0 9936 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1676037725
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1676037725
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1676037725
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1676037725
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_149
timestamp 1676037725
transform 1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1676037725
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1676037725
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1676037725
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1676037725
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1676037725
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_206
timestamp 1676037725
transform 1 0 20056 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_213
timestamp 1676037725
transform 1 0 20700 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1676037725
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_239
timestamp 1676037725
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1676037725
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_271
timestamp 1676037725
transform 1 0 26036 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1676037725
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1676037725
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_286
timestamp 1676037725
transform 1 0 27416 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_294
timestamp 1676037725
transform 1 0 28152 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1676037725
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1676037725
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_343
timestamp 1676037725
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_355
timestamp 1676037725
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_383
timestamp 1676037725
transform 1 0 36340 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1676037725
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_393
timestamp 1676037725
transform 1 0 37260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1676037725
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1676037725
transform 1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1676037725
transform 1 0 19596 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1676037725
transform -1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1676037725
transform -1 0 16100 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1676037725
transform 1 0 15088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_8  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_8  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10580 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_4  _0841_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7176 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8832 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_4  _0844_
timestamp 1676037725
transform -1 0 6072 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13708 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0846_
timestamp 1676037725
transform 1 0 12236 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1676037725
transform 1 0 7636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27324 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0849_
timestamp 1676037725
transform -1 0 23644 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0855_
timestamp 1676037725
transform 1 0 24564 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27416 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27784 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1676037725
transform 1 0 27048 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform -1 0 24748 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0862_
timestamp 1676037725
transform 1 0 26036 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26496 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0866_
timestamp 1676037725
transform -1 0 20792 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0867_
timestamp 1676037725
transform -1 0 23276 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_4  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0869_
timestamp 1676037725
transform -1 0 22724 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1676037725
transform 1 0 25116 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26864 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21344 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25484 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19688 0 -1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1676037725
transform -1 0 19412 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0878_
timestamp 1676037725
transform 1 0 27232 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0879_
timestamp 1676037725
transform -1 0 18860 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0880_
timestamp 1676037725
transform -1 0 26312 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0881_
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0882_
timestamp 1676037725
transform -1 0 23000 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1676037725
transform -1 0 20700 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0884_
timestamp 1676037725
transform -1 0 22448 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1676037725
transform -1 0 21528 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0887_
timestamp 1676037725
transform 1 0 22632 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1676037725
transform -1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0889_
timestamp 1676037725
transform 1 0 24564 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1676037725
transform -1 0 24104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25576 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0892_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1676037725
transform 1 0 36708 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0894_
timestamp 1676037725
transform -1 0 24104 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0895_
timestamp 1676037725
transform -1 0 19872 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1676037725
transform -1 0 25484 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0897_
timestamp 1676037725
transform -1 0 18400 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0898_
timestamp 1676037725
transform -1 0 19320 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1676037725
transform -1 0 23644 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0900_
timestamp 1676037725
transform -1 0 22080 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0901_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0903_
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1676037725
transform -1 0 20424 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0905_
timestamp 1676037725
transform -1 0 25668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27416 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0908_
timestamp 1676037725
transform -1 0 24656 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0909_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21068 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23828 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20976 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1676037725
transform -1 0 20332 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0915_
timestamp 1676037725
transform -1 0 19688 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18492 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0917_
timestamp 1676037725
transform 1 0 24840 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1676037725
transform -1 0 21528 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0920_
timestamp 1676037725
transform -1 0 16468 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25392 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1676037725
transform 1 0 27048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0925_
timestamp 1676037725
transform 1 0 18032 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__o22ai_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0930_
timestamp 1676037725
transform -1 0 23276 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0931_
timestamp 1676037725
transform 1 0 26956 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0932_
timestamp 1676037725
transform -1 0 27416 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21160 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_4  _0936_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26956 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_8  _0940_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__and4_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1676037725
transform 1 0 34132 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 35512 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _0945_
timestamp 1676037725
transform 1 0 29900 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _0946_
timestamp 1676037725
transform -1 0 35144 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__a221oi_4  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35052 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0948_
timestamp 1676037725
transform -1 0 28060 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0949_
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0950_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0951_
timestamp 1676037725
transform -1 0 24104 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform -1 0 24104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22540 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0954_
timestamp 1676037725
transform -1 0 23736 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1676037725
transform 1 0 22540 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _0957_
timestamp 1676037725
transform 1 0 25576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28428 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0959_
timestamp 1676037725
transform -1 0 25944 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform -1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1676037725
transform 1 0 33948 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1676037725
transform -1 0 35420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0963_
timestamp 1676037725
transform 1 0 35052 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1676037725
transform -1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _0965_
timestamp 1676037725
transform 1 0 27600 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0966_
timestamp 1676037725
transform -1 0 27232 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _0967_
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0968_
timestamp 1676037725
transform -1 0 21160 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21804 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1676037725
transform -1 0 19872 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20700 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20240 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0973_
timestamp 1676037725
transform 1 0 21160 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0974_
timestamp 1676037725
transform 1 0 22080 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20608 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _0978_
timestamp 1676037725
transform -1 0 17020 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0980_
timestamp 1676037725
transform -1 0 18676 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1676037725
transform -1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0982_
timestamp 1676037725
transform 1 0 17296 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1676037725
transform 1 0 17204 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1676037725
transform -1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0987_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22264 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1676037725
transform -1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0990_
timestamp 1676037725
transform 1 0 11500 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1676037725
transform -1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1676037725
transform 1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0994_
timestamp 1676037725
transform -1 0 15824 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1676037725
transform -1 0 14812 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0996_
timestamp 1676037725
transform -1 0 14536 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1676037725
transform -1 0 34316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0999_
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28152 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1002_
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1003_
timestamp 1676037725
transform -1 0 22080 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21712 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1005_
timestamp 1676037725
transform -1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1676037725
transform -1 0 22632 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1009_
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1676037725
transform -1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1012_
timestamp 1676037725
transform 1 0 20884 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1676037725
transform 1 0 19964 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1676037725
transform -1 0 20056 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1676037725
transform 1 0 33764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1016_
timestamp 1676037725
transform -1 0 35604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1017_
timestamp 1676037725
transform 1 0 35512 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1676037725
transform -1 0 28796 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1019_
timestamp 1676037725
transform -1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1020_
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1021_
timestamp 1676037725
transform -1 0 22080 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1676037725
transform -1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1023_
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1676037725
transform -1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1025_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1026_
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20884 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1028_
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1676037725
transform 1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1031_
timestamp 1676037725
transform -1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1032_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 1676037725
transform 1 0 24380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1676037725
transform 1 0 25760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1035_
timestamp 1676037725
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1036_
timestamp 1676037725
transform -1 0 26588 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1676037725
transform -1 0 28704 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1038_
timestamp 1676037725
transform -1 0 26128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1039_
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1040_
timestamp 1676037725
transform -1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1676037725
transform -1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1042_
timestamp 1676037725
transform 1 0 20148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1676037725
transform -1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 1676037725
transform -1 0 19780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1046_
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1047_
timestamp 1676037725
transform -1 0 19596 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1048_
timestamp 1676037725
transform -1 0 18952 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1676037725
transform -1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1676037725
transform -1 0 29992 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1676037725
transform 1 0 30360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1052_
timestamp 1676037725
transform -1 0 30820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1054_
timestamp 1676037725
transform 1 0 28152 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1055_
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1056_
timestamp 1676037725
transform -1 0 22724 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1676037725
transform -1 0 18492 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1059_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1676037725
transform -1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 1676037725
transform -1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1063_
timestamp 1676037725
transform -1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21160 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1066_
timestamp 1676037725
transform 1 0 25944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1676037725
transform -1 0 25392 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1676037725
transform -1 0 25944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1069_
timestamp 1676037725
transform -1 0 26128 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1676037725
transform -1 0 26588 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1071_
timestamp 1676037725
transform -1 0 26036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1073_
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1075_
timestamp 1676037725
transform 1 0 15364 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _1076_
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1077_
timestamp 1676037725
transform 1 0 14352 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15916 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _1079_
timestamp 1676037725
transform -1 0 13800 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1080_
timestamp 1676037725
transform -1 0 15456 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1676037725
transform -1 0 14720 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1082_
timestamp 1676037725
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1676037725
transform -1 0 16744 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1085_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1676037725
transform 1 0 22816 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1087_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1089_
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1090_
timestamp 1676037725
transform -1 0 14720 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1676037725
transform -1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1092_
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _1093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _1094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _1095_
timestamp 1676037725
transform -1 0 15824 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1096_
timestamp 1676037725
transform -1 0 16652 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _1097_
timestamp 1676037725
transform -1 0 20056 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1098_
timestamp 1676037725
transform -1 0 18952 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1099_
timestamp 1676037725
transform 1 0 17848 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1676037725
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1104_
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1105_
timestamp 1676037725
transform -1 0 16192 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1106_
timestamp 1676037725
transform 1 0 16652 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1676037725
transform -1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1108_
timestamp 1676037725
transform -1 0 21160 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__o211ai_4  _1110_
timestamp 1676037725
transform -1 0 14904 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1676037725
transform 1 0 28244 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1676037725
transform -1 0 29716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1113_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1676037725
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1676037725
transform -1 0 27416 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1116_
timestamp 1676037725
transform 1 0 26496 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _1117_
timestamp 1676037725
transform -1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1676037725
transform -1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1676037725
transform 1 0 19596 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1120_
timestamp 1676037725
transform -1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1122_
timestamp 1676037725
transform -1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1124_
timestamp 1676037725
transform -1 0 13892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1676037725
transform -1 0 14260 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1126_
timestamp 1676037725
transform -1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1676037725
transform 1 0 11776 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1130_
timestamp 1676037725
transform -1 0 22724 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1132_
timestamp 1676037725
transform -1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1133_
timestamp 1676037725
transform 1 0 16836 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1676037725
transform 1 0 14536 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1676037725
transform -1 0 12880 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1138_
timestamp 1676037725
transform -1 0 13064 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1676037725
transform -1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1140_
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1141_
timestamp 1676037725
transform -1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1676037725
transform -1 0 10764 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1143_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1676037725
transform -1 0 13156 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1145_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1148_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1676037725
transform -1 0 20240 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1151_
timestamp 1676037725
transform 1 0 29716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1676037725
transform -1 0 27232 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1153_
timestamp 1676037725
transform 1 0 28336 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1154_
timestamp 1676037725
transform 1 0 25760 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1155_
timestamp 1676037725
transform -1 0 29072 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _1156_
timestamp 1676037725
transform 1 0 31280 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1157_
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__o31ai_4  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_8  _1159_
timestamp 1676037725
transform 1 0 28980 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1676037725
transform -1 0 32292 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1161_
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1676037725
transform 1 0 25944 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1164_
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1166_
timestamp 1676037725
transform 1 0 25852 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1676037725
transform -1 0 27048 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1676037725
transform -1 0 28152 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1676037725
transform 1 0 28704 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28428 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1172_
timestamp 1676037725
transform -1 0 27416 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_2  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31004 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32016 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1676037725
transform 1 0 32568 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1676037725
transform 1 0 32660 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1676037725
transform -1 0 33764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1178_
timestamp 1676037725
transform -1 0 29256 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1676037725
transform 1 0 31188 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _1180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 34132 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__or3b_2  _1181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33304 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1676037725
transform 1 0 33028 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30636 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1676037725
transform 1 0 32752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1185_
timestamp 1676037725
transform -1 0 33580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1676037725
transform -1 0 33672 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1187_
timestamp 1676037725
transform 1 0 33304 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1188_
timestamp 1676037725
transform 1 0 32292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1189_
timestamp 1676037725
transform -1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1676037725
transform 1 0 33120 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1191_
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1192_
timestamp 1676037725
transform -1 0 33120 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1193_
timestamp 1676037725
transform 1 0 32568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1196_
timestamp 1676037725
transform 1 0 32660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1197_
timestamp 1676037725
transform 1 0 33764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1676037725
transform 1 0 33764 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1199_
timestamp 1676037725
transform 1 0 33580 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1200_
timestamp 1676037725
transform 1 0 31924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1201_
timestamp 1676037725
transform -1 0 33672 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1202_
timestamp 1676037725
transform -1 0 34408 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1676037725
transform -1 0 35328 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1676037725
transform -1 0 34408 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1205_
timestamp 1676037725
transform -1 0 31280 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1676037725
transform -1 0 31464 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1676037725
transform 1 0 29808 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1208_
timestamp 1676037725
transform 1 0 31648 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1209_
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1210_
timestamp 1676037725
transform 1 0 29716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1676037725
transform 1 0 31004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1676037725
transform 1 0 32108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1676037725
transform 1 0 32476 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1216_
timestamp 1676037725
transform 1 0 30728 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1676037725
transform 1 0 32108 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1218_
timestamp 1676037725
transform 1 0 29716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1676037725
transform 1 0 30636 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1220_
timestamp 1676037725
transform 1 0 32292 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1676037725
transform -1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1676037725
transform 1 0 32752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1223_
timestamp 1676037725
transform 1 0 30084 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1224_
timestamp 1676037725
transform 1 0 31004 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1225_
timestamp 1676037725
transform 1 0 33120 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1226_
timestamp 1676037725
transform -1 0 31556 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1227_
timestamp 1676037725
transform 1 0 31188 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1228_
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1676037725
transform 1 0 32660 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1230_
timestamp 1676037725
transform -1 0 33580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1231_
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1232_
timestamp 1676037725
transform 1 0 30820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1676037725
transform 1 0 32476 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1676037725
transform 1 0 32752 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1676037725
transform 1 0 33580 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1236_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1676037725
transform 1 0 30636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp 1676037725
transform 1 0 31372 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1240_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1676037725
transform -1 0 19964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1676037725
transform 1 0 9476 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1243_
timestamp 1676037725
transform -1 0 6072 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1676037725
transform 1 0 6808 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1245_
timestamp 1676037725
transform 1 0 11224 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1246_
timestamp 1676037725
transform -1 0 10948 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1247_
timestamp 1676037725
transform 1 0 7176 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1676037725
transform -1 0 6164 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1676037725
transform 1 0 5244 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1250_
timestamp 1676037725
transform 1 0 5152 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1676037725
transform 1 0 4416 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1252_
timestamp 1676037725
transform 1 0 6532 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _1253_
timestamp 1676037725
transform 1 0 4784 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1254_
timestamp 1676037725
transform -1 0 6072 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1676037725
transform -1 0 9568 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1256_
timestamp 1676037725
transform -1 0 8648 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _1257_
timestamp 1676037725
transform -1 0 8832 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1258_
timestamp 1676037725
transform 1 0 9844 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1676037725
transform 1 0 6532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1260_
timestamp 1676037725
transform -1 0 7268 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1261_
timestamp 1676037725
transform 1 0 13248 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1676037725
transform 1 0 25760 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1264_
timestamp 1676037725
transform -1 0 16008 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 1676037725
transform -1 0 16376 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1676037725
transform 1 0 4784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1268_
timestamp 1676037725
transform 1 0 9936 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1269_
timestamp 1676037725
transform 1 0 7360 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1270_
timestamp 1676037725
transform 1 0 10304 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1676037725
transform 1 0 13064 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1676037725
transform 1 0 15180 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1676037725
transform -1 0 7544 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1676037725
transform 1 0 12512 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1676037725
transform -1 0 6808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1277_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1676037725
transform -1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1279_
timestamp 1676037725
transform 1 0 11684 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1280_
timestamp 1676037725
transform 1 0 10396 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1676037725
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1283_
timestamp 1676037725
transform -1 0 24104 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1676037725
transform 1 0 16468 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1285_
timestamp 1676037725
transform -1 0 18952 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1676037725
transform -1 0 18124 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1676037725
transform -1 0 17940 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1288_
timestamp 1676037725
transform 1 0 12604 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1289_
timestamp 1676037725
transform 1 0 20240 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1290_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1676037725
transform 1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1676037725
transform -1 0 16100 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1293_
timestamp 1676037725
transform -1 0 5336 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1294_
timestamp 1676037725
transform 1 0 8924 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1676037725
transform 1 0 10212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1297_
timestamp 1676037725
transform 1 0 14076 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1676037725
transform -1 0 18584 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1676037725
transform -1 0 5704 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1676037725
transform -1 0 4784 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1301_
timestamp 1676037725
transform -1 0 8648 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1676037725
transform 1 0 10304 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1676037725
transform 1 0 12696 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1305_
timestamp 1676037725
transform 1 0 8832 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1306_
timestamp 1676037725
transform -1 0 6072 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1307_
timestamp 1676037725
transform 1 0 5704 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1676037725
transform 1 0 11868 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1309_
timestamp 1676037725
transform -1 0 12236 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1676037725
transform -1 0 10396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_2  _1312_
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1313_
timestamp 1676037725
transform 1 0 21528 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1314_
timestamp 1676037725
transform 1 0 10304 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1315_
timestamp 1676037725
transform 1 0 19228 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14352 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 1676037725
transform -1 0 12788 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1676037725
transform 1 0 7452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1676037725
transform 1 0 10396 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1321_
timestamp 1676037725
transform 1 0 8648 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1322_
timestamp 1676037725
transform -1 0 4416 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1676037725
transform 1 0 5796 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1324_
timestamp 1676037725
transform 1 0 7728 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1325_
timestamp 1676037725
transform -1 0 8280 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1326_
timestamp 1676037725
transform -1 0 6992 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1327_
timestamp 1676037725
transform -1 0 6072 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11500 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1329_
timestamp 1676037725
transform -1 0 12512 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1676037725
transform -1 0 9936 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1331_
timestamp 1676037725
transform -1 0 10028 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1332_
timestamp 1676037725
transform 1 0 9752 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1333_
timestamp 1676037725
transform 1 0 11868 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1334_
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1337_
timestamp 1676037725
transform 1 0 19136 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1338_
timestamp 1676037725
transform 1 0 14076 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1339_
timestamp 1676037725
transform -1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1676037725
transform 1 0 14720 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1676037725
transform 1 0 15272 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1676037725
transform 1 0 11960 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1676037725
transform 1 0 13432 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1344_
timestamp 1676037725
transform 1 0 10764 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1676037725
transform 1 0 16836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1676037725
transform 1 0 13524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1348_
timestamp 1676037725
transform 1 0 14076 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1676037725
transform 1 0 15364 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1350_
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1676037725
transform -1 0 19964 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1676037725
transform 1 0 15088 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1353_
timestamp 1676037725
transform 1 0 15364 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1676037725
transform 1 0 22080 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1355_
timestamp 1676037725
transform 1 0 20976 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1356_
timestamp 1676037725
transform -1 0 24288 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1676037725
transform -1 0 17848 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1676037725
transform -1 0 17756 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1676037725
transform -1 0 12420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1676037725
transform 1 0 17296 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1361_
timestamp 1676037725
transform -1 0 13800 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_4  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1676037725
transform 1 0 18400 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1365_
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1366_
timestamp 1676037725
transform 1 0 18216 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1367_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1368_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _1369_
timestamp 1676037725
transform 1 0 29440 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _1370_
timestamp 1676037725
transform 1 0 27600 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_4  _1371_
timestamp 1676037725
transform 1 0 27784 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1372_
timestamp 1676037725
transform 1 0 28244 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1676037725
transform 1 0 28980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1374_
timestamp 1676037725
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1375_
timestamp 1676037725
transform 1 0 28428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1376_
timestamp 1676037725
transform -1 0 26680 0 -1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1377_
timestamp 1676037725
transform 1 0 30084 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_4  _1378_
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1676037725
transform 1 0 30912 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _1380_
timestamp 1676037725
transform 1 0 30820 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _1381_
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1382_
timestamp 1676037725
transform -1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1383_
timestamp 1676037725
transform -1 0 32936 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1676037725
transform -1 0 35604 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1385_
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1386_
timestamp 1676037725
transform -1 0 35236 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1387_
timestamp 1676037725
transform 1 0 35144 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_
timestamp 1676037725
transform -1 0 35696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1389_
timestamp 1676037725
transform -1 0 36340 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1390_
timestamp 1676037725
transform 1 0 34960 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1391_
timestamp 1676037725
transform -1 0 36156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1392_
timestamp 1676037725
transform -1 0 36708 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1394_
timestamp 1676037725
transform -1 0 33948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1395_
timestamp 1676037725
transform -1 0 35880 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1397_
timestamp 1676037725
transform -1 0 36156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1398_
timestamp 1676037725
transform -1 0 36156 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1399_
timestamp 1676037725
transform 1 0 34868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1400_
timestamp 1676037725
transform -1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1676037725
transform -1 0 36616 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1402_
timestamp 1676037725
transform 1 0 31188 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1403_
timestamp 1676037725
transform -1 0 31740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1404_
timestamp 1676037725
transform -1 0 32936 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1405_
timestamp 1676037725
transform -1 0 31280 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1406_
timestamp 1676037725
transform 1 0 29808 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1676037725
transform -1 0 34132 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1676037725
transform -1 0 32936 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 1676037725
transform 1 0 33948 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1410_
timestamp 1676037725
transform -1 0 35604 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1676037725
transform -1 0 35420 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 1676037725
transform 1 0 34868 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1413_
timestamp 1676037725
transform 1 0 35512 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 1676037725
transform 1 0 34868 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1676037725
transform 1 0 35604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1417_
timestamp 1676037725
transform 1 0 35236 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 1676037725
transform 1 0 34868 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1676037725
transform 1 0 35696 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 1676037725
transform 1 0 34500 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1421_
timestamp 1676037725
transform 1 0 35512 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1676037725
transform 1 0 31924 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1676037725
transform 1 0 33028 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 26680 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__o21bai_4  _1425_
timestamp 1676037725
transform -1 0 27600 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1676037725
transform -1 0 27784 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1676037725
transform 1 0 26128 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1431_
timestamp 1676037725
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1432_
timestamp 1676037725
transform -1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1676037725
transform -1 0 30360 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1676037725
transform -1 0 29256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1436_
timestamp 1676037725
transform -1 0 29440 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 1676037725
transform -1 0 28612 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1676037725
transform 1 0 28336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _1439_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29440 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 1676037725
transform -1 0 28152 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1676037725
transform -1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1442_
timestamp 1676037725
transform -1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1443_
timestamp 1676037725
transform -1 0 29072 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1444_
timestamp 1676037725
transform -1 0 29072 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1445_
timestamp 1676037725
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 1676037725
transform -1 0 29808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1676037725
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1448_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1676037725
transform 1 0 26128 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1450_
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _1451_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29992 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1676037725
transform -1 0 29072 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1453_
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1454_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _1455_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _1457_
timestamp 1676037725
transform -1 0 29532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1458_
timestamp 1676037725
transform -1 0 24932 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1676037725
transform 1 0 22632 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1461_
timestamp 1676037725
transform 1 0 23092 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1462_
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1463_
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1466_
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1676037725
transform 1 0 30084 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1676037725
transform -1 0 24012 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1469_
timestamp 1676037725
transform -1 0 23736 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1470_
timestamp 1676037725
transform -1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1471_
timestamp 1676037725
transform 1 0 23460 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1676037725
transform -1 0 26588 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1474_
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1475_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1676037725
transform 1 0 30728 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1477_
timestamp 1676037725
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1478_
timestamp 1676037725
transform 1 0 32568 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1479_
timestamp 1676037725
transform -1 0 31648 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1676037725
transform 1 0 32660 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1482_
timestamp 1676037725
transform 1 0 23368 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1676037725
transform -1 0 23828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1676037725
transform -1 0 25024 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1485_
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31372 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1676037725
transform 1 0 33120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1676037725
transform 1 0 23000 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1490_
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1491_
timestamp 1676037725
transform -1 0 25208 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1676037725
transform 1 0 33396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1494_
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1676037725
transform 1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1497_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _1498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25116 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1676037725
transform 1 0 27140 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1500_
timestamp 1676037725
transform -1 0 30728 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1676037725
transform 1 0 24748 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1676037725
transform 1 0 27876 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1676037725
transform 1 0 23184 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1676037725
transform 1 0 35236 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1676037725
transform 1 0 30728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1676037725
transform 1 0 35052 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1509_
timestamp 1676037725
transform -1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1510_
timestamp 1676037725
transform -1 0 21528 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1676037725
transform 1 0 27600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1512_
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1513_
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1676037725
transform 1 0 20792 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1515_
timestamp 1676037725
transform 1 0 20148 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1516_
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1517_
timestamp 1676037725
transform -1 0 27876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1518_
timestamp 1676037725
transform 1 0 26128 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1676037725
transform 1 0 31004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1676037725
transform 1 0 37076 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1527_
timestamp 1676037725
transform -1 0 16928 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1528_
timestamp 1676037725
transform 1 0 14628 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1529_
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1530_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1536_
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1537_
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1539_
timestamp 1676037725
transform -1 0 22540 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1540_
timestamp 1676037725
transform 1 0 20976 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1676037725
transform 1 0 18584 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1545_
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 1676037725
transform -1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1676037725
transform 1 0 12052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1555_
timestamp 1676037725
transform -1 0 18952 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1556_
timestamp 1676037725
transform -1 0 20792 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1676037725
transform 1 0 19872 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1676037725
transform -1 0 20608 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1676037725
transform 1 0 21068 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1560_
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 1676037725
transform 1 0 9200 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1676037725
transform 1 0 9936 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1564_
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1565_
timestamp 1676037725
transform 1 0 14352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1566_
timestamp 1676037725
transform -1 0 16100 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1676037725
transform -1 0 16284 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1568_
timestamp 1676037725
transform -1 0 23920 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1676037725
transform 1 0 5152 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1676037725
transform 1 0 5152 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1676037725
transform 1 0 7084 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1676037725
transform 1 0 9476 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1574_
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1676037725
transform -1 0 13524 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1676037725
transform 1 0 22080 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1676037725
transform -1 0 27416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1578_
timestamp 1676037725
transform 1 0 26312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1579_
timestamp 1676037725
transform -1 0 12144 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1580_
timestamp 1676037725
transform -1 0 6992 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1581_
timestamp 1676037725
transform 1 0 7820 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1676037725
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1583_
timestamp 1676037725
transform -1 0 8464 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1676037725
transform -1 0 5428 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1676037725
transform 1 0 5612 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1586_
timestamp 1676037725
transform -1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1676037725
transform -1 0 9568 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1588_
timestamp 1676037725
transform -1 0 8648 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1676037725
transform 1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1590_
timestamp 1676037725
transform 1 0 6532 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1591_
timestamp 1676037725
transform -1 0 7360 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1592_
timestamp 1676037725
transform 1 0 5060 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1593_
timestamp 1676037725
transform -1 0 5612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 1676037725
transform 1 0 4048 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1595_
timestamp 1676037725
transform 1 0 28244 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1596_
timestamp 1676037725
transform 1 0 4784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1598_
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1599_
timestamp 1676037725
transform -1 0 5612 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1600_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1676037725
transform -1 0 13248 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1602_
timestamp 1676037725
transform 1 0 5428 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1676037725
transform 1 0 5152 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1604_
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 1676037725
transform -1 0 8004 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1676037725
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1676037725
transform 1 0 6532 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1609_
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1610_
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1676037725
transform -1 0 4692 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1612_
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1676037725
transform -1 0 8372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1614_
timestamp 1676037725
transform -1 0 9568 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1615_
timestamp 1676037725
transform -1 0 9476 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1616_
timestamp 1676037725
transform 1 0 14720 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1617_
timestamp 1676037725
transform 1 0 2944 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1618_
timestamp 1676037725
transform 1 0 3956 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1619_
timestamp 1676037725
transform 1 0 9200 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp 1676037725
transform -1 0 6256 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1624_
timestamp 1676037725
transform -1 0 11224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1676037725
transform 1 0 10304 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1626_
timestamp 1676037725
transform 1 0 8280 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1627_
timestamp 1676037725
transform 1 0 9936 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1630_
timestamp 1676037725
transform -1 0 7268 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1676037725
transform -1 0 6808 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1676037725
transform 1 0 6532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1676037725
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 1676037725
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1636_
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1637_
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1638_
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1639_
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1640_
timestamp 1676037725
transform -1 0 6900 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1641_
timestamp 1676037725
transform -1 0 7912 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1642_
timestamp 1676037725
transform 1 0 7728 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1643_
timestamp 1676037725
transform -1 0 7820 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1676037725
transform -1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1645_
timestamp 1676037725
transform -1 0 8464 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1646_
timestamp 1676037725
transform 1 0 7728 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1676037725
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1676037725
transform 1 0 8280 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1651_
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1652_
timestamp 1676037725
transform 1 0 9292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1676037725
transform 1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1676037725
transform 1 0 10580 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1676037725
transform 1 0 8372 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp 1676037725
transform 1 0 10212 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1657_
timestamp 1676037725
transform 1 0 10120 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1658_
timestamp 1676037725
transform -1 0 9752 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1676037725
transform 1 0 10580 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1676037725
transform -1 0 9752 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1676037725
transform 1 0 13248 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1676037725
transform -1 0 13432 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1663_
timestamp 1676037725
transform -1 0 30544 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1664_
timestamp 1676037725
transform 1 0 28888 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1676037725
transform 1 0 32752 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1676037725
transform 1 0 37444 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1676037725
transform -1 0 36984 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1676037725
transform 1 0 37444 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1676037725
transform 1 0 37444 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1676037725
transform 1 0 37444 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1673_
timestamp 1676037725
transform -1 0 30544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1676037725
transform 1 0 30360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1676037725
transform 1 0 24472 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1676037725
transform 1 0 35512 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1676037725
transform 1 0 27508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1682_
timestamp 1676037725
transform -1 0 30360 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1676037725
transform 1 0 24748 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1676037725
transform 1 0 28244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1676037725
transform 1 0 32292 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1676037725
transform 1 0 28428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1676037725
transform -1 0 14996 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1676037725
transform -1 0 17112 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1676037725
transform -1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1676037725
transform -1 0 19688 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1676037725
transform -1 0 25760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1698_
timestamp 1676037725
transform 1 0 15548 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1701_
timestamp 1676037725
transform -1 0 25944 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1676037725
transform 1 0 29716 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1676037725
transform -1 0 27876 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1676037725
transform 1 0 32292 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1676037725
transform 1 0 30820 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1676037725
transform 1 0 32660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1676037725
transform 1 0 32936 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1676037725
transform 1 0 26404 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1676037725
transform 1 0 24380 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1676037725
transform 1 0 27324 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1676037725
transform 1 0 34960 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1676037725
transform 1 0 32936 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1676037725
transform 1 0 26496 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9384 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1719_
timestamp 1676037725
transform 1 0 8740 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1676037725
transform 1 0 21528 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1721_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1722_
timestamp 1676037725
transform 1 0 16192 0 1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1723_
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1724_
timestamp 1676037725
transform -1 0 18860 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1725_
timestamp 1676037725
transform 1 0 20700 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1726_
timestamp 1676037725
transform 1 0 10580 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1727_
timestamp 1676037725
transform 1 0 12052 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1676037725
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1676037725
transform 1 0 7544 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 27784 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1731_
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1732_
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1733_
timestamp 1676037725
transform 1 0 34592 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1734_
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1735_
timestamp 1676037725
transform 1 0 33672 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1736_
timestamp 1676037725
transform 1 0 34684 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1737_
timestamp 1676037725
transform -1 0 36708 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1738_
timestamp 1676037725
transform 1 0 34132 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1739_
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1740_
timestamp 1676037725
transform 1 0 33580 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1741_
timestamp 1676037725
transform 1 0 32752 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1742_
timestamp 1676037725
transform 1 0 34224 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1743_
timestamp 1676037725
transform 1 0 34868 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1744_
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1745_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1676037725
transform 1 0 30360 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1748_
timestamp 1676037725
transform 1 0 36708 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1676037725
transform 1 0 36708 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1676037725
transform 1 0 36708 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1676037725
transform 1 0 36800 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1676037725
transform 1 0 36800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1676037725
transform 1 0 36616 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1754_
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1676037725
transform -1 0 23460 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1759_
timestamp 1676037725
transform 1 0 11500 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1760_
timestamp 1676037725
transform 1 0 20700 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1676037725
transform 1 0 4600 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1676037725
transform 1 0 4324 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1676037725
transform 1 0 6440 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1676037725
transform 1 0 10488 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1676037725
transform 1 0 9108 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1676037725
transform 1 0 8188 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1676037725
transform -1 0 13524 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1676037725
transform 1 0 22080 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1770_
timestamp 1676037725
transform 1 0 26128 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1676037725
transform 1 0 27508 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1676037725
transform 1 0 12328 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1676037725
transform 1 0 2760 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1676037725
transform 1 0 2760 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1676037725
transform 1 0 14536 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1778_
timestamp 1676037725
transform 1 0 2760 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1779_
timestamp 1676037725
transform 1 0 8372 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1780_
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1676037725
transform 1 0 4600 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1676037725
transform 1 0 11316 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1676037725
transform 1 0 12696 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1676037725
transform 1 0 7820 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1789_
timestamp 1676037725
transform -1 0 7912 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1676037725
transform 1 0 4416 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1676037725
transform 1 0 11040 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1676037725
transform -1 0 11592 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1800_
timestamp 1676037725
transform 1 0 14260 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1676037725
transform 1 0 16560 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1676037725
transform -1 0 31096 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1806_
timestamp 1676037725
transform 1 0 28796 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1676037725
transform -1 0 32384 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1676037725
transform 1 0 36524 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1676037725
transform 1 0 36616 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1810_
timestamp 1676037725
transform 1 0 36800 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1811_
timestamp 1676037725
transform 1 0 36340 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1812_
timestamp 1676037725
transform 1 0 36800 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1813_
timestamp 1676037725
transform 1 0 36340 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1814_
timestamp 1676037725
transform 1 0 36800 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1676037725
transform 1 0 30176 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1676037725
transform 1 0 35052 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1676037725
transform 1 0 30912 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1676037725
transform 1 0 36708 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1676037725
transform 1 0 36800 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1676037725
transform 1 0 27508 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1676037725
transform 1 0 22172 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1676037725
transform 1 0 36800 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22448 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform -1 0 8464 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform 1 0 11960 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform -1 0 13800 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform -1 0 8280 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform -1 0 8832 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform -1 0 13524 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform -1 0 14352 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform -1 0 26772 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform -1 0 28152 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform -1 0 33856 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform -1 0 33948 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 32568 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform -1 0 31832 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 34960 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform 1 0 34776 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 33120 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1676037725
transform -1 0 19412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1676037725
transform -1 0 30912 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19596 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout45
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1676037725
transform -1 0 12052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 1676037725
transform -1 0 6072 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout49
timestamp 1676037725
transform -1 0 21712 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1676037725
transform -1 0 9752 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1676037725
transform -1 0 29072 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout52
timestamp 1676037725
transform -1 0 7912 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout53
timestamp 1676037725
transform -1 0 25484 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1676037725
transform 1 0 28336 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout55
timestamp 1676037725
transform -1 0 11776 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1676037725
transform -1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout57
timestamp 1676037725
transform -1 0 14444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1676037725
transform -1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1676037725
transform -1 0 16376 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout60
timestamp 1676037725
transform 1 0 27140 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout61
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout62
timestamp 1676037725
transform 1 0 14260 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1676037725
transform -1 0 14720 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout64
timestamp 1676037725
transform 1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout65
timestamp 1676037725
transform -1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout66
timestamp 1676037725
transform 1 0 24564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1676037725
transform -1 0 29624 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout69
timestamp 1676037725
transform 1 0 29716 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  fanout70
timestamp 1676037725
transform -1 0 10948 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout71
timestamp 1676037725
transform -1 0 30268 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1676037725
transform 1 0 6992 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout73
timestamp 1676037725
transform -1 0 26036 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout74
timestamp 1676037725
transform 1 0 27324 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout76
timestamp 1676037725
transform -1 0 27968 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout77
timestamp 1676037725
transform 1 0 27140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout78
timestamp 1676037725
transform -1 0 27968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout79
timestamp 1676037725
transform 1 0 28520 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 1676037725
transform -1 0 14904 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout81
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout82
timestamp 1676037725
transform 1 0 20148 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout83
timestamp 1676037725
transform 1 0 22080 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1676037725
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout85
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout86
timestamp 1676037725
transform -1 0 19964 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout87
timestamp 1676037725
transform 1 0 23644 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout88
timestamp 1676037725
transform 1 0 17480 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout89
timestamp 1676037725
transform 1 0 26036 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout90
timestamp 1676037725
transform 1 0 18032 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1676037725
transform 1 0 1840 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1676037725
transform 1 0 6532 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1676037725
transform -1 0 8648 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input4
timestamp 1676037725
transform 1 0 11776 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input5
timestamp 1676037725
transform 1 0 15088 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  input7
timestamp 1676037725
transform 1 0 21988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  input8
timestamp 1676037725
transform 1 0 25024 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform -1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input11
timestamp 1676037725
transform -1 0 38364 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 36432 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 37812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 37812 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 37812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1676037725
transform 1 0 37812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1676037725
transform 1 0 37812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1676037725
transform 1 0 37812 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1676037725
transform 1 0 37812 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1676037725
transform 1 0 37812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp 1676037725
transform 1 0 37812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp 1676037725
transform 1 0 37812 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp 1676037725
transform 1 0 37812 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp 1676037725
transform -1 0 36984 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp 1676037725
transform 1 0 37812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp 1676037725
transform 1 0 37812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp 1676037725
transform 1 0 37812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp 1676037725
transform 1 0 37812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp 1676037725
transform 1 0 37812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp 1676037725
transform 1 0 37812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_92
timestamp 1676037725
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
<< labels >>
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 39200 38224 40000 38344 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal3 s 39200 1504 40000 1624 0 FreeSans 480 0 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal3 s 39200 15104 40000 15224 0 FreeSans 480 0 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal3 s 39200 16464 40000 16584 0 FreeSans 480 0 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal3 s 39200 17824 40000 17944 0 FreeSans 480 0 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal3 s 39200 19184 40000 19304 0 FreeSans 480 0 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal3 s 39200 20544 40000 20664 0 FreeSans 480 0 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal3 s 39200 21904 40000 22024 0 FreeSans 480 0 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal3 s 39200 23264 40000 23384 0 FreeSans 480 0 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal3 s 39200 24624 40000 24744 0 FreeSans 480 0 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal3 s 39200 25984 40000 26104 0 FreeSans 480 0 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal3 s 39200 27344 40000 27464 0 FreeSans 480 0 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal3 s 39200 2864 40000 2984 0 FreeSans 480 0 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal3 s 39200 28704 40000 28824 0 FreeSans 480 0 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal3 s 39200 30064 40000 30184 0 FreeSans 480 0 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal3 s 39200 31424 40000 31544 0 FreeSans 480 0 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal3 s 39200 32784 40000 32904 0 FreeSans 480 0 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal3 s 39200 34144 40000 34264 0 FreeSans 480 0 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal3 s 39200 35504 40000 35624 0 FreeSans 480 0 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal3 s 39200 36864 40000 36984 0 FreeSans 480 0 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal3 s 39200 4224 40000 4344 0 FreeSans 480 0 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal3 s 39200 5584 40000 5704 0 FreeSans 480 0 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal3 s 39200 6944 40000 7064 0 FreeSans 480 0 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal3 s 39200 8304 40000 8424 0 FreeSans 480 0 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal3 s 39200 9664 40000 9784 0 FreeSans 480 0 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal3 s 39200 11024 40000 11144 0 FreeSans 480 0 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal3 s 39200 12384 40000 12504 0 FreeSans 480 0 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal3 s 39200 13744 40000 13864 0 FreeSans 480 0 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
